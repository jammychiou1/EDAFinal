module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43);

  input in1, in3, in4, in6, in7, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90;

  input [1:0] in2, in8;

  input [4:0] in5;

  output [6:0] out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27;

  output [5:0] out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43;
  wire in1, in3, in4, in6, in7, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90;
  wire [1:0] in2, in8;
  wire [4:0] in5;
  wire [6:0] out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27;
  wire [5:0] out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43;
  wire w__1113, w__1117, w__1117, w__1145, w__1149, w__1149, w__7, w__1124;
  wire w__9, w__10, w__11, w__12, w__13, w__14, w__15, w__16;
  wire w__17, w__18, w__19, w__20, w__21, w__22, w__23, w__24;
  wire w__25, w__26, w__91, w__28, w__29, w__30, w__31, w__32;
  wire w__33, w__34, w__35, w__36, w__37, w__38, w__39, w__40;
  wire w__41, w__42, w__91, w__28, w__29, w__46, w__47, w__48;
  wire w__49, w__50, w__51, w__52, w__53, w__54, w__55, w__56;
  wire w__57, w__58, w__91, w__60, w__29, w__62, w__63, w__64;
  wire w__65, w__66, w__67, w__68, w__69, w__70, w__71, w__72;
  wire w__73, w__74, w__75, w__28, w__29, w__78, w__79, w__80;
  wire w__81, w__82, w__83, w__84, w__85, w__86, w__87, w__88;
  wire w__89, w__90, w__91, w__28, w__29, w__94, w__95, w__96;
  wire w__97, w__98, w__99, w__100, w__101, w__102, w__103, w__104;
  wire w__105, w__106, w__91, w__28, w__29, w__110, w__111, w__112;
  wire w__113, w__114, w__115, w__116, w__117, w__118, w__119, w__120;
  wire w__121, w__122, w__91, w__28, w__29, w__126, w__127, w__128;
  wire w__129, w__130, w__131, w__132, w__133, w__134, w__135, w__136;
  wire w__137, w__138, w__91, w__140, w__29, w__142, w__143, w__144;
  wire w__145, w__146, w__147, w__148, w__149, w__150, w__151, w__152;
  wire w__153, w__154, w__155, w__156, w__29, w__158, w__159, w__160;
  wire w__161, w__162, w__163, w__164, w__165, w__166, w__167, w__168;
  wire w__169, w__170, w__91, w__172, w__29, w__174, w__175, w__176;
  wire w__177, w__178, w__179, w__180, w__181, w__182, w__183, w__184;
  wire w__185, w__186, w__187, w__28, w__29, w__190, w__191, w__192;
  wire w__193, w__194, w__195, w__196, w__197, w__198, w__199, w__200;
  wire w__201, w__202, w__91, w__28, w__29, w__206, w__207, w__208;
  wire w__209, w__210, w__211, w__212, w__213, w__214, w__215, w__216;
  wire w__217, w__218, w__219, w__220, w__29, w__222, w__223, w__224;
  wire w__225, w__226, w__227, w__228, w__229, w__230, w__231, w__232;
  wire w__233, w__234, w__235, w__236, w__29, w__238, w__239, w__240;
  wire w__241, w__242, w__243, w__244, w__245, w__246, w__247, w__248;
  wire w__249, w__250, w__91, w__28, w__29, w__254, w__255, w__256;
  wire w__257, w__258, w__259, w__260, w__261, w__262, w__263, w__264;
  wire w__265, w__266, w__91, w__28, w__29, w__270, w__271, w__272;
  wire w__273, w__274, w__275, w__276, w__277, w__278, w__279, w__280;
  wire w__281, w__282, w__283, w__284, w__29, w__286, w__287, w__288;
  wire w__289, w__290, w__291, w__292, w__293, w__294, w__295, w__296;
  wire w__297, w__298, w__299, w__300, w__29, w__302, w__303, w__304;
  wire w__305, w__306, w__307, w__308, w__309, w__310, w__311, w__312;
  wire w__313, w__314, w__91, w__316, w__29, w__318, w__319, w__320;
  wire w__321, w__322, w__323, w__324, w__325, w__326, w__327, w__328;
  wire w__329, w__330, w__331, w__28, w__29, w__334, w__335, w__336;
  wire w__337, w__338, w__339, w__340, w__341, w__342, w__343, w__344;
  wire w__345, w__346, w__347, w__348, w__29, w__350, w__351, w__352;
  wire w__353, w__354, w__355, w__356, w__357, w__358, w__359, w__360;
  wire w__361, w__362, w__363, w__28, w__29, w__366, w__367, w__368;
  wire w__369, w__370, w__371, w__372, w__373, w__374, w__375, w__376;
  wire w__377, w__378, w__379, w__380, w__29, w__382, w__383, w__384;
  wire w__385, w__386, w__387, w__388, w__389, w__390, w__391, w__392;
  wire w__393, w__394, w__91, w__396, w__29, w__398, w__399, w__400;
  wire w__401, w__402, w__403, w__404, w__405, w__406, w__407, w__408;
  wire w__409, w__410, w__411, w__28, w__29, w__414, w__415, w__416;
  wire w__417, w__418, w__419, w__420, w__421, w__422, w__423, w__424;
  wire w__425, w__426, w__91, w__28, w__29, w__430, w__431, w__432;
  wire w__433, w__434, w__435, w__436, w__437, w__438, w__439, w__440;
  wire w__441, w__442, w__91, w__28, w__29, w__446, w__447, w__448;
  wire w__449, w__450, w__451, w__452, w__453, w__454, w__455, w__456;
  wire w__457, w__458, w__459, w__477, w__29, w__462, w__463, w__464;
  wire w__465, w__466, w__467, w__468, w__469, w__470, w__471, w__472;
  wire w__473, w__474, w__475, w__459, w__477, w__29, w__479, w__480;
  wire w__481, w__482, w__483, w__484, w__485, w__486, w__487, w__488;
  wire w__489, w__490, w__491, w__492, w__493, w__494, w__29, w__496;
  wire w__497, w__498, w__499, w__500, w__501, w__502, w__503, w__504;
  wire w__505, w__506, w__507, w__508, w__509, w__459, w__477, w__29;
  wire w__513, w__514, w__515, w__516, w__517, w__518, w__519, w__520;
  wire w__521, w__522, w__523, w__524, w__525, w__526, w__459, w__477;
  wire w__29, w__530, w__531, w__532, w__533, w__534, w__535, w__536;
  wire w__537, w__538, w__539, w__540, w__541, w__542, w__543, w__544;
  wire w__545, w__29, w__547, w__548, w__549, w__550, w__551, w__552;
  wire w__553, w__554, w__555, w__556, w__557, w__558, w__559, w__560;
  wire w__459, w__477, w__29, w__564, w__565, w__566, w__567, w__568;
  wire w__569, w__570, w__571, w__572, w__573, w__574, w__575, w__576;
  wire w__577, w__459, w__477, w__29, w__581, w__582, w__583, w__584;
  wire w__585, w__586, w__587, w__588, w__589, w__590, w__591, w__592;
  wire w__593, w__594, w__595, w__477, w__29, w__598, w__599, w__600;
  wire w__601, w__602, w__603, w__604, w__605, w__606, w__607, w__608;
  wire w__609, w__610, w__611, w__459, w__477, w__29, w__615, w__616;
  wire w__617, w__618, w__619, w__620, w__621, w__622, w__623, w__624;
  wire w__625, w__626, w__627, w__628, w__459, w__630, w__29, w__632;
  wire w__633, w__634, w__635, w__636, w__637, w__638, w__639, w__640;
  wire w__641, w__642, w__643, w__644, w__645, w__646, w__647, w__29;
  wire w__649, w__650, w__651, w__652, w__653, w__654, w__655, w__656;
  wire w__657, w__658, w__659, w__660, w__661, w__662, w__663, w__664;
  wire w__29, w__666, w__667, w__668, w__669, w__670, w__671, w__672;
  wire w__673, w__674, w__675, w__676, w__677, w__678, w__679, w__459;
  wire w__477, w__29, w__683, w__684, w__685, w__686, w__687, w__688;
  wire w__689, w__690, w__691, w__692, w__693, w__694, w__695, w__696;
  wire w__459, w__477, w__29, w__700, w__701, w__702, w__703, w__704;
  wire w__705, w__706, w__707, w__708, w__709, w__710, w__711, w__712;
  wire w__713, w__459, w__477, w__29, w__717, w__718, w__719, w__720;
  wire w__721, w__722, w__723, w__724, w__725, w__726, w__727, w__728;
  wire w__729, w__730, w__29, w__732, w__733, w__734, w__735, w__736;
  wire w__29, w__732, w__739, w__740, w__741, w__742, w__743, inc_add_183_20_n_1;
  wire inc_add_183_20_n_2, inc_add_183_20_n_3, inc_add_183_20_n_4, inc_add_183_20_n_5, inc_add_183_20_n_6, w__778, w__779, w__746;
  wire w__747, w__746, w__747, w__750, w__751, w__750, w__751, w__754;
  wire w__755, w__754, w__755, w__758, w__759, w__758, w__759, w__762;
  wire w__763, w__762, w__763, w__762, w__763, w__758, w__759, w__750;
  wire w__751, w__778, w__779, w__746, w__747, w__754, w__755, w__778;
  wire w__779, w__1081, w__1077, w__1079, w__1075, w__1083, w__1085, w__855;
  wire w__857, w__857, w__804, w__806, w__806, w__855, w__857, w__857;
  wire w__819, w__821, w__821, w__828, w__830, w__830, w__843, w__845;
  wire w__845, w__804, w__806, w__806, w__843, w__845, w__845, w__819;
  wire w__821, w__821, w__804, w__806, w__806, w__819, w__821, w__821;
  wire w__819, w__821, w__821, w__843, w__845, w__845, w__831, w__833;
  wire w__833, w__828, w__830, w__830, w__831, w__833, w__833, w__828;
  wire w__830, w__830, w__831, w__833, w__833, w__855, w__857, w__857;
  wire w__843, w__845, w__845, w__831, w__833, w__833, w__828, w__830;
  wire w__830, w__804, w__806, w__806, w__855, w__857, w__857, w__855;
  wire w__857, w__857, w__855, w__857, w__857, w__819, w__821, w__821;
  wire w__819, w__821, w__821, w__843, w__845, w__845, w__819, w__821;
  wire w__821, w__831, w__833, w__833, w__843, w__845, w__845, w__828;
  wire w__830, w__830, w__831, w__833, w__833, w__828, w__830, w__830;
  wire w__828, w__830, w__830, w__828, w__830, w__830, w__831, w__833;
  wire w__833, w__804, w__806, w__806, w__831, w__833, w__833, w__804;
  wire w__806, w__806, w__855, w__857, w__857, w__855, w__857, w__857;
  wire w__804, w__806, w__806, w__843, w__845, w__845, w__804, w__806;
  wire w__806, w__843, w__845, w__845, w__819, w__821, w__821, w__819;
  wire w__821, w__821, w__855, w__857, w__857, w__843, w__845, w__845;
  wire w__828, w__830, w__830, w__831, w__833, w__833, w__804, w__806;
  wire w__806, w__804, w__806, w__806, w__831, w__833, w__833, w__819;
  wire w__821, w__821, w__828, w__830, w__830, w__855, w__857, w__857;
  wire w__843, w__845, w__845, w__976, w__980, w__983, w__1023, w__1025;
  wire w__1050, w__1052, w__1053, w__1055, w__975, w__976, w__1128, w__1117;
  wire w__979, w__980, w__1149, w__982, w__983, w__976, w__1129, w__1129;
  wire w__1023, w__1025, w__1025, w__983, w__1150, w__1150, w__1050, w__1052;
  wire w__1052, w__1053, w__1055, w__1055, w__980, w__1118, w__1118, w__976;
  wire w__1129, w__1129, w__976, w__1129, w__1129, w__976, w__1129, w__1129;
  wire w__976, w__1129, w__1129, w__1023, w__1025, w__1025, w__1023, w__1025;
  wire w__1025, w__1023, w__1025, w__1025, w__1023, w__1025, w__1025, w__1053;
  wire w__1055, w__1055, w__983, w__1150, w__1150, w__983, w__1150, w__1150;
  wire w__983, w__1150, w__1150, w__983, w__1150, w__1150, w__1050, w__1052;
  wire w__1052, w__1050, w__1052, w__1052, w__1050, w__1052, w__1052, w__1050;
  wire w__1052, w__1052, w__1053, w__1055, w__1055, w__980, w__1118, w__1118;
  wire w__980, w__1118, w__1118, w__980, w__1118, w__1118, w__980, w__1118;
  wire w__1118, w__1053, w__1055, w__1055, w__1053, w__1055, w__1055, w__1074;
  wire w__1075, w__1076, w__1077, w__1078, w__1079, w__1080, w__1081, w__1082;
  wire w__1083, w__1084, w__1085, w__1075, w__1123, w__1077, w__1134, w__1079;
  wire w__1139, w__1085, w__1144, w__1081, w__1155, w__1083, w__1160, w__979;
  wire w__979, w__1118, w__1074, w__975, w__975, w__1129, w__1076, w__1078;
  wire w__1084, w__982, w__982, w__1150, w__1080, w__1082, w__1113, w__979;
  wire w__1118, w__1118, w__1117, w__1118, w__1123, w__1123, w__1123, w__1122;
  wire w__1123, w__1124, w__975, w__1129, w__1129, w__1128, w__1129, w__1134;
  wire w__1134, w__1134, w__1133, w__1134, w__1139, w__1139, w__1139, w__1138;
  wire w__1139, w__1144, w__1144, w__1144, w__1143, w__1144, w__1145, w__982;
  wire w__1150, w__1150, w__1149, w__1150, w__1155, w__1155, w__1155, w__1154;
  wire w__1155, w__1160, w__1160, w__1160, w__1159, w__1160, w__1161, w__1162;
  wire w__1163, w__1164, w__1165, w__1166, w__1167, w__1168, w__1169, w__1170;
  wire w__1171, w__1172, w__1173, w__1174, w__1175, w__1176, w__1177, w__1178;
  wire w__1179, w__1180, w__1181, w__1182, w__1183, w__1184, w__1185, w__1186;
  wire w__1187, w__1188, w__1189, w__1190, w__1191, w__1192, w__1193, w__1194;
  wire w__1195, w__1196, w__1197, w__1198, w__1199, w__1200, w__1201, w__1202;
  wire w__1203, w__1204, w__1205, w__1206, w__1207, w__1208, w__1209, w__1210;
  wire w__1211, w__1212, w__1213, w__1214, w__1215, w__1216, w__1217, w__1218;
  wire w__1219, w__1220, w__1221, w__1222, w__1223, w__1224, w__1225, w__1226;
  wire w__1227, w__1228, w__1229, w__1230, w__1231, w__1232, w__1233, w__1234;
  wire w__1235, w__1236, w__1237, w__1238, w__1239, w__1240, w__1241, w__1242;
  wire w__1243, w__1244, w__1245, w__1246, w__1247, w__1248, w__1249, w__1250;
  wire w__1251, w__1252, w__1253, w__1254, w__1255, w__1256, w__1257, w__1258;
  wire w__1259, w__1260, w__1261, w__1262, w__1263, w__1264, w__1265, w__1266;
  wire w__1267, w__1268, w__1269, w__1270, w__1271, w__1272, w__1273, w__1274;
  wire w__1275, w__1276, w__1277, w__1278, w__1279, w__1280, w__1281, w__1282;
  wire w__1283, w__1284, w__1285, w__1286, w__1287, w__1288, w__1289, w__1290;
  wire w__1291, w__1292, w__1293, w__1294, w__1295, w__1296, w__1297, w__1298;
  wire w__1299, w__1300, w__1301, w__1302, w__1303, w__1304, w__1305, w__1306;
  wire w__1307, w__1308, w__1309, w__1310, w__1311, w__1312, w__1313, w__1314;
  wire w__1315, w__1316, w__1317, w__1318, w__1319, w__1320, w__1321, w__1322;
  wire w__1323, w__1324, w__1325, w__1326, w__1327, w__1328, w__1329, w__1330;
  wire w__1331, w__1332, w__1333, w__1334, w__1335, w__1336, w__1337, w__1338;
  wire w__1339, w__1340, w__1341, w__1342, w__1343, w__1344, w__1345, w__1346;
  wire w__1347, w__1348, w__1349, w__1350, w__1351, w__1352, w__1353, w__1354;
  wire w__1355, w__1356, w__1357, w__1358, w__1359, w__1360, w__1361, w__1362;
  wire w__1363, w__1364, w__1365, w__1366, w__1367, w__1368, w__1369, w__1370;
  wire w__1371, w__1372, w__1373, w__1374, w__1375, w__1376, w__1377, w__1378;
  wire w__1379, w__1380, w__1381, w__1382, w__1383, w__1384, w__1385, w__1386;
  wire w__1387, w__1388, w__1389, w__1390, w__1391, w__1392, w__1393, w__1394;
  wire w__1395, w__1396, w__1397, w__1398, w__1399, w__1400, w__1401, w__1402;
  wire w__1403, w__1404, w__1405, w__1406, w__1407, w__1408, w__1409, w__1410;
  wire w__1411, w__1412, w__1413, w__1414, w__1415, w__1416, w__1417, w__1418;
  wire w__1419, w__1420, w__1421, w__1422, w__1423, w__1424, w__1425, w__1426;
  wire w__1427, w__1428, w__1429, w__1430, w__1431, w__1432, w__1433, w__1434;
  wire w__1435, w__1436, w__1437, w__1438, w__1439, w__1440, w__1441, w__1442;
  wire w__1443, w__1444, w__1445, w__1446, w__1447, w__1448, w__1449, w__1450;
  wire w__1451, w__1452, w__1453, w__1454, w__1455, w__1456, w__1457, w__1458;
  wire w__1459, w__1460, w__1461, w__1462, w__1463, w__1464, w__1465, w__1466;
  wire w__1467, w__1468, w__1469, w__1470, w__1471, w__1472, w__1473, w__1474;
  wire w__1475, w__1476, w__1477, w__1478, w__1479, w__1480, w__1481, w__1482;
  wire w__1483, w__1484, w__1485, w__1486, w__1487, w__1488, w__1489, w__1490;
  wire w__1491, w__1492, w__1493, w__1494, w__1495, w__1496, w__1497, w__1498;
  wire w__1499, w__1500, w__1501, w__1502, w__1503, w__1504, w__1505, w__1506;
  wire w__1507, w__1508, w__1509, w__1516, w__1509, w__1516, w__1513, w__1514;
  wire w__1509, w__1516, w__1527, w__1518, w__1519, w__1520, w__1527, w__1530;
  wire w__1523, w__1524, w__1525, w__1530, w__1527, w__1530, w__1527, w__1530;
  wire w__1531, w__1532, w__1533, w__1534, w__1535, w__1536, w__1537, w__1538;
  wire w__1539, w__1540, w__1541, w__1542, w__1543, w__1544, w__1545, w__1546;
  wire w__1547, w__1548, w__1549, w__1550, w__1551, w__1552, w__1553, w__1554;
  wire w__1555, w__1556, w__1557, w__1558, w__1559, w__1560, w__1561, w__1562;
  wire w__1563, w__1564, w__1565, w__1566, w__1567, w__1568, w__1569, w__1570;
  wire w__1571, w__1572, w__1573, w__1574, w__1575, w__1576, w__1577, w__1578;
  wire w__1579, w__1580, w__1581, w__1582, w__1583, w__1584, w__1585, w__1586;
  wire w__1587, w__1588, w__1589, w__1590, w__1591, w__1592, w__1593, w__1594;
  wire w__1595, w__1596, w__1597, w__1598, w__1599, w__1600, w__1601, w__1602;
  wire w__1603, w__1604, w__1605, w__1606, w__1607, w__1608, w__1609, w__1610;
  wire w__1611, w__1612, w__1613, w__1614, w__1615, w__1616, w__1617, w__1618;
  wire w__1619, w__1620, w__1621, w__1622, w__1623, w__1624, w__1625, w__1626;
  wire w__1627, w__1628, w__1629, w__1630, w__1631, w__1632, w__1633, w__1634;
  wire w__1635, w__1636, w__1637, w__1638, w__1639, w__1640, w__1641, w__1642;
  wire w__1643, w__1644, w__1645, w__1646, w__1647, w__1648, w__1649, w__1650;
  wire w__1651, w__1652, w__1653, w__1654, w__1655, w__1656, w__1657, w__1658;
  wire w__1659, w__1660, w__1661, w__1662, w__1663, w__1664, w__1665, w__1666;
  wire w__1667, w__1668, w__1669, w__1670, w__1671, w__1672, w__1673, w__1674;
  wire w__1675, w__1676, w__1677, w__1678, w__1679, w__1680, w__1681, w__1682;
  wire w__1683, w__1684, w__1685, w__1686, w__1687, w__1688, w__1689, w__1690;
  not g__1(w__1527 ,w__1507);
  not g__2(w__1530 ,w__1508);
  not g__5(w__1520 ,w__1508);
  not g__6(w__1509 ,w__1506);
  not g__7(w__1519 ,w__1507);
  not g__10(w__1516 ,w__1505);
  not g__12(w__1524 ,w__1508);
  not g__13(w__1523 ,w__1507);
  not g__14(w__1513 ,w__1506);
  not g__18(w__1514 ,w__1505);
  not g__19(w__1518 ,w__1508);
  not g__21(w__1525 ,w__1507);
  not g__23(w__1505 ,w__1592);
  not g__24(w__1507 ,w__1676);
  not g__25(w__1506 ,w__1591);
  not g__26(w__1508 ,w__1677);
  or g__27(out32[0] ,w__1373 ,w__1472);
  or g__28(out2[2] ,w__1285 ,w__1455);
  or g__29(out3[0] ,w__1308 ,w__1479);
  or g__30(out6[0] ,w__1348 ,w__1498);
  or g__31(out7[2] ,w__1343 ,w__1488);
  or g__32(out13[1] ,w__1333 ,w__1500);
  or g__33(out26[2] ,w__1356 ,w__1502);
  or g__34(out26[1] ,w__1337 ,w__1501);
  or g__35(out13[0] ,w__1341 ,w__1494);
  or g__36(out26[0] ,w__1332 ,w__1499);
  or g__37(out27[2] ,w__1329 ,w__1496);
  or g__38(out27[1] ,w__1342 ,w__1495);
  or g__39(out7[1] ,w__1290 ,w__1485);
  or g__40(out14[2] ,w__1346 ,w__1490);
  or g__41(out27[0] ,w__1344 ,w__1493);
  or g__42(out28[1] ,w__1314 ,w__1491);
  or g__43(out14[1] ,w__1303 ,w__1487);
  or g__44(out28[0] ,w__1349 ,w__1489);
  or g__45(out29[1] ,w__1351 ,w__1486);
  or g__46(out4[2] ,w__1371 ,w__1461);
  or g__47(out7[0] ,w__1364 ,w__1474);
  or g__48(out14[0] ,w__1355 ,w__1482);
  or g__49(out29[0] ,w__1293 ,w__1484);
  or g__50(out30[1] ,w__1289 ,w__1483);
  or g__51(out15[2] ,w__1360 ,w__1477);
  or g__52(out30[0] ,w__1359 ,w__1481);
  or g__53(out15[1] ,w__1244 ,w__1476);
  or g__54(out31[1] ,w__1362 ,w__1480);
  or g__55(out31[0] ,w__1366 ,w__1475);
  or g__56(out8[2] ,w__1246 ,w__1464);
  or g__57(out15[0] ,w__1374 ,w__1471);
  or g__58(out32[1] ,w__1369 ,w__1473);
  or g__59(out1[2] ,w__1237 ,w__1497);
  or g__60(out16[2] ,w__1247 ,w__1466);
  or g__61(out33[1] ,w__1188 ,w__1470);
  or g__62(out33[0] ,w__1168 ,w__1469);
  or g__63(out34[1] ,w__1236 ,w__1467);
  or g__64(out2[1] ,w__1197 ,w__1444);
  or g__65(out4[1] ,w__1257 ,w__1449);
  or g__66(out8[1] ,w__1169 ,w__1458);
  or g__67(out16[1] ,w__1163 ,w__1463);
  or g__68(out34[0] ,w__1323 ,w__1465);
  or g__69(out35[1] ,w__1319 ,w__1462);
  or g__70(out16[0] ,w__1164 ,w__1459);
  or g__71(out35[0] ,w__1216 ,w__1460);
  or g__72(out17[2] ,w__1231 ,w__1454);
  or g__73(out36[1] ,w__1174 ,w__1457);
  or g__74(out8[0] ,w__1180 ,w__1452);
  or g__75(out17[1] ,w__1261 ,w__1450);
  or g__76(out36[0] ,w__1187 ,w__1456);
  or g__77(out37[1] ,w__1177 ,w__1453);
  or g__78(out9[2] ,w__1186 ,w__1441);
  or g__79(out37[0] ,w__1211 ,w__1451);
  or g__80(out38[1] ,w__1262 ,w__1448);
  or g__81(out17[0] ,w__1178 ,w__1446);
  or g__82(out38[0] ,w__1225 ,w__1447);
  or g__83(out4[0] ,w__1267 ,w__1433);
  or g__84(out9[1] ,w__1271 ,w__1437);
  or g__85(out18[2] ,w__1265 ,w__1442);
  or g__86(out39[1] ,w__1183 ,w__1445);
  or g__87(out39[0] ,w__1204 ,w__1443);
  or g__88(out18[1] ,w__1185 ,w__1439);
  or g__89(out40[1] ,w__1268 ,w__1440);
  or g__90(out40[0] ,w__1200 ,w__1438);
  or g__91(out25[0] ,w__1328 ,w__1408);
  or g__92(out18[0] ,w__1189 ,w__1434);
  or g__93(out41[1] ,w__1228 ,w__1436);
  or g__94(out19[2] ,w__1196 ,w__1430);
  or g__95(out41[0] ,w__1275 ,w__1435);
  or g__96(out42[1] ,w__1195 ,w__1432);
  or g__97(out9[0] ,w__1270 ,w__1427);
  or g__98(out42[0] ,w__1192 ,w__1431);
  or g__99(out19[1] ,w__1227 ,w__1428);
  or g__100(out43[1] ,w__1269 ,w__1429);
  or g__101(out1[1] ,w__1336 ,w__1468);
  or g__102(out1[0] ,w__1310 ,w__1388);
  or g__103(out2[0] ,w__1256 ,w__1504);
  or g__104(out10[2] ,w__1230 ,w__1421);
  or g__105(out19[0] ,w__1279 ,w__1425);
  or g__106(out43[0] ,w__1238 ,w__1426);
  or g__107(out20[2] ,w__1281 ,w__1423);
  or g__108(w__1531 ,w__1260 ,w__1424);
  or g__109(out5[1] ,w__1205 ,w__1414);
  or g__110(out10[1] ,w__1273 ,w__1415);
  or g__111(out20[1] ,w__1202 ,w__1420);
  or g__112(w__1535 ,w__1255 ,w__1422);
  or g__113(w__1539 ,w__1300 ,w__1418);
  or g__114(out20[0] ,w__1203 ,w__1416);
  or g__115(out21[2] ,w__1179 ,w__1412);
  or g__116(w__1543 ,w__1243 ,w__1478);
  or g__117(out3[2] ,w__1214 ,w__1380);
  or g__118(out10[0] ,w__1276 ,w__1409);
  or g__119(out21[1] ,w__1368 ,w__1411);
  or g__120(w__1547 ,w__1282 ,w__1413);
  or g__121(out11[2] ,w__1350 ,w__1403);
  or g__122(w__1551 ,w__1325 ,w__1410);
  or g__123(out21[0] ,w__1309 ,w__1406);
  or g__124(w__1555 ,w__1305 ,w__1407);
  or g__125(out5[0] ,w__1210 ,w__1395);
  or g__126(out22[2] ,w__1298 ,w__1404);
  or g__127(w__1559 ,w__1327 ,w__1405);
  or g__128(out11[1] ,w__1306 ,w__1400);
  or g__129(out22[1] ,w__1222 ,w__1401);
  or g__130(w__1563 ,w__1162 ,w__1402);
  or g__131(out3[1] ,w__1338 ,w__1492);
  or g__132(out6[2] ,w__1206 ,w__1383);
  or g__133(out11[0] ,w__1172 ,w__1392);
  or g__134(out22[0] ,w__1322 ,w__1398);
  or g__135(w__1567 ,w__1212 ,w__1399);
  or g__136(out23[2] ,w__1217 ,w__1394);
  or g__137(w__1571 ,w__1315 ,w__1397);
  or g__138(out23[1] ,w__1171 ,w__1393);
  or g__139(w__1575 ,w__1170 ,w__1396);
  or g__140(out12[2] ,w__1299 ,w__1385);
  or g__141(out23[0] ,w__1313 ,w__1390);
  or g__142(w__1579 ,w__1198 ,w__1391);
  or g__143(out24[2] ,w__1316 ,w__1386);
  or g__144(w__1583 ,w__1176 ,w__1389);
  or g__145(w__1587 ,w__1292 ,w__1387);
  or g__146(out6[1] ,w__1161 ,w__1376);
  or g__147(out12[1] ,w__1220 ,w__1381);
  or g__148(out24[1] ,w__1181 ,w__1384);
  or g__149(w__1594 ,w__1264 ,w__1417);
  or g__150(out24[0] ,w__1321 ,w__1382);
  or g__151(out25[2] ,w__1167 ,w__1379);
  or g__152(out12[0] ,w__1324 ,w__1378);
  or g__153(out25[1] ,w__1326 ,w__1377);
  or g__154(out13[2] ,w__1357 ,w__1503);
  or g__155(out5[2] ,w__1232 ,w__1419);
  nor g__156(w__1504 ,w__1025 ,in9);
  nor g__157(w__1503 ,w__1055 ,in31);
  nor g__158(w__1502 ,w__1118 ,in57);
  nor g__159(w__1501 ,w__1052 ,in57);
  nor g__160(w__1500 ,w__1150 ,in31);
  nor g__161(w__1499 ,w__1129 ,in57);
  nor g__162(w__1498 ,w__1025 ,in17);
  nor g__163(w__1497 ,w__1055 ,in6);
  nor g__164(w__1496 ,w__1118 ,in59);
  nor g__165(w__1495 ,w__1052 ,in59);
  nor g__166(w__1494 ,w__1129 ,in31);
  nor g__167(w__1493 ,w__1025 ,in59);
  nor g__168(w__1492 ,w__1150 ,in11);
  nor g__169(w__1491 ,w__1052 ,in61);
  nor g__170(w__1490 ,w__1055 ,in33);
  nor g__171(w__1489 ,w__1129 ,in61);
  nor g__172(w__1488 ,w__1118 ,in19);
  nor g__173(w__1487 ,w__1150 ,in33);
  nor g__174(w__1486 ,w__1150 ,in3);
  nor g__175(w__1485 ,w__1150 ,in19);
  nor g__176(w__1484 ,w__1129 ,in3);
  nor g__177(w__1483 ,w__1052 ,in63);
  nor g__178(w__1482 ,w__1129 ,in33);
  nor g__179(w__1481 ,w__1025 ,in63);
  nor g__180(w__1480 ,w__1052 ,in65);
  nor g__181(w__1479 ,w__1025 ,in11);
  nor g__182(w__1478 ,w__1118 ,in83);
  nor g__183(w__1477 ,w__1118 ,in35);
  nor g__184(w__1476 ,w__1150 ,in35);
  nor g__185(w__1475 ,w__1129 ,in65);
  nor g__186(w__1474 ,w__1129 ,in19);
  nor g__187(w__1473 ,w__1150 ,in67);
  nor g__188(w__1472 ,w__1025 ,in67);
  nor g__189(w__1471 ,w__1129 ,in35);
  nor g__190(w__1470 ,w__1052 ,in69);
  nor g__191(w__1469 ,w__1129 ,in69);
  nor g__192(w__1468 ,w__1150 ,in6);
  nor g__193(w__1467 ,w__1150 ,in71);
  nor g__194(w__1466 ,w__1055 ,in37);
  nor g__195(w__1465 ,w__1025 ,in71);
  nor g__196(w__1464 ,w__1055 ,in21);
  nor g__197(w__1463 ,w__1052 ,in37);
  nor g__198(w__1462 ,w__1150 ,in73);
  nor g__199(w__1461 ,w__1118 ,in13);
  nor g__200(w__1460 ,w__1129 ,in73);
  nor g__201(w__1459 ,w__1025 ,in37);
  nor g__202(w__1458 ,w__1052 ,in21);
  nor g__203(w__1457 ,w__1150 ,in75);
  nor g__204(w__1456 ,w__1129 ,in75);
  nor g__205(w__1455 ,w__1118 ,in9);
  nor g__206(w__1454 ,w__1055 ,in39);
  nor g__207(w__1453 ,w__1052 ,in77);
  nor g__208(w__1452 ,w__1025 ,in21);
  nor g__209(w__1451 ,w__1025 ,in77);
  nor g__210(w__1450 ,w__1052 ,in39);
  nor g__211(w__1449 ,w__1150 ,in13);
  nor g__212(w__1448 ,w__1052 ,in79);
  nor g__213(w__1447 ,w__1129 ,in79);
  nor g__214(w__1446 ,w__1025 ,in39);
  nor g__215(w__1445 ,w__1052 ,in81);
  nor g__216(w__1444 ,w__1052 ,in9);
  nor g__217(w__1443 ,w__1025 ,in81);
  nor g__218(w__1442 ,w__1118 ,in41);
  nor g__219(w__1441 ,w__1118 ,in23);
  nor g__220(w__1440 ,w__1150 ,in83);
  nor g__221(w__1439 ,w__1150 ,in41);
  nor g__222(w__1438 ,w__1025 ,in83);
  nor g__223(w__1437 ,w__1052 ,in23);
  nor g__224(w__1436 ,w__1052 ,in85);
  nor g__225(w__1435 ,w__1129 ,in85);
  nor g__226(w__1434 ,w__1129 ,in41);
  nor g__227(w__1433 ,w__1025 ,in13);
  nor g__228(w__1432 ,w__1150 ,in87);
  nor g__229(w__1431 ,w__1025 ,in87);
  nor g__230(w__1430 ,w__1055 ,in43);
  nor g__231(w__1429 ,w__1150 ,in89);
  nor g__232(w__1428 ,w__1052 ,in43);
  nor g__233(w__1427 ,w__1129 ,in23);
  nor g__234(w__1426 ,w__1129 ,in89);
  nor g__235(w__1425 ,w__1025 ,in43);
  nor g__236(w__1424 ,w__1118 ,in89);
  nor g__237(w__1423 ,w__1055 ,in45);
  nor g__238(w__1422 ,w__1118 ,in87);
  nor g__239(w__1421 ,w__1055 ,in25);
  nor g__240(w__1420 ,w__1150 ,in45);
  nor g__241(w__1419 ,w__1055 ,in15);
  nor g__242(w__1418 ,w__1118 ,in85);
  nor g__243(w__1417 ,w__1055 ,in61);
  nor g__244(w__1416 ,w__1129 ,in45);
  nor g__245(w__1415 ,w__1052 ,in25);
  nor g__246(w__1414 ,w__1150 ,in15);
  nor g__247(w__1413 ,w__1055 ,in81);
  nor g__248(w__1412 ,w__1055 ,in47);
  nor g__249(w__1411 ,w__1150 ,in47);
  nor g__250(w__1410 ,w__1118 ,in79);
  nor g__251(w__1409 ,w__1025 ,in25);
  nor g__252(w__1408 ,w__1129 ,in55);
  nor g__253(w__1407 ,w__1118 ,in77);
  nor g__254(w__1406 ,w__1129 ,in47);
  nor g__255(w__1405 ,w__1055 ,in75);
  nor g__256(w__1404 ,w__1055 ,in49);
  nor g__257(w__1403 ,w__1118 ,in27);
  nor g__258(w__1402 ,w__1118 ,in73);
  nor g__259(w__1401 ,w__1052 ,in49);
  nor g__260(w__1400 ,w__1052 ,in27);
  nor g__261(w__1399 ,w__1055 ,in71);
  nor g__262(w__1398 ,w__1025 ,in49);
  nor g__263(w__1397 ,w__1118 ,in69);
  nor g__264(w__1396 ,w__1055 ,in67);
  nor g__265(w__1395 ,w__1025 ,in15);
  nor g__266(w__1394 ,w__1118 ,in51);
  nor g__267(w__1393 ,w__1052 ,in51);
  nor g__268(w__1392 ,w__1025 ,in27);
  nor g__269(w__1391 ,w__1118 ,in65);
  nor g__270(w__1390 ,w__1025 ,in51);
  nor g__271(w__1389 ,w__1055 ,in63);
  nor g__272(w__1388 ,w__1129 ,in6);
  nor g__273(w__1387 ,w__1055 ,in3);
  nor g__274(w__1386 ,w__1055 ,in53);
  nor g__275(w__1385 ,w__1055 ,in29);
  nor g__276(w__1384 ,w__1052 ,in53);
  nor g__277(w__1383 ,w__1118 ,in17);
  nor g__278(w__1382 ,w__1025 ,in53);
  nor g__279(w__1381 ,w__1150 ,in29);
  nor g__280(w__1380 ,w__1055 ,in11);
  nor g__281(w__1379 ,w__1118 ,in55);
  nor g__282(w__1378 ,w__1129 ,in29);
  nor g__283(w__1377 ,w__1052 ,in55);
  nor g__284(w__1376 ,w__1150 ,in17);
  and g__285(w__1375 ,in49 ,w__830);
  and g__286(w__1374 ,in35 ,w__821);
  and g__287(w__1373 ,in67 ,w__821);
  and g__288(w__1372 ,in23 ,w__845);
  and g__289(w__1371 ,in13 ,w__806);
  and g__290(w__1370 ,in59 ,w__845);
  and g__291(w__1369 ,in67 ,w__833);
  and g__292(w__1368 ,in47 ,w__833);
  and g__293(w__1367 ,in53 ,w__830);
  and g__294(w__1366 ,in65 ,w__821);
  and g__295(w__1365 ,in6 ,w__845);
  and g__296(w__1364 ,in19 ,w__821);
  and g__297(w__1363 ,in43 ,w__830);
  and g__298(w__1362 ,in65 ,w__833);
  and g__299(w__1361 ,in43 ,w__845);
  and g__300(w__1360 ,in35 ,w__806);
  and g__301(w__1359 ,in63 ,w__821);
  and g__302(w__1658 ,in19 ,w__857);
  and g__303(w__1358 ,in17 ,w__830);
  and g__304(w__1357 ,in31 ,w__806);
  and g__305(w__1356 ,in57 ,w__806);
  and g__306(w__1661 ,in17 ,w__857);
  and g__307(w__1355 ,in33 ,w__821);
  and g__308(w__1354 ,in41 ,w__845);
  and g__309(w__1353 ,in39 ,w__830);
  and g__310(w__1352 ,in77 ,w__857);
  and g__311(w__1643 ,in29 ,w__857);
  and g__312(w__1351 ,in3 ,w__833);
  and g__313(w__1670 ,in11 ,w__857);
  and g__314(w__1350 ,in27 ,w__806);
  and g__315(w__1349 ,in61 ,w__821);
  and g__316(w__1348 ,in17 ,w__821);
  and g__317(w__1679 ,in6 ,w__857);
  and g__318(w__1347 ,in13 ,w__845);
  and g__319(w__1664 ,in15 ,w__857);
  and g__320(w__1346 ,in33 ,w__806);
  and g__321(w__1345 ,in17 ,w__845);
  and g__322(w__1344 ,in59 ,w__821);
  and g__323(w__1343 ,in19 ,w__806);
  and g__324(w__1342 ,in59 ,w__833);
  and g__325(w__1652 ,in23 ,w__857);
  and g__326(w__1566 ,in73 ,w__830);
  and g__327(w__1341 ,in31 ,w__821);
  and g__328(w__1646 ,in27 ,w__857);
  and g__329(w__1340 ,in15 ,w__830);
  and g__330(w__1339 ,in6 ,w__830);
  and g__331(w__1338 ,in11 ,w__833);
  and g__332(w__1337 ,in57 ,w__833);
  and g__333(w__1336 ,in6 ,w__833);
  and g__334(w__1335 ,in75 ,w__857);
  and g__335(w__1334 ,in73 ,w__845);
  and g__336(w__1673 ,in9 ,w__857);
  and g__337(w__1333 ,in31 ,w__833);
  and g__338(w__1332 ,in57 ,w__821);
  and g__339(w__1331 ,in9 ,w__830);
  and g__340(w__1330 ,in9 ,w__845);
  and g__341(w__1329 ,in59 ,w__806);
  and g__342(w__1328 ,in55 ,w__821);
  and g__343(w__1327 ,in75 ,w__806);
  and g__344(w__1570 ,in71 ,w__830);
  and g__345(w__1326 ,in55 ,w__833);
  and g__346(w__1325 ,in79 ,w__806);
  and g__347(w__1324 ,in29 ,w__821);
  and g__348(w__1562 ,in75 ,w__830);
  and g__349(w__1550 ,in81 ,w__830);
  and g__350(w__1323 ,in71 ,w__821);
  and g__351(w__1322 ,in49 ,w__821);
  and g__352(w__1321 ,in53 ,w__821);
  and g__353(w__1320 ,in11 ,w__845);
  and g__354(w__1319 ,in73 ,w__833);
  and g__355(w__1667 ,in13 ,w__857);
  and g__356(w__1318 ,in75 ,w__845);
  and g__357(w__1317 ,in11 ,w__830);
  and g__358(w__1316 ,in53 ,w__806);
  and g__359(w__1590 ,in3 ,w__830);
  and g__360(w__1315 ,in69 ,w__806);
  and g__361(w__1314 ,in61 ,w__833);
  and g__362(w__1313 ,in51 ,w__821);
  and g__363(w__1312 ,in65 ,w__857);
  and g__364(w__1311 ,in67 ,w__857);
  and g__365(w__1582 ,in65 ,w__830);
  and g__366(w__1310 ,in6 ,w__821);
  and g__367(w__1309 ,in47 ,w__821);
  and g__368(w__1578 ,in67 ,w__830);
  and g__369(w__1308 ,in11 ,w__821);
  and g__370(w__1307 ,in65 ,w__845);
  and g__371(w__1306 ,in27 ,w__833);
  and g__372(w__1305 ,in77 ,w__806);
  and g__373(w__1304 ,in13 ,w__830);
  and g__374(w__1303 ,in33 ,w__833);
  and g__375(w__1302 ,in77 ,w__845);
  and g__376(w__1301 ,in73 ,w__857);
  and g__377(w__1300 ,in85 ,w__806);
  and g__378(w__1299 ,in29 ,w__806);
  and g__379(w__1298 ,in49 ,w__806);
  and g__380(w__1297 ,in79 ,w__845);
  and g__381(w__1296 ,in21 ,w__830);
  and g__382(w__1295 ,in3 ,w__857);
  and g__383(w__1558 ,in77 ,w__830);
  and g__384(w__1294 ,in3 ,w__845);
  and g__385(w__1293 ,in3 ,w__821);
  and g__386(w__1554 ,in79 ,w__830);
  and g__387(w__1292 ,in3 ,w__806);
  and g__388(w__1291 ,in19 ,w__845);
  and g__389(w__1290 ,in19 ,w__833);
  and g__390(w__1289 ,in63 ,w__833);
  and g__391(w__1288 ,in27 ,w__830);
  and g__392(w__1287 ,in81 ,w__857);
  and g__393(w__1286 ,in21 ,w__845);
  and g__394(w__1285 ,in9 ,w__806);
  and g__395(w__1284 ,in19 ,w__830);
  and g__396(w__1283 ,in59 ,w__830);
  and g__397(w__1282 ,in81 ,w__806);
  and g__398(w__1538 ,in87 ,w__830);
  and g__399(w__1281 ,in45 ,w__806);
  and g__400(w__1280 ,in55 ,w__830);
  and g__401(w__1655 ,in21 ,w__857);
  and g__402(w__1279 ,in43 ,w__821);
  and g__403(w__1278 ,in61 ,w__845);
  and g__404(w__1277 ,in55 ,w__845);
  and g__405(w__1276 ,in25 ,w__821);
  and g__406(w__1275 ,in85 ,w__821);
  and g__407(w__1610 ,in51 ,w__857);
  and g__408(w__1274 ,in51 ,w__845);
  and g__409(w__1273 ,in25 ,w__833);
  and g__410(w__1272 ,in47 ,w__845);
  and g__411(w__1616 ,in47 ,w__857);
  and g__412(w__1613 ,in49 ,w__857);
  and g__413(w__1271 ,in23 ,w__833);
  and g__414(w__1270 ,in23 ,w__821);
  and g__415(w__1269 ,in89 ,w__833);
  and g__416(w__1268 ,in83 ,w__833);
  and g__417(w__1267 ,in13 ,w__821);
  and g__418(w__1266 ,in41 ,w__830);
  and g__419(w__1265 ,in41 ,w__806);
  and g__420(w__1622 ,in43 ,w__857);
  and g__421(w__1264 ,in61 ,w__806);
  and g__422(w__1263 ,in89 ,w__845);
  and g__423(w__1262 ,in79 ,w__833);
  and g__424(w__1631 ,in37 ,w__857);
  and g__425(w__1261 ,in39 ,w__833);
  and g__426(w__1260 ,in89 ,w__806);
  and g__427(w__1259 ,in35 ,w__845);
  and g__428(w__1258 ,in35 ,w__830);
  and g__429(w__1257 ,in13 ,w__833);
  and g__430(w__1256 ,in9 ,w__821);
  and g__431(w__1255 ,in87 ,w__806);
  and g__432(w__1254 ,in33 ,w__845);
  and g__433(w__1253 ,in31 ,w__845);
  and g__434(w__1252 ,in85 ,w__857);
  and g__435(w__1251 ,in29 ,w__830);
  and g__436(w__1250 ,in33 ,w__751);
  and g__437(w__1249 ,in27 ,w__845);
  and g__438(w__1248 ,in25 ,w__751);
  and g__439(w__1247 ,in37 ,w__806);
  and g__440(w__1246 ,in21 ,w__806);
  and g__441(w__1649 ,in25 ,w__857);
  and g__442(w__1245 ,in23 ,w__830);
  and g__443(w__1244 ,in35 ,w__833);
  and g__444(w__1243 ,in83 ,w__806);
  and g__445(w__1242 ,in81 ,w__845);
  and g__446(w__1241 ,in15 ,w__845);
  and g__447(w__1546 ,in83 ,w__751);
  and g__448(w__1240 ,in83 ,w__857);
  and g__449(w__1239 ,in83 ,w__779);
  and g__450(w__1238 ,in89 ,w__821);
  and g__451(w__1542 ,in85 ,w__830);
  and g__452(w__1625 ,in41 ,w__857);
  and g__453(w__1237 ,in6 ,w__806);
  and g__454(w__1236 ,in71 ,w__833);
  and g__455(w__1235 ,in85 ,w__779);
  and g__456(w__1234 ,in87 ,w__845);
  and g__457(w__1598 ,in59 ,w__857);
  and g__458(w__1233 ,in87 ,w__747);
  and g__459(w__1232 ,in15 ,w__763);
  and g__460(w__1634 ,in35 ,w__747);
  and g__461(w__1231 ,in39 ,w__763);
  and g__462(w__1230 ,in25 ,w__806);
  and g__463(w__1534 ,in89 ,w__830);
  and g__464(w__1229 ,in37 ,w__779);
  and g__465(w__1628 ,in39 ,w__857);
  and g__466(w__1228 ,in85 ,w__833);
  and g__467(w__1227 ,in43 ,w__833);
  and g__468(w__1226 ,in45 ,w__845);
  and g__469(w__1225 ,in79 ,w__755);
  and g__470(w__1224 ,in71 ,w__845);
  and g__471(w__1223 ,in25 ,w__845);
  and g__472(w__1222 ,in49 ,w__833);
  and g__473(w__1221 ,in53 ,w__845);
  and g__474(w__1640 ,in31 ,w__747);
  and g__475(w__1220 ,in29 ,w__759);
  and g__476(w__1219 ,in69 ,w__779);
  and g__477(w__1218 ,in71 ,w__857);
  and g__478(w__1217 ,in51 ,w__763);
  and g__479(w__1216 ,in73 ,w__755);
  and g__480(w__1637 ,in33 ,w__857);
  and g__481(w__1215 ,in67 ,w__845);
  and g__482(w__1607 ,in53 ,w__857);
  and g__483(w__1214 ,in11 ,w__806);
  and g__484(w__1213 ,in69 ,w__857);
  and g__485(w__1212 ,in71 ,w__806);
  and g__486(w__1211 ,in77 ,w__821);
  and g__487(w__1210 ,in15 ,w__755);
  and g__488(w__1209 ,in39 ,w__779);
  and g__489(w__1586 ,in63 ,w__830);
  and g__490(w__1208 ,in37 ,w__830);
  and g__491(w__1207 ,in79 ,w__747);
  and g__492(w__1206 ,in17 ,w__806);
  and g__493(w__1205 ,in15 ,w__759);
  and g__494(w__1204 ,in81 ,w__821);
  and g__495(w__1203 ,in45 ,w__821);
  and g__496(w__1202 ,in45 ,w__833);
  and g__497(w__1201 ,in57 ,w__751);
  and g__498(w__1200 ,in83 ,w__821);
  and g__499(w__1199 ,in89 ,w__857);
  and g__500(w__1198 ,in65 ,w__806);
  and g__501(w__1604 ,in55 ,w__747);
  and g__502(w__1197 ,in9 ,w__759);
  and g__503(w__1196 ,in43 ,w__763);
  and g__504(w__1195 ,in87 ,w__833);
  and g__505(w__1194 ,in45 ,w__830);
  and g__506(w__1193 ,in49 ,w__845);
  and g__507(w__1619 ,in45 ,w__857);
  and g__508(w__1192 ,in87 ,w__821);
  and g__509(w__1191 ,in47 ,w__751);
  and g__510(w__1190 ,in51 ,w__830);
  and g__511(w__1189 ,in41 ,w__755);
  and g__512(w__1188 ,in69 ,w__833);
  and g__513(w__1187 ,in75 ,w__821);
  and g__514(w__1186 ,in23 ,w__806);
  and g__515(w__1185 ,in41 ,w__833);
  and g__516(w__1184 ,in57 ,w__779);
  and g__517(w__1601 ,in57 ,w__747);
  and g__518(w__1183 ,in81 ,w__833);
  and g__519(w__1182 ,in61 ,w__857);
  and g__520(w__1181 ,in53 ,w__759);
  and g__521(w__1180 ,in21 ,w__755);
  and g__522(w__1597 ,in61 ,w__751);
  and g__523(w__1179 ,in47 ,w__763);
  and g__524(w__1178 ,in39 ,w__821);
  and g__525(w__1177 ,in77 ,w__833);
  and g__526(w__1176 ,in63 ,w__806);
  and g__527(w__1175 ,in63 ,w__845);
  and g__528(w__1174 ,in75 ,w__759);
  and g__529(w__1173 ,in63 ,w__857);
  and g__530(w__1172 ,in27 ,w__755);
  and g__531(w__1171 ,in51 ,w__833);
  and g__532(w__1170 ,in67 ,w__763);
  and g__533(w__1169 ,in21 ,w__759);
  and g__534(w__1168 ,in69 ,w__821);
  and g__535(w__1167 ,in55 ,w__806);
  and g__536(w__1166 ,in29 ,w__845);
  and g__537(w__1574 ,in69 ,w__830);
  and g__538(w__1165 ,in31 ,w__830);
  and g__539(w__1164 ,in37 ,w__821);
  and g__540(w__1163 ,in37 ,w__833);
  and g__541(w__1162 ,in73 ,w__806);
  and g__542(w__1161 ,in17 ,w__833);
  not g__543(w__1160 ,w__1083);
  not g__547(w__1159 ,w__1686);
  not g__548(w__1155 ,w__1081);
  not g__552(w__1154 ,w__1683);
  not g__553(w__1150 ,w__983);
  not g__555(w__1149 ,w__1145);
  not g__560(w__1145 ,w__1689);
  not g__561(w__1144 ,w__1085);
  not g__565(w__1143 ,w__1685);
  not g__566(w__1139 ,w__1079);
  not g__570(w__1138 ,w__1684);
  not g__571(w__1134 ,w__1077);
  not g__575(w__1133 ,w__1687);
  not g__576(w__1129 ,w__976);
  not g__578(w__1128 ,w__1124);
  not g__583(w__1124 ,w__1688);
  not g__584(w__1123 ,w__1075);
  not g__588(w__1122 ,w__1682);
  not g__589(w__1118 ,w__980);
  not g__591(w__1117 ,w__1113);
  not g__596(w__1113 ,w__1690);
  not g__609(w__1085 ,w__1084);
  not g__610(w__1084 ,w__1143);
  not g__611(w__1083 ,w__1082);
  not g__612(w__1082 ,w__1159);
  not g__613(w__1081 ,w__1080);
  not g__614(w__1080 ,w__1154);
  not g__615(w__1079 ,w__1078);
  not g__616(w__1078 ,w__1138);
  not g__617(w__1077 ,w__1076);
  not g__618(w__1076 ,w__1133);
  not g__619(w__1075 ,w__1074);
  not g__620(w__1074 ,w__1122);
  not g__639(w__1055 ,w__1053);
  not g__641(w__1053 ,w__1118);
  not g__642(w__1052 ,w__1050);
  not g__644(w__1050 ,w__1150);
  not g__669(w__1025 ,w__1023);
  not g__671(w__1023 ,w__1129);
  not g__711(w__983 ,w__982);
  not g__712(w__982 ,w__1149);
  not g__714(w__980 ,w__979);
  not g__715(w__979 ,w__1117);
  not g__718(w__976 ,w__975);
  not g__719(w__975 ,w__1128);
  buf g__732(w__1632 ,w__1229);
  buf g__733(w__1548 ,w__1287);
  buf g__734(w__1536 ,w__1233);
  buf g__735(w__1656 ,w__1286);
  buf g__736(w__1629 ,w__1209);
  buf g__737(w__1552 ,w__1207);
  buf g__738(w__1605 ,w__1277);
  buf g__739(w__1611 ,w__1274);
  buf g__740(w__1602 ,w__1184);
  buf g__741(w__1641 ,w__1253);
  buf g__742(w__1644 ,w__1166);
  buf g__743(w__1560 ,w__1335);
  buf g__744(w__1614 ,w__1193);
  buf g__745(w__1659 ,w__1291);
  buf g__746(w__1588 ,w__1295);
  buf g__747(w__1638 ,w__1254);
  buf g__748(w__1572 ,w__1213);
  buf g__749(w__1599 ,w__1370);
  buf g__750(w__1568 ,w__1218);
  buf g__751(w__1620 ,w__1226);
  buf g__752(w__1674 ,w__1330);
  buf g__753(w__1584 ,w__1173);
  buf g__754(w__1671 ,w__1320);
  buf g__755(w__1626 ,w__1354);
  buf g__756(w__1617 ,w__1272);
  buf g__757(w__1556 ,w__1352);
  buf g__758(w__1595 ,w__1182);
  buf g__759(w__1662 ,w__1345);
  buf g__760(w__1635 ,w__1259);
  buf g__761(w__1532 ,w__1199);
  buf g__762(w__1680 ,w__1365);
  buf g__763(w__1580 ,w__1312);
  buf g__764(w__1650 ,w__1223);
  buf g__765(w__1576 ,w__1311);
  buf g__766(w__1540 ,w__1252);
  buf g__767(w__1647 ,w__1249);
  buf g__768(w__1544 ,w__1240);
  buf g__769(w__1665 ,w__1241);
  buf g__770(w__1668 ,w__1347);
  buf g__771(w__1608 ,w__1221);
  buf g__772(w__1564 ,w__1301);
  buf g__773(w__1623 ,w__1361);
  buf g__774(w__1653 ,w__1372);
  buf g__775(w__1537 ,w__1234);
  buf g__776(w__1573 ,w__1219);
  buf g__777(w__1669 ,w__1304);
  buf g__778(w__1654 ,w__1245);
  buf g__779(w__1545 ,w__1239);
  buf g__780(w__1651 ,w__1248);
  buf g__781(w__1618 ,w__1191);
  buf g__782(w__1606 ,w__1280);
  buf g__783(w__1541 ,w__1235);
  buf g__784(w__1603 ,w__1201);
  buf g__785(w__1639 ,w__1250);
  buf g__786(w__1577 ,w__1215);
  buf g__787(w__1663 ,w__1358);
  buf g__788(w__1612 ,w__1190);
  buf g__789(w__1533 ,w__1263);
  buf g__790(w__1633 ,w__1208);
  buf g__791(w__1657 ,w__1296);
  buf g__792(w__1672 ,w__1317);
  buf g__793(w__1681 ,w__1339);
  buf g__794(w__1553 ,w__1297);
  buf g__795(w__1589 ,w__1294);
  buf g__796(w__1561 ,w__1318);
  buf g__797(w__1642 ,w__1165);
  buf g__798(w__1660 ,w__1284);
  buf g__799(w__1557 ,w__1302);
  buf g__800(w__1621 ,w__1194);
  buf g__801(w__1549 ,w__1242);
  buf g__802(w__1645 ,w__1251);
  buf g__803(w__1600 ,w__1283);
  buf g__804(w__1630 ,w__1353);
  buf g__805(w__1581 ,w__1307);
  buf g__806(w__1666 ,w__1340);
  buf g__807(w__1609 ,w__1367);
  buf g__808(w__1627 ,w__1266);
  buf g__809(w__1648 ,w__1288);
  buf g__810(w__1675 ,w__1331);
  buf g__811(w__1624 ,w__1363);
  buf g__812(w__1569 ,w__1224);
  buf g__813(w__1615 ,w__1375);
  buf g__814(w__1585 ,w__1175);
  buf g__815(w__1565 ,w__1334);
  buf g__816(w__1596 ,w__1278);
  buf g__817(w__1636 ,w__1258);
  not g__926(w__857 ,w__855);
  not g__928(w__855 ,w__1144);
  not g__938(w__845 ,w__843);
  not g__940(w__843 ,w__1160);
  not g__950(w__833 ,w__831);
  not g__952(w__831 ,w__1155);
  not g__953(w__830 ,w__828);
  not g__955(w__828 ,w__1134);
  not g__962(w__821 ,w__819);
  not g__964(w__819 ,w__1123);
  not g__977(w__806 ,w__804);
  not g__979(w__804 ,w__1139);
  not g__1010(w__779 ,w__778);
  not g__1011(w__778 ,w__845);
  not g__1026(w__763 ,w__762);
  not g__1027(w__762 ,w__806);
  not g__1030(w__759 ,w__758);
  not g__1031(w__758 ,w__833);
  not g__1034(w__755 ,w__754);
  not g__1035(w__754 ,w__821);
  not g__1038(w__751 ,w__750);
  not g__1039(w__750 ,w__830);
  not g__1042(w__747 ,w__746);
  not g__1043(w__746 ,w__857);
  xnor g__1046(w__1686 ,w__23 ,in5[4]);
  and g__1047(w__1687 ,in5[4] ,w__24);
  nor g__1048(w__26 ,w__24 ,w__25);
  nor g__1049(w__25 ,in5[3] ,w__21);
  not g__1050(w__24 ,w__23);
  or g__1051(w__23 ,w__9 ,w__22);
  not g__1052(w__22 ,w__21);
  or g__1053(w__21 ,w__14 ,w__20);
  xnor g__1054(w__1684 ,w__19 ,w__16);
  and g__1055(w__20 ,w__15 ,w__19);
  xor g__1056(w__1683 ,w__13 ,w__17);
  or g__1057(w__19 ,w__10 ,w__18);
  nor g__1058(w__18 ,w__13 ,w__12);
  and g__1059(w__1682 ,w__13 ,w__11);
  xnor g__1060(w__17 ,w__1149 ,in5[1]);
  xnor g__1061(w__16 ,w__1117 ,in5[2]);
  or g__1062(w__15 ,w__1117 ,in5[2]);
  and g__1063(w__14 ,w__1117 ,in5[2]);
  or g__1064(w__13 ,w__1124 ,w__7);
  nor g__1065(w__12 ,w__1149 ,in5[1]);
  or g__1066(w__11 ,w__1688 ,in5[0]);
  and g__1067(w__10 ,w__1149 ,in5[1]);
  not g__1068(w__9 ,in5[3]);
  not g__1070(w__7 ,in5[0]);
  buf g__1077(w__1685 ,w__26);
  xnor g__1078(out1[6] ,w__1678 ,w__42);
  nor g__1079(w__42 ,w__33 ,w__41);
  xnor g__1080(out1[5] ,w__40 ,w__38);
  and g__1081(w__41 ,w__34 ,w__40);
  xor g__1082(out1[4] ,w__31 ,w__37);
  or g__1083(w__40 ,w__32 ,w__39);
  nor g__1084(w__39 ,w__31 ,w__35);
  and g__1085(out1[3] ,w__31 ,w__36);
  xnor g__1086(w__38 ,w__91 ,w__1681);
  xnor g__1087(w__37 ,w__28 ,w__1680);
  or g__1088(w__36 ,w__1679 ,in8[0]);
  nor g__1089(w__35 ,w__1680 ,w__28);
  or g__1090(w__34 ,w__1681 ,w__91);
  and g__1091(w__33 ,w__1681 ,w__91);
  and g__1092(w__32 ,w__1680 ,w__28);
  or g__1093(w__31 ,w__30 ,w__29);
  not g__1094(w__30 ,w__1679);
  not g__1095(w__29 ,in8[0]);
  buf g__1096(w__28 ,w__1527);
  xnor g__1098(out2[6] ,w__1678 ,w__58);
  nor g__1099(w__58 ,w__49 ,w__57);
  xnor g__1100(out2[5] ,w__56 ,w__54);
  and g__1101(w__57 ,w__50 ,w__56);
  xor g__1102(out2[4] ,w__47 ,w__53);
  or g__1103(w__56 ,w__48 ,w__55);
  nor g__1104(w__55 ,w__47 ,w__51);
  and g__1105(out2[3] ,w__47 ,w__52);
  xnor g__1106(w__54 ,w__91 ,w__1675);
  xnor g__1107(w__53 ,w__28 ,w__1674);
  or g__1108(w__52 ,w__1673 ,in8[0]);
  nor g__1109(w__51 ,w__1674 ,w__28);
  or g__1110(w__50 ,w__1675 ,w__91);
  and g__1111(w__49 ,w__1675 ,w__91);
  and g__1112(w__48 ,w__1674 ,w__28);
  or g__1113(w__47 ,w__46 ,w__29);
  not g__1114(w__46 ,w__1673);
  xnor g__1118(out3[6] ,w__1678 ,w__74);
  nor g__1119(w__74 ,w__65 ,w__73);
  xnor g__1120(out3[5] ,w__72 ,w__70);
  and g__1121(w__73 ,w__66 ,w__72);
  xor g__1122(out3[4] ,w__63 ,w__69);
  or g__1123(w__72 ,w__64 ,w__71);
  nor g__1124(w__71 ,w__63 ,w__67);
  and g__1125(out3[3] ,w__63 ,w__68);
  xnor g__1126(w__70 ,w__91 ,w__1672);
  xnor g__1127(w__69 ,w__60 ,w__1671);
  or g__1128(w__68 ,w__1670 ,in8[0]);
  nor g__1129(w__67 ,w__1671 ,w__60);
  or g__1130(w__66 ,w__1672 ,w__91);
  and g__1131(w__65 ,w__1672 ,w__91);
  and g__1132(w__64 ,w__1671 ,w__60);
  or g__1133(w__63 ,w__62 ,w__29);
  not g__1134(w__62 ,w__1670);
  buf g__1136(w__60 ,w__1525);
  xnor g__1138(out4[6] ,w__1678 ,w__90);
  nor g__1139(w__90 ,w__81 ,w__89);
  xnor g__1140(out4[5] ,w__88 ,w__86);
  and g__1141(w__89 ,w__82 ,w__88);
  xor g__1142(out4[4] ,w__79 ,w__85);
  or g__1143(w__88 ,w__80 ,w__87);
  nor g__1144(w__87 ,w__79 ,w__83);
  and g__1145(out4[3] ,w__79 ,w__84);
  xnor g__1146(w__86 ,w__75 ,w__1669);
  xnor g__1147(w__85 ,w__28 ,w__1668);
  or g__1148(w__84 ,w__1667 ,in8[0]);
  nor g__1149(w__83 ,w__1668 ,w__28);
  or g__1150(w__82 ,w__1669 ,w__75);
  and g__1151(w__81 ,w__1669 ,w__75);
  and g__1152(w__80 ,w__1668 ,w__28);
  or g__1153(w__79 ,w__78 ,w__29);
  not g__1154(w__78 ,w__1667);
  buf g__1157(w__75 ,w__1518);
  xnor g__1158(out5[6] ,w__1678 ,w__106);
  nor g__1159(w__106 ,w__97 ,w__105);
  xnor g__1160(out5[5] ,w__104 ,w__102);
  and g__1161(w__105 ,w__98 ,w__104);
  xor g__1162(out5[4] ,w__95 ,w__101);
  or g__1163(w__104 ,w__96 ,w__103);
  nor g__1164(w__103 ,w__95 ,w__99);
  and g__1165(out5[3] ,w__95 ,w__100);
  xnor g__1166(w__102 ,w__91 ,w__1666);
  xnor g__1167(w__101 ,w__28 ,w__1665);
  or g__1168(w__100 ,w__1664 ,in8[0]);
  nor g__1169(w__99 ,w__1665 ,w__28);
  or g__1170(w__98 ,w__1666 ,w__91);
  and g__1171(w__97 ,w__1666 ,w__91);
  and g__1172(w__96 ,w__1665 ,w__28);
  or g__1173(w__95 ,w__94 ,w__29);
  not g__1174(w__94 ,w__1664);
  buf g__1177(w__91 ,w__1530);
  xnor g__1178(out6[6] ,w__1678 ,w__122);
  nor g__1179(w__122 ,w__113 ,w__121);
  xnor g__1180(out6[5] ,w__120 ,w__118);
  and g__1181(w__121 ,w__114 ,w__120);
  xor g__1182(out6[4] ,w__111 ,w__117);
  or g__1183(w__120 ,w__112 ,w__119);
  nor g__1184(w__119 ,w__111 ,w__115);
  and g__1185(out6[3] ,w__111 ,w__116);
  xnor g__1186(w__118 ,w__91 ,w__1663);
  xnor g__1187(w__117 ,w__28 ,w__1662);
  or g__1188(w__116 ,w__1661 ,in8[0]);
  nor g__1189(w__115 ,w__1662 ,w__28);
  or g__1190(w__114 ,w__1663 ,w__91);
  and g__1191(w__113 ,w__1663 ,w__91);
  and g__1192(w__112 ,w__1662 ,w__28);
  or g__1193(w__111 ,w__110 ,w__29);
  not g__1194(w__110 ,w__1661);
  xnor g__1198(out7[6] ,w__1678 ,w__138);
  nor g__1199(w__138 ,w__129 ,w__137);
  xnor g__1200(out7[5] ,w__136 ,w__134);
  and g__1201(w__137 ,w__130 ,w__136);
  xor g__1202(out7[4] ,w__127 ,w__133);
  or g__1203(w__136 ,w__128 ,w__135);
  nor g__1204(w__135 ,w__127 ,w__131);
  and g__1205(out7[3] ,w__127 ,w__132);
  xnor g__1206(w__134 ,w__91 ,w__1660);
  xnor g__1207(w__133 ,w__28 ,w__1659);
  or g__1208(w__132 ,w__1658 ,in8[0]);
  nor g__1209(w__131 ,w__1659 ,w__28);
  or g__1210(w__130 ,w__1660 ,w__91);
  and g__1211(w__129 ,w__1660 ,w__91);
  and g__1212(w__128 ,w__1659 ,w__28);
  or g__1213(w__127 ,w__126 ,w__29);
  not g__1214(w__126 ,w__1658);
  xnor g__1218(out8[6] ,w__1678 ,w__154);
  nor g__1219(w__154 ,w__145 ,w__153);
  xnor g__1220(out8[5] ,w__152 ,w__150);
  and g__1221(w__153 ,w__146 ,w__152);
  xor g__1222(out8[4] ,w__143 ,w__149);
  or g__1223(w__152 ,w__144 ,w__151);
  nor g__1224(w__151 ,w__143 ,w__147);
  and g__1225(out8[3] ,w__143 ,w__148);
  xnor g__1226(w__150 ,w__91 ,w__1657);
  xnor g__1227(w__149 ,w__140 ,w__1656);
  or g__1228(w__148 ,w__1655 ,in8[0]);
  nor g__1229(w__147 ,w__1656 ,w__140);
  or g__1230(w__146 ,w__1657 ,w__91);
  and g__1231(w__145 ,w__1657 ,w__91);
  and g__1232(w__144 ,w__1656 ,w__140);
  or g__1233(w__143 ,w__142 ,w__29);
  not g__1234(w__142 ,w__1655);
  buf g__1236(w__140 ,w__1525);
  xnor g__1238(out9[6] ,w__1678 ,w__170);
  nor g__1239(w__170 ,w__161 ,w__169);
  xnor g__1240(out9[5] ,w__168 ,w__166);
  and g__1241(w__169 ,w__162 ,w__168);
  xor g__1242(out9[4] ,w__159 ,w__165);
  or g__1243(w__168 ,w__160 ,w__167);
  nor g__1244(w__167 ,w__159 ,w__163);
  and g__1245(out9[3] ,w__159 ,w__164);
  xnor g__1246(w__166 ,w__155 ,w__1654);
  xnor g__1247(w__165 ,w__156 ,w__1653);
  or g__1248(w__164 ,w__1652 ,in8[0]);
  nor g__1249(w__163 ,w__1653 ,w__156);
  or g__1250(w__162 ,w__1654 ,w__155);
  and g__1251(w__161 ,w__1654 ,w__155);
  and g__1252(w__160 ,w__1653 ,w__156);
  or g__1253(w__159 ,w__158 ,w__29);
  not g__1254(w__158 ,w__1652);
  buf g__1256(w__156 ,w__1519);
  buf g__1257(w__155 ,w__1520);
  xnor g__1258(out10[6] ,w__1678 ,w__186);
  nor g__1259(w__186 ,w__177 ,w__185);
  xnor g__1260(out10[5] ,w__184 ,w__182);
  and g__1261(w__185 ,w__178 ,w__184);
  xor g__1262(out10[4] ,w__175 ,w__181);
  or g__1263(w__184 ,w__176 ,w__183);
  nor g__1264(w__183 ,w__175 ,w__179);
  and g__1265(out10[3] ,w__175 ,w__180);
  xnor g__1266(w__182 ,w__91 ,w__1651);
  xnor g__1267(w__181 ,w__172 ,w__1650);
  or g__1268(w__180 ,w__1649 ,in8[0]);
  nor g__1269(w__179 ,w__1650 ,w__172);
  or g__1270(w__178 ,w__1651 ,w__91);
  and g__1271(w__177 ,w__1651 ,w__91);
  and g__1272(w__176 ,w__1650 ,w__172);
  or g__1273(w__175 ,w__174 ,w__29);
  not g__1274(w__174 ,w__1649);
  buf g__1276(w__172 ,w__1525);
  xnor g__1278(out11[6] ,w__1678 ,w__202);
  nor g__1279(w__202 ,w__193 ,w__201);
  xnor g__1280(out11[5] ,w__200 ,w__198);
  and g__1281(w__201 ,w__194 ,w__200);
  xor g__1282(out11[4] ,w__191 ,w__197);
  or g__1283(w__200 ,w__192 ,w__199);
  nor g__1284(w__199 ,w__191 ,w__195);
  and g__1285(out11[3] ,w__191 ,w__196);
  xnor g__1286(w__198 ,w__187 ,w__1648);
  xnor g__1287(w__197 ,w__28 ,w__1647);
  or g__1288(w__196 ,w__1646 ,in8[0]);
  nor g__1289(w__195 ,w__1647 ,w__28);
  or g__1290(w__194 ,w__1648 ,w__187);
  and g__1291(w__193 ,w__1648 ,w__187);
  and g__1292(w__192 ,w__1647 ,w__28);
  or g__1293(w__191 ,w__190 ,w__29);
  not g__1294(w__190 ,w__1646);
  buf g__1297(w__187 ,w__1530);
  xnor g__1298(out12[6] ,w__1678 ,w__218);
  nor g__1299(w__218 ,w__209 ,w__217);
  xnor g__1300(out12[5] ,w__216 ,w__214);
  and g__1301(w__217 ,w__210 ,w__216);
  xor g__1302(out12[4] ,w__207 ,w__213);
  or g__1303(w__216 ,w__208 ,w__215);
  nor g__1304(w__215 ,w__207 ,w__211);
  and g__1305(out12[3] ,w__207 ,w__212);
  xnor g__1306(w__214 ,w__91 ,w__1645);
  xnor g__1307(w__213 ,w__28 ,w__1644);
  or g__1308(w__212 ,w__1643 ,in8[0]);
  nor g__1309(w__211 ,w__1644 ,w__28);
  or g__1310(w__210 ,w__1645 ,w__91);
  and g__1311(w__209 ,w__1645 ,w__91);
  and g__1312(w__208 ,w__1644 ,w__28);
  or g__1313(w__207 ,w__206 ,w__29);
  not g__1314(w__206 ,w__1643);
  xnor g__1318(out13[6] ,w__1678 ,w__234);
  nor g__1319(w__234 ,w__225 ,w__233);
  xnor g__1320(out13[5] ,w__232 ,w__230);
  and g__1321(w__233 ,w__226 ,w__232);
  xor g__1322(out13[4] ,w__223 ,w__229);
  or g__1323(w__232 ,w__224 ,w__231);
  nor g__1324(w__231 ,w__223 ,w__227);
  and g__1325(out13[3] ,w__223 ,w__228);
  xnor g__1326(w__230 ,w__219 ,w__1642);
  xnor g__1327(w__229 ,w__220 ,w__1641);
  or g__1328(w__228 ,w__1640 ,in8[0]);
  nor g__1329(w__227 ,w__1641 ,w__220);
  or g__1330(w__226 ,w__1642 ,w__219);
  and g__1331(w__225 ,w__1642 ,w__219);
  and g__1332(w__224 ,w__1641 ,w__220);
  or g__1333(w__223 ,w__222 ,w__29);
  not g__1334(w__222 ,w__1640);
  buf g__1336(w__220 ,w__1523);
  buf g__1337(w__219 ,w__1524);
  xnor g__1338(out14[6] ,w__1678 ,w__250);
  nor g__1339(w__250 ,w__241 ,w__249);
  xnor g__1340(out14[5] ,w__248 ,w__246);
  and g__1341(w__249 ,w__242 ,w__248);
  xor g__1342(out14[4] ,w__239 ,w__245);
  or g__1343(w__248 ,w__240 ,w__247);
  nor g__1344(w__247 ,w__239 ,w__243);
  and g__1345(out14[3] ,w__239 ,w__244);
  xnor g__1346(w__246 ,w__235 ,w__1639);
  xnor g__1347(w__245 ,w__236 ,w__1638);
  or g__1348(w__244 ,w__1637 ,in8[0]);
  nor g__1349(w__243 ,w__1638 ,w__236);
  or g__1350(w__242 ,w__1639 ,w__235);
  and g__1351(w__241 ,w__1639 ,w__235);
  and g__1352(w__240 ,w__1638 ,w__236);
  or g__1353(w__239 ,w__238 ,w__29);
  not g__1354(w__238 ,w__1637);
  buf g__1356(w__236 ,w__1523);
  buf g__1357(w__235 ,w__1524);
  xnor g__1358(out15[6] ,w__1678 ,w__266);
  nor g__1359(w__266 ,w__257 ,w__265);
  xnor g__1360(out15[5] ,w__264 ,w__262);
  and g__1361(w__265 ,w__258 ,w__264);
  xor g__1362(out15[4] ,w__255 ,w__261);
  or g__1363(w__264 ,w__256 ,w__263);
  nor g__1364(w__263 ,w__255 ,w__259);
  and g__1365(out15[3] ,w__255 ,w__260);
  xnor g__1366(w__262 ,w__91 ,w__1636);
  xnor g__1367(w__261 ,w__28 ,w__1635);
  or g__1368(w__260 ,w__1634 ,in8[0]);
  nor g__1369(w__259 ,w__1635 ,w__28);
  or g__1370(w__258 ,w__1636 ,w__91);
  and g__1371(w__257 ,w__1636 ,w__91);
  and g__1372(w__256 ,w__1635 ,w__28);
  or g__1373(w__255 ,w__254 ,w__29);
  not g__1374(w__254 ,w__1634);
  xnor g__1378(out16[6] ,w__1678 ,w__282);
  nor g__1379(w__282 ,w__273 ,w__281);
  xnor g__1380(out16[5] ,w__280 ,w__278);
  and g__1381(w__281 ,w__274 ,w__280);
  xor g__1382(out16[4] ,w__271 ,w__277);
  or g__1383(w__280 ,w__272 ,w__279);
  nor g__1384(w__279 ,w__271 ,w__275);
  and g__1385(out16[3] ,w__271 ,w__276);
  xnor g__1386(w__278 ,w__91 ,w__1633);
  xnor g__1387(w__277 ,w__28 ,w__1632);
  or g__1388(w__276 ,w__1631 ,in8[0]);
  nor g__1389(w__275 ,w__1632 ,w__28);
  or g__1390(w__274 ,w__1633 ,w__91);
  and g__1391(w__273 ,w__1633 ,w__91);
  and g__1392(w__272 ,w__1632 ,w__28);
  or g__1393(w__271 ,w__270 ,w__29);
  not g__1394(w__270 ,w__1631);
  xnor g__1398(out17[6] ,w__1678 ,w__298);
  nor g__1399(w__298 ,w__289 ,w__297);
  xnor g__1400(out17[5] ,w__296 ,w__294);
  and g__1401(w__297 ,w__290 ,w__296);
  xor g__1402(out17[4] ,w__287 ,w__293);
  or g__1403(w__296 ,w__288 ,w__295);
  nor g__1404(w__295 ,w__287 ,w__291);
  and g__1405(out17[3] ,w__287 ,w__292);
  xnor g__1406(w__294 ,w__283 ,w__1630);
  xnor g__1407(w__293 ,w__284 ,w__1629);
  or g__1408(w__292 ,w__1628 ,in8[0]);
  nor g__1409(w__291 ,w__1629 ,w__284);
  or g__1410(w__290 ,w__1630 ,w__283);
  and g__1411(w__289 ,w__1630 ,w__283);
  and g__1412(w__288 ,w__1629 ,w__284);
  or g__1413(w__287 ,w__286 ,w__29);
  not g__1414(w__286 ,w__1628);
  buf g__1416(w__284 ,w__1519);
  buf g__1417(w__283 ,w__1520);
  xnor g__1418(out18[6] ,w__1678 ,w__314);
  nor g__1419(w__314 ,w__305 ,w__313);
  xnor g__1420(out18[5] ,w__312 ,w__310);
  and g__1421(w__313 ,w__306 ,w__312);
  xor g__1422(out18[4] ,w__303 ,w__309);
  or g__1423(w__312 ,w__304 ,w__311);
  nor g__1424(w__311 ,w__303 ,w__307);
  and g__1425(out18[3] ,w__303 ,w__308);
  xnor g__1426(w__310 ,w__299 ,w__1627);
  xnor g__1427(w__309 ,w__300 ,w__1626);
  or g__1428(w__308 ,w__1625 ,in8[0]);
  nor g__1429(w__307 ,w__1626 ,w__300);
  or g__1430(w__306 ,w__1627 ,w__299);
  and g__1431(w__305 ,w__1627 ,w__299);
  and g__1432(w__304 ,w__1626 ,w__300);
  or g__1433(w__303 ,w__302 ,w__29);
  not g__1434(w__302 ,w__1625);
  buf g__1436(w__300 ,w__1519);
  buf g__1437(w__299 ,w__1520);
  xnor g__1438(out19[6] ,w__1678 ,w__330);
  nor g__1439(w__330 ,w__321 ,w__329);
  xnor g__1440(out19[5] ,w__328 ,w__326);
  and g__1441(w__329 ,w__322 ,w__328);
  xor g__1442(out19[4] ,w__319 ,w__325);
  or g__1443(w__328 ,w__320 ,w__327);
  nor g__1444(w__327 ,w__319 ,w__323);
  and g__1445(out19[3] ,w__319 ,w__324);
  xnor g__1446(w__326 ,w__91 ,w__1624);
  xnor g__1447(w__325 ,w__316 ,w__1623);
  or g__1448(w__324 ,w__1622 ,in8[0]);
  nor g__1449(w__323 ,w__1623 ,w__316);
  or g__1450(w__322 ,w__1624 ,w__91);
  and g__1451(w__321 ,w__1624 ,w__91);
  and g__1452(w__320 ,w__1623 ,w__316);
  or g__1453(w__319 ,w__318 ,w__29);
  not g__1454(w__318 ,w__1622);
  buf g__1456(w__316 ,w__1527);
  xnor g__1458(out20[6] ,w__1678 ,w__346);
  nor g__1459(w__346 ,w__337 ,w__345);
  xnor g__1460(out20[5] ,w__344 ,w__342);
  and g__1461(w__345 ,w__338 ,w__344);
  xor g__1462(out20[4] ,w__335 ,w__341);
  or g__1463(w__344 ,w__336 ,w__343);
  nor g__1464(w__343 ,w__335 ,w__339);
  and g__1465(out20[3] ,w__335 ,w__340);
  xnor g__1466(w__342 ,w__331 ,w__1621);
  xnor g__1467(w__341 ,w__28 ,w__1620);
  or g__1468(w__340 ,w__1619 ,in8[0]);
  nor g__1469(w__339 ,w__1620 ,w__28);
  or g__1470(w__338 ,w__1621 ,w__331);
  and g__1471(w__337 ,w__1621 ,w__331);
  and g__1472(w__336 ,w__1620 ,w__28);
  or g__1473(w__335 ,w__334 ,w__29);
  not g__1474(w__334 ,w__1619);
  buf g__1477(w__331 ,w__1518);
  xnor g__1478(out21[6] ,w__1678 ,w__362);
  nor g__1479(w__362 ,w__353 ,w__361);
  xnor g__1480(out21[5] ,w__360 ,w__358);
  and g__1481(w__361 ,w__354 ,w__360);
  xor g__1482(out21[4] ,w__351 ,w__357);
  or g__1483(w__360 ,w__352 ,w__359);
  nor g__1484(w__359 ,w__351 ,w__355);
  and g__1485(out21[3] ,w__351 ,w__356);
  xnor g__1486(w__358 ,w__347 ,w__1618);
  xnor g__1487(w__357 ,w__348 ,w__1617);
  or g__1488(w__356 ,w__1616 ,in8[0]);
  nor g__1489(w__355 ,w__1617 ,w__348);
  or g__1490(w__354 ,w__1618 ,w__347);
  and g__1491(w__353 ,w__1618 ,w__347);
  and g__1492(w__352 ,w__1617 ,w__348);
  or g__1493(w__351 ,w__350 ,w__29);
  not g__1494(w__350 ,w__1616);
  buf g__1496(w__348 ,w__1523);
  buf g__1497(w__347 ,w__1524);
  xnor g__1498(out22[6] ,w__1678 ,w__378);
  nor g__1499(w__378 ,w__369 ,w__377);
  xnor g__1500(out22[5] ,w__376 ,w__374);
  and g__1501(w__377 ,w__370 ,w__376);
  xor g__1502(out22[4] ,w__367 ,w__373);
  or g__1503(w__376 ,w__368 ,w__375);
  nor g__1504(w__375 ,w__367 ,w__371);
  and g__1505(out22[3] ,w__367 ,w__372);
  xnor g__1506(w__374 ,w__363 ,w__1615);
  xnor g__1507(w__373 ,w__28 ,w__1614);
  or g__1508(w__372 ,w__1613 ,in8[0]);
  nor g__1509(w__371 ,w__1614 ,w__28);
  or g__1510(w__370 ,w__1615 ,w__363);
  and g__1511(w__369 ,w__1615 ,w__363);
  and g__1512(w__368 ,w__1614 ,w__28);
  or g__1513(w__367 ,w__366 ,w__29);
  not g__1514(w__366 ,w__1613);
  buf g__1517(w__363 ,w__1518);
  xnor g__1518(out23[6] ,w__1678 ,w__394);
  nor g__1519(w__394 ,w__385 ,w__393);
  xnor g__1520(out23[5] ,w__392 ,w__390);
  and g__1521(w__393 ,w__386 ,w__392);
  xor g__1522(out23[4] ,w__383 ,w__389);
  or g__1523(w__392 ,w__384 ,w__391);
  nor g__1524(w__391 ,w__383 ,w__387);
  and g__1525(out23[3] ,w__383 ,w__388);
  xnor g__1526(w__390 ,w__379 ,w__1612);
  xnor g__1527(w__389 ,w__380 ,w__1611);
  or g__1528(w__388 ,w__1610 ,in8[0]);
  nor g__1529(w__387 ,w__1611 ,w__380);
  or g__1530(w__386 ,w__1612 ,w__379);
  and g__1531(w__385 ,w__1612 ,w__379);
  and g__1532(w__384 ,w__1611 ,w__380);
  or g__1533(w__383 ,w__382 ,w__29);
  not g__1534(w__382 ,w__1610);
  buf g__1536(w__380 ,w__1519);
  buf g__1537(w__379 ,w__1520);
  xnor g__1538(out24[6] ,w__1678 ,w__410);
  nor g__1539(w__410 ,w__401 ,w__409);
  xnor g__1540(out24[5] ,w__408 ,w__406);
  and g__1541(w__409 ,w__402 ,w__408);
  xor g__1542(out24[4] ,w__399 ,w__405);
  or g__1543(w__408 ,w__400 ,w__407);
  nor g__1544(w__407 ,w__399 ,w__403);
  and g__1545(out24[3] ,w__399 ,w__404);
  xnor g__1546(w__406 ,w__91 ,w__1609);
  xnor g__1547(w__405 ,w__396 ,w__1608);
  or g__1548(w__404 ,w__1607 ,in8[0]);
  nor g__1549(w__403 ,w__1608 ,w__396);
  or g__1550(w__402 ,w__1609 ,w__91);
  and g__1551(w__401 ,w__1609 ,w__91);
  and g__1552(w__400 ,w__1608 ,w__396);
  or g__1553(w__399 ,w__398 ,w__29);
  not g__1554(w__398 ,w__1607);
  buf g__1556(w__396 ,w__1525);
  xnor g__1558(out25[6] ,w__1678 ,w__426);
  nor g__1559(w__426 ,w__417 ,w__425);
  xnor g__1560(out25[5] ,w__424 ,w__422);
  and g__1561(w__425 ,w__418 ,w__424);
  xor g__1562(out25[4] ,w__415 ,w__421);
  or g__1563(w__424 ,w__416 ,w__423);
  nor g__1564(w__423 ,w__415 ,w__419);
  and g__1565(out25[3] ,w__415 ,w__420);
  xnor g__1566(w__422 ,w__411 ,w__1606);
  xnor g__1567(w__421 ,w__28 ,w__1605);
  or g__1568(w__420 ,w__1604 ,in8[0]);
  nor g__1569(w__419 ,w__1605 ,w__28);
  or g__1570(w__418 ,w__1606 ,w__411);
  and g__1571(w__417 ,w__1606 ,w__411);
  and g__1572(w__416 ,w__1605 ,w__28);
  or g__1573(w__415 ,w__414 ,w__29);
  not g__1574(w__414 ,w__1604);
  buf g__1577(w__411 ,w__1518);
  xnor g__1578(out26[6] ,w__1678 ,w__442);
  nor g__1579(w__442 ,w__433 ,w__441);
  xnor g__1580(out26[5] ,w__440 ,w__438);
  and g__1581(w__441 ,w__434 ,w__440);
  xor g__1582(out26[4] ,w__431 ,w__437);
  or g__1583(w__440 ,w__432 ,w__439);
  nor g__1584(w__439 ,w__431 ,w__435);
  and g__1585(out26[3] ,w__431 ,w__436);
  xnor g__1586(w__438 ,w__91 ,w__1603);
  xnor g__1587(w__437 ,w__28 ,w__1602);
  or g__1588(w__436 ,w__1601 ,in8[0]);
  nor g__1589(w__435 ,w__1602 ,w__28);
  or g__1590(w__434 ,w__1603 ,w__91);
  and g__1591(w__433 ,w__1603 ,w__91);
  and g__1592(w__432 ,w__1602 ,w__28);
  or g__1593(w__431 ,w__430 ,w__29);
  not g__1594(w__430 ,w__1601);
  xnor g__1598(out27[6] ,w__1678 ,w__458);
  nor g__1599(w__458 ,w__449 ,w__457);
  xnor g__1600(out27[5] ,w__456 ,w__454);
  and g__1601(w__457 ,w__450 ,w__456);
  xor g__1602(out27[4] ,w__447 ,w__453);
  or g__1603(w__456 ,w__448 ,w__455);
  nor g__1604(w__455 ,w__447 ,w__451);
  and g__1605(out27[3] ,w__447 ,w__452);
  xnor g__1606(w__454 ,w__91 ,w__1600);
  xnor g__1607(w__453 ,w__28 ,w__1599);
  or g__1608(w__452 ,w__1598 ,in8[0]);
  nor g__1609(w__451 ,w__1599 ,w__28);
  or g__1610(w__450 ,w__1600 ,w__91);
  and g__1611(w__449 ,w__1600 ,w__91);
  and g__1612(w__448 ,w__1599 ,w__28);
  or g__1613(w__447 ,w__446 ,w__29);
  not g__1614(w__446 ,w__1598);
  xnor g__1618(out28[5] ,w__470 ,w__475);
  or g__1619(w__475 ,w__466 ,w__474);
  xnor g__1620(out28[4] ,w__473 ,w__469);
  and g__1621(w__474 ,w__468 ,w__473);
  xor g__1622(out28[3] ,w__463 ,w__471);
  or g__1623(w__473 ,w__467 ,w__472);
  nor g__1624(w__472 ,w__463 ,w__465);
  and g__1625(out28[2] ,w__463 ,w__464);
  xnor g__1626(w__471 ,w__477 ,w__1595);
  xnor g__1627(w__470 ,w__1593 ,w__1597);
  xnor g__1628(w__469 ,w__459 ,w__1596);
  or g__1629(w__468 ,w__1596 ,w__459);
  and g__1630(w__467 ,w__1595 ,w__477);
  and g__1631(w__466 ,w__1596 ,w__459);
  nor g__1632(w__465 ,w__1595 ,w__477);
  or g__1633(w__464 ,w__1594 ,in8[0]);
  or g__1634(w__463 ,w__462 ,w__29);
  not g__1635(w__462 ,w__1594);
  buf g__1638(w__459 ,w__1516);
  xnor g__1639(out29[5] ,w__487 ,w__492);
  or g__1640(w__492 ,w__483 ,w__491);
  xnor g__1641(out29[4] ,w__490 ,w__486);
  and g__1642(w__491 ,w__485 ,w__490);
  xor g__1643(out29[3] ,w__480 ,w__488);
  or g__1644(w__490 ,w__484 ,w__489);
  nor g__1645(w__489 ,w__480 ,w__482);
  and g__1646(out29[2] ,w__480 ,w__481);
  xnor g__1647(w__488 ,w__477 ,w__1588);
  xnor g__1648(w__487 ,w__1593 ,w__1590);
  xnor g__1649(w__486 ,w__459 ,w__1589);
  or g__1650(w__485 ,w__1589 ,w__459);
  and g__1651(w__484 ,w__1588 ,w__477);
  and g__1652(w__483 ,w__1589 ,w__459);
  nor g__1653(w__482 ,w__1588 ,w__477);
  or g__1654(w__481 ,w__1587 ,in8[0]);
  or g__1655(w__480 ,w__479 ,w__29);
  not g__1656(w__479 ,w__1587);
  buf g__1658(w__477 ,w__1509);
  xnor g__1660(out30[5] ,w__504 ,w__509);
  or g__1661(w__509 ,w__500 ,w__508);
  xnor g__1662(out30[4] ,w__507 ,w__503);
  and g__1663(w__508 ,w__502 ,w__507);
  xor g__1664(out30[3] ,w__497 ,w__505);
  or g__1665(w__507 ,w__501 ,w__506);
  nor g__1666(w__506 ,w__497 ,w__499);
  and g__1667(out30[2] ,w__497 ,w__498);
  xnor g__1668(w__505 ,w__494 ,w__1584);
  xnor g__1669(w__504 ,w__1593 ,w__1586);
  xnor g__1670(w__503 ,w__493 ,w__1585);
  or g__1671(w__502 ,w__1585 ,w__493);
  and g__1672(w__501 ,w__1584 ,w__494);
  and g__1673(w__500 ,w__1585 ,w__493);
  nor g__1674(w__499 ,w__1584 ,w__494);
  or g__1675(w__498 ,w__1583 ,in8[0]);
  or g__1676(w__497 ,w__496 ,w__29);
  not g__1677(w__496 ,w__1583);
  buf g__1679(w__494 ,w__1513);
  buf g__1680(w__493 ,w__1514);
  xnor g__1681(out31[5] ,w__521 ,w__526);
  or g__1682(w__526 ,w__517 ,w__525);
  xnor g__1683(out31[4] ,w__524 ,w__520);
  and g__1684(w__525 ,w__519 ,w__524);
  xor g__1685(out31[3] ,w__514 ,w__522);
  or g__1686(w__524 ,w__518 ,w__523);
  nor g__1687(w__523 ,w__514 ,w__516);
  and g__1688(out31[2] ,w__514 ,w__515);
  xnor g__1689(w__522 ,w__477 ,w__1580);
  xnor g__1690(w__521 ,w__1593 ,w__1582);
  xnor g__1691(w__520 ,w__459 ,w__1581);
  or g__1692(w__519 ,w__1581 ,w__459);
  and g__1693(w__518 ,w__1580 ,w__477);
  and g__1694(w__517 ,w__1581 ,w__459);
  nor g__1695(w__516 ,w__1580 ,w__477);
  or g__1696(w__515 ,w__1579 ,in8[0]);
  or g__1697(w__514 ,w__513 ,w__29);
  not g__1698(w__513 ,w__1579);
  xnor g__1702(out32[5] ,w__538 ,w__543);
  or g__1703(w__543 ,w__534 ,w__542);
  xnor g__1704(out32[4] ,w__541 ,w__537);
  and g__1705(w__542 ,w__536 ,w__541);
  xor g__1706(out32[3] ,w__531 ,w__539);
  or g__1707(w__541 ,w__535 ,w__540);
  nor g__1708(w__540 ,w__531 ,w__533);
  and g__1709(out32[2] ,w__531 ,w__532);
  xnor g__1710(w__539 ,w__477 ,w__1576);
  xnor g__1711(w__538 ,w__1593 ,w__1578);
  xnor g__1712(w__537 ,w__459 ,w__1577);
  or g__1713(w__536 ,w__1577 ,w__459);
  and g__1714(w__535 ,w__1576 ,w__477);
  and g__1715(w__534 ,w__1577 ,w__459);
  nor g__1716(w__533 ,w__1576 ,w__477);
  or g__1717(w__532 ,w__1575 ,in8[0]);
  or g__1718(w__531 ,w__530 ,w__29);
  not g__1719(w__530 ,w__1575);
  xnor g__1723(out33[5] ,w__555 ,w__560);
  or g__1724(w__560 ,w__551 ,w__559);
  xnor g__1725(out33[4] ,w__558 ,w__554);
  and g__1726(w__559 ,w__553 ,w__558);
  xor g__1727(out33[3] ,w__548 ,w__556);
  or g__1728(w__558 ,w__552 ,w__557);
  nor g__1729(w__557 ,w__548 ,w__550);
  and g__1730(out33[2] ,w__548 ,w__549);
  xnor g__1731(w__556 ,w__545 ,w__1572);
  xnor g__1732(w__555 ,w__1593 ,w__1574);
  xnor g__1733(w__554 ,w__544 ,w__1573);
  or g__1734(w__553 ,w__1573 ,w__544);
  and g__1735(w__552 ,w__1572 ,w__545);
  and g__1736(w__551 ,w__1573 ,w__544);
  nor g__1737(w__550 ,w__1572 ,w__545);
  or g__1738(w__549 ,w__1571 ,in8[0]);
  or g__1739(w__548 ,w__547 ,w__29);
  not g__1740(w__547 ,w__1571);
  buf g__1742(w__545 ,w__1513);
  buf g__1743(w__544 ,w__1514);
  xnor g__1744(out34[5] ,w__572 ,w__577);
  or g__1745(w__577 ,w__568 ,w__576);
  xnor g__1746(out34[4] ,w__575 ,w__571);
  and g__1747(w__576 ,w__570 ,w__575);
  xor g__1748(out34[3] ,w__565 ,w__573);
  or g__1749(w__575 ,w__569 ,w__574);
  nor g__1750(w__574 ,w__565 ,w__567);
  and g__1751(out34[2] ,w__565 ,w__566);
  xnor g__1752(w__573 ,w__477 ,w__1568);
  xnor g__1753(w__572 ,w__1593 ,w__1570);
  xnor g__1754(w__571 ,w__459 ,w__1569);
  or g__1755(w__570 ,w__1569 ,w__459);
  and g__1756(w__569 ,w__1568 ,w__477);
  and g__1757(w__568 ,w__1569 ,w__459);
  nor g__1758(w__567 ,w__1568 ,w__477);
  or g__1759(w__566 ,w__1567 ,in8[0]);
  or g__1760(w__565 ,w__564 ,w__29);
  not g__1761(w__564 ,w__1567);
  xnor g__1765(out35[5] ,w__589 ,w__594);
  or g__1766(w__594 ,w__585 ,w__593);
  xnor g__1767(out35[4] ,w__592 ,w__588);
  and g__1768(w__593 ,w__587 ,w__592);
  xor g__1769(out35[3] ,w__582 ,w__590);
  or g__1770(w__592 ,w__586 ,w__591);
  nor g__1771(w__591 ,w__582 ,w__584);
  and g__1772(out35[2] ,w__582 ,w__583);
  xnor g__1773(w__590 ,w__477 ,w__1564);
  xnor g__1774(w__589 ,w__1593 ,w__1566);
  xnor g__1775(w__588 ,w__459 ,w__1565);
  or g__1776(w__587 ,w__1565 ,w__459);
  and g__1777(w__586 ,w__1564 ,w__477);
  and g__1778(w__585 ,w__1565 ,w__459);
  nor g__1779(w__584 ,w__1564 ,w__477);
  or g__1780(w__583 ,w__1563 ,in8[0]);
  or g__1781(w__582 ,w__581 ,w__29);
  not g__1782(w__581 ,w__1563);
  xnor g__1786(out36[5] ,w__606 ,w__611);
  or g__1787(w__611 ,w__602 ,w__610);
  xnor g__1788(out36[4] ,w__609 ,w__605);
  and g__1789(w__610 ,w__604 ,w__609);
  xor g__1790(out36[3] ,w__599 ,w__607);
  or g__1791(w__609 ,w__603 ,w__608);
  nor g__1792(w__608 ,w__599 ,w__601);
  and g__1793(out36[2] ,w__599 ,w__600);
  xnor g__1794(w__607 ,w__477 ,w__1560);
  xnor g__1795(w__606 ,w__1593 ,w__1562);
  xnor g__1796(w__605 ,w__595 ,w__1561);
  or g__1797(w__604 ,w__1561 ,w__595);
  and g__1798(w__603 ,w__1560 ,w__477);
  and g__1799(w__602 ,w__1561 ,w__595);
  nor g__1800(w__601 ,w__1560 ,w__477);
  or g__1801(w__600 ,w__1559 ,in8[0]);
  or g__1802(w__599 ,w__598 ,w__29);
  not g__1803(w__598 ,w__1559);
  buf g__1806(w__595 ,w__1516);
  xnor g__1807(out37[5] ,w__623 ,w__628);
  or g__1808(w__628 ,w__619 ,w__627);
  xnor g__1809(out37[4] ,w__626 ,w__622);
  and g__1810(w__627 ,w__621 ,w__626);
  xor g__1811(out37[3] ,w__616 ,w__624);
  or g__1812(w__626 ,w__620 ,w__625);
  nor g__1813(w__625 ,w__616 ,w__618);
  and g__1814(out37[2] ,w__616 ,w__617);
  xnor g__1815(w__624 ,w__477 ,w__1556);
  xnor g__1816(w__623 ,w__1593 ,w__1558);
  xnor g__1817(w__622 ,w__459 ,w__1557);
  or g__1818(w__621 ,w__1557 ,w__459);
  and g__1819(w__620 ,w__1556 ,w__477);
  and g__1820(w__619 ,w__1557 ,w__459);
  nor g__1821(w__618 ,w__1556 ,w__477);
  or g__1822(w__617 ,w__1555 ,in8[0]);
  or g__1823(w__616 ,w__615 ,w__29);
  not g__1824(w__615 ,w__1555);
  xnor g__1828(out38[5] ,w__640 ,w__645);
  or g__1829(w__645 ,w__636 ,w__644);
  xnor g__1830(out38[4] ,w__643 ,w__639);
  and g__1831(w__644 ,w__638 ,w__643);
  xor g__1832(out38[3] ,w__633 ,w__641);
  or g__1833(w__643 ,w__637 ,w__642);
  nor g__1834(w__642 ,w__633 ,w__635);
  and g__1835(out38[2] ,w__633 ,w__634);
  xnor g__1836(w__641 ,w__630 ,w__1552);
  xnor g__1837(w__640 ,w__1593 ,w__1554);
  xnor g__1838(w__639 ,w__459 ,w__1553);
  or g__1839(w__638 ,w__1553 ,w__459);
  and g__1840(w__637 ,w__1552 ,w__630);
  and g__1841(w__636 ,w__1553 ,w__459);
  nor g__1842(w__635 ,w__1552 ,w__630);
  or g__1843(w__634 ,w__1551 ,in8[0]);
  or g__1844(w__633 ,w__632 ,w__29);
  not g__1845(w__632 ,w__1551);
  buf g__1847(w__630 ,w__1509);
  xnor g__1849(out39[5] ,w__657 ,w__662);
  or g__1850(w__662 ,w__653 ,w__661);
  xnor g__1851(out39[4] ,w__660 ,w__656);
  and g__1852(w__661 ,w__655 ,w__660);
  xor g__1853(out39[3] ,w__650 ,w__658);
  or g__1854(w__660 ,w__654 ,w__659);
  nor g__1855(w__659 ,w__650 ,w__652);
  and g__1856(out39[2] ,w__650 ,w__651);
  xnor g__1857(w__658 ,w__647 ,w__1548);
  xnor g__1858(w__657 ,w__1593 ,w__1550);
  xnor g__1859(w__656 ,w__646 ,w__1549);
  or g__1860(w__655 ,w__1549 ,w__646);
  and g__1861(w__654 ,w__1548 ,w__647);
  and g__1862(w__653 ,w__1549 ,w__646);
  nor g__1863(w__652 ,w__1548 ,w__647);
  or g__1864(w__651 ,w__1547 ,in8[0]);
  or g__1865(w__650 ,w__649 ,w__29);
  not g__1866(w__649 ,w__1547);
  buf g__1868(w__647 ,w__1513);
  buf g__1869(w__646 ,w__1514);
  xnor g__1870(out40[5] ,w__674 ,w__679);
  or g__1871(w__679 ,w__670 ,w__678);
  xnor g__1872(out40[4] ,w__677 ,w__673);
  and g__1873(w__678 ,w__672 ,w__677);
  xor g__1874(out40[3] ,w__667 ,w__675);
  or g__1875(w__677 ,w__671 ,w__676);
  nor g__1876(w__676 ,w__667 ,w__669);
  and g__1877(out40[2] ,w__667 ,w__668);
  xnor g__1878(w__675 ,w__664 ,w__1544);
  xnor g__1879(w__674 ,w__1593 ,w__1546);
  xnor g__1880(w__673 ,w__663 ,w__1545);
  or g__1881(w__672 ,w__1545 ,w__663);
  and g__1882(w__671 ,w__1544 ,w__664);
  and g__1883(w__670 ,w__1545 ,w__663);
  nor g__1884(w__669 ,w__1544 ,w__664);
  or g__1885(w__668 ,w__1543 ,in8[0]);
  or g__1886(w__667 ,w__666 ,w__29);
  not g__1887(w__666 ,w__1543);
  buf g__1889(w__664 ,w__1513);
  buf g__1890(w__663 ,w__1514);
  xnor g__1891(out41[5] ,w__691 ,w__696);
  or g__1892(w__696 ,w__687 ,w__695);
  xnor g__1893(out41[4] ,w__694 ,w__690);
  and g__1894(w__695 ,w__689 ,w__694);
  xor g__1895(out41[3] ,w__684 ,w__692);
  or g__1896(w__694 ,w__688 ,w__693);
  nor g__1897(w__693 ,w__684 ,w__686);
  and g__1898(out41[2] ,w__684 ,w__685);
  xnor g__1899(w__692 ,w__477 ,w__1540);
  xnor g__1900(w__691 ,w__1593 ,w__1542);
  xnor g__1901(w__690 ,w__459 ,w__1541);
  or g__1902(w__689 ,w__1541 ,w__459);
  and g__1903(w__688 ,w__1540 ,w__477);
  and g__1904(w__687 ,w__1541 ,w__459);
  nor g__1905(w__686 ,w__1540 ,w__477);
  or g__1906(w__685 ,w__1539 ,in8[0]);
  or g__1907(w__684 ,w__683 ,w__29);
  not g__1908(w__683 ,w__1539);
  xnor g__1912(out42[5] ,w__708 ,w__713);
  or g__1913(w__713 ,w__704 ,w__712);
  xnor g__1914(out42[4] ,w__711 ,w__707);
  and g__1915(w__712 ,w__706 ,w__711);
  xor g__1916(out42[3] ,w__701 ,w__709);
  or g__1917(w__711 ,w__705 ,w__710);
  nor g__1918(w__710 ,w__701 ,w__703);
  and g__1919(out42[2] ,w__701 ,w__702);
  xnor g__1920(w__709 ,w__477 ,w__1536);
  xnor g__1921(w__708 ,w__1593 ,w__1538);
  xnor g__1922(w__707 ,w__459 ,w__1537);
  or g__1923(w__706 ,w__1537 ,w__459);
  and g__1924(w__705 ,w__1536 ,w__477);
  and g__1925(w__704 ,w__1537 ,w__459);
  nor g__1926(w__703 ,w__1536 ,w__477);
  or g__1927(w__702 ,w__1535 ,in8[0]);
  or g__1928(w__701 ,w__700 ,w__29);
  not g__1929(w__700 ,w__1535);
  xnor g__1933(out43[5] ,w__725 ,w__730);
  or g__1934(w__730 ,w__721 ,w__729);
  xnor g__1935(out43[4] ,w__728 ,w__724);
  and g__1936(w__729 ,w__723 ,w__728);
  xor g__1937(out43[3] ,w__718 ,w__726);
  or g__1938(w__728 ,w__722 ,w__727);
  nor g__1939(w__727 ,w__718 ,w__720);
  and g__1940(out43[2] ,w__718 ,w__719);
  xnor g__1941(w__726 ,w__477 ,w__1532);
  xnor g__1942(w__725 ,w__1593 ,w__1534);
  xnor g__1943(w__724 ,w__459 ,w__1533);
  or g__1944(w__723 ,w__1533 ,w__459);
  and g__1945(w__722 ,w__1532 ,w__477);
  and g__1946(w__721 ,w__1533 ,w__459);
  nor g__1947(w__720 ,w__1532 ,w__477);
  or g__1948(w__719 ,w__1531 ,in8[0]);
  or g__1949(w__718 ,w__717 ,w__29);
  not g__1950(w__717 ,w__1531);
  xnor g__1954(w__1677 ,w__733 ,in8[1]);
  not g__1955(w__736 ,w__735);
  and g__1956(w__1676 ,w__733 ,w__734);
  or g__1957(w__734 ,in8[1] ,in8[0]);
  or g__1958(w__733 ,w__732 ,w__29);
  not g__1959(w__732 ,in8[1]);
  buf g__1961(w__1678 ,w__736);
  xnor g__1962(w__1592 ,w__739 ,in8[1]);
  and g__1963(w__743 ,in8[1] ,w__740);
  nor g__1964(w__742 ,w__740 ,w__741);
  nor g__1965(w__741 ,in8[1] ,in8[0]);
  not g__1966(w__740 ,w__739);
  or g__1967(w__739 ,w__732 ,w__29);
  buf g__1970(w__1593 ,w__743);
  buf g__1971(w__1591 ,w__742);
  xnor g__1972(w__1689 ,inc_add_183_20_n_4 ,in2[1]);
  and g__1973(w__1690 ,in2[1] ,inc_add_183_20_n_3);
  and g__1974(inc_add_183_20_n_6 ,inc_add_183_20_n_4 ,inc_add_183_20_n_5);
  or g__1975(inc_add_183_20_n_5 ,in2[0] ,in1);
  not g__1976(inc_add_183_20_n_3 ,inc_add_183_20_n_4);
  or g__1977(inc_add_183_20_n_4 ,inc_add_183_20_n_1 ,inc_add_183_20_n_2);
  not g__1978(inc_add_183_20_n_2 ,in1);
  not g__1979(inc_add_183_20_n_1 ,in2[0]);
  buf g__1980(w__1688 ,inc_add_183_20_n_6);
  buf g__1981(w__735 ,w__733);

endmodule

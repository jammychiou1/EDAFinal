module top(in1, in2, in3, in4, in5, in6, out1, out2, out3, out4, out5);
  input [1:0] in1;
  input [1:0] in2;
  input [4:0] in3;
  input [2:0] in4;
  input [4:0] in5;
  input [2:0] in6;
  output [4:0] out1;
  output out2;
  output [4:0] out3;
  output out4;
  output [4:0] out5;
  wire [1:0] in1;
  wire [1:0] in2;
  wire [4:0] in3;
  wire [2:0] in4;
  wire [4:0] in5;
  wire [2:0] in6;
  wire [4:0] out1;
  wire out2;
  wire [4:0] out3;
  wire out4;
  wire [4:0] out5;
  assign out1 = 1 + in2 - 5 * in1 - 4 * in1 * in1 + 8 * in1 * in1 * in1;

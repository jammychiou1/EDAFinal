module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, out1);

  input [10:0] in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24;

  output [25:0] out1;
  wire [10:0] in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24;
  wire [25:0] out1;
  wire csa_tree_add_51_79_groupi_n_0, csa_tree_add_51_79_groupi_n_1, csa_tree_add_51_79_groupi_n_2, csa_tree_add_51_79_groupi_n_3, csa_tree_add_51_79_groupi_n_4, csa_tree_add_51_79_groupi_n_5, csa_tree_add_51_79_groupi_n_6, csa_tree_add_51_79_groupi_n_7;
  wire csa_tree_add_51_79_groupi_n_8, csa_tree_add_51_79_groupi_n_9, csa_tree_add_51_79_groupi_n_10, csa_tree_add_51_79_groupi_n_11, csa_tree_add_51_79_groupi_n_12, csa_tree_add_51_79_groupi_n_13, csa_tree_add_51_79_groupi_n_14, csa_tree_add_51_79_groupi_n_15;
  wire csa_tree_add_51_79_groupi_n_16, csa_tree_add_51_79_groupi_n_17, csa_tree_add_51_79_groupi_n_18, csa_tree_add_51_79_groupi_n_19, csa_tree_add_51_79_groupi_n_20, csa_tree_add_51_79_groupi_n_21, csa_tree_add_51_79_groupi_n_22, csa_tree_add_51_79_groupi_n_23;
  wire csa_tree_add_51_79_groupi_n_24, csa_tree_add_51_79_groupi_n_25, csa_tree_add_51_79_groupi_n_26, csa_tree_add_51_79_groupi_n_27, csa_tree_add_51_79_groupi_n_28, csa_tree_add_51_79_groupi_n_29, csa_tree_add_51_79_groupi_n_30, csa_tree_add_51_79_groupi_n_31;
  wire csa_tree_add_51_79_groupi_n_32, csa_tree_add_51_79_groupi_n_33, csa_tree_add_51_79_groupi_n_34, csa_tree_add_51_79_groupi_n_35, csa_tree_add_51_79_groupi_n_36, csa_tree_add_51_79_groupi_n_37, csa_tree_add_51_79_groupi_n_38, csa_tree_add_51_79_groupi_n_39;
  wire csa_tree_add_51_79_groupi_n_40, csa_tree_add_51_79_groupi_n_41, csa_tree_add_51_79_groupi_n_42, csa_tree_add_51_79_groupi_n_43, csa_tree_add_51_79_groupi_n_44, csa_tree_add_51_79_groupi_n_45, csa_tree_add_51_79_groupi_n_46, csa_tree_add_51_79_groupi_n_47;
  wire csa_tree_add_51_79_groupi_n_48, csa_tree_add_51_79_groupi_n_49, csa_tree_add_51_79_groupi_n_1036, csa_tree_add_51_79_groupi_n_1038, csa_tree_add_51_79_groupi_n_1038, csa_tree_add_51_79_groupi_n_53, csa_tree_add_51_79_groupi_n_54, csa_tree_add_51_79_groupi_n_55;
  wire csa_tree_add_51_79_groupi_n_1024, csa_tree_add_51_79_groupi_n_1026, csa_tree_add_51_79_groupi_n_1026, csa_tree_add_51_79_groupi_n_59, csa_tree_add_51_79_groupi_n_60, csa_tree_add_51_79_groupi_n_61, csa_tree_add_51_79_groupi_n_1018, csa_tree_add_51_79_groupi_n_1020;
  wire csa_tree_add_51_79_groupi_n_1020, csa_tree_add_51_79_groupi_n_65, csa_tree_add_51_79_groupi_n_66, csa_tree_add_51_79_groupi_n_67, csa_tree_add_51_79_groupi_n_1015, csa_tree_add_51_79_groupi_n_1017, csa_tree_add_51_79_groupi_n_1017, csa_tree_add_51_79_groupi_n_71;
  wire csa_tree_add_51_79_groupi_n_72, csa_tree_add_51_79_groupi_n_73, csa_tree_add_51_79_groupi_n_1009, csa_tree_add_51_79_groupi_n_1011, csa_tree_add_51_79_groupi_n_1011, csa_tree_add_51_79_groupi_n_77, csa_tree_add_51_79_groupi_n_78, csa_tree_add_51_79_groupi_n_79;
  wire csa_tree_add_51_79_groupi_n_1006, csa_tree_add_51_79_groupi_n_1008, csa_tree_add_51_79_groupi_n_1008, csa_tree_add_51_79_groupi_n_83, csa_tree_add_51_79_groupi_n_84, csa_tree_add_51_79_groupi_n_85, csa_tree_add_51_79_groupi_n_1063, csa_tree_add_51_79_groupi_n_1065;
  wire csa_tree_add_51_79_groupi_n_1065, csa_tree_add_51_79_groupi_n_89, csa_tree_add_51_79_groupi_n_90, csa_tree_add_51_79_groupi_n_91, csa_tree_add_51_79_groupi_n_1003, csa_tree_add_51_79_groupi_n_1005, csa_tree_add_51_79_groupi_n_1005, csa_tree_add_51_79_groupi_n_95;
  wire csa_tree_add_51_79_groupi_n_96, csa_tree_add_51_79_groupi_n_97, csa_tree_add_51_79_groupi_n_1000, csa_tree_add_51_79_groupi_n_1002, csa_tree_add_51_79_groupi_n_1002, csa_tree_add_51_79_groupi_n_101, csa_tree_add_51_79_groupi_n_102, csa_tree_add_51_79_groupi_n_103;
  wire csa_tree_add_51_79_groupi_n_1060, csa_tree_add_51_79_groupi_n_1062, csa_tree_add_51_79_groupi_n_1062, csa_tree_add_51_79_groupi_n_107, csa_tree_add_51_79_groupi_n_108, csa_tree_add_51_79_groupi_n_109, csa_tree_add_51_79_groupi_n_1057, csa_tree_add_51_79_groupi_n_1059;
  wire csa_tree_add_51_79_groupi_n_1059, csa_tree_add_51_79_groupi_n_113, csa_tree_add_51_79_groupi_n_114, csa_tree_add_51_79_groupi_n_115, csa_tree_add_51_79_groupi_n_997, csa_tree_add_51_79_groupi_n_999, csa_tree_add_51_79_groupi_n_999, csa_tree_add_51_79_groupi_n_119;
  wire csa_tree_add_51_79_groupi_n_120, csa_tree_add_51_79_groupi_n_121, csa_tree_add_51_79_groupi_n_991, csa_tree_add_51_79_groupi_n_993, csa_tree_add_51_79_groupi_n_993, csa_tree_add_51_79_groupi_n_125, csa_tree_add_51_79_groupi_n_126, csa_tree_add_51_79_groupi_n_127;
  wire csa_tree_add_51_79_groupi_n_994, csa_tree_add_51_79_groupi_n_996, csa_tree_add_51_79_groupi_n_996, csa_tree_add_51_79_groupi_n_131, csa_tree_add_51_79_groupi_n_132, csa_tree_add_51_79_groupi_n_133, csa_tree_add_51_79_groupi_n_982, csa_tree_add_51_79_groupi_n_984;
  wire csa_tree_add_51_79_groupi_n_984, csa_tree_add_51_79_groupi_n_137, csa_tree_add_51_79_groupi_n_138, csa_tree_add_51_79_groupi_n_139, csa_tree_add_51_79_groupi_n_988, csa_tree_add_51_79_groupi_n_990, csa_tree_add_51_79_groupi_n_990, csa_tree_add_51_79_groupi_n_143;
  wire csa_tree_add_51_79_groupi_n_144, csa_tree_add_51_79_groupi_n_145, csa_tree_add_51_79_groupi_n_985, csa_tree_add_51_79_groupi_n_987, csa_tree_add_51_79_groupi_n_987, csa_tree_add_51_79_groupi_n_149, csa_tree_add_51_79_groupi_n_150, csa_tree_add_51_79_groupi_n_151;
  wire csa_tree_add_51_79_groupi_n_1054, csa_tree_add_51_79_groupi_n_1056, csa_tree_add_51_79_groupi_n_1056, csa_tree_add_51_79_groupi_n_155, csa_tree_add_51_79_groupi_n_156, csa_tree_add_51_79_groupi_n_157, csa_tree_add_51_79_groupi_n_1051, csa_tree_add_51_79_groupi_n_1053;
  wire csa_tree_add_51_79_groupi_n_1053, csa_tree_add_51_79_groupi_n_161, csa_tree_add_51_79_groupi_n_162, csa_tree_add_51_79_groupi_n_163, csa_tree_add_51_79_groupi_n_973, csa_tree_add_51_79_groupi_n_975, csa_tree_add_51_79_groupi_n_975, csa_tree_add_51_79_groupi_n_167;
  wire csa_tree_add_51_79_groupi_n_168, csa_tree_add_51_79_groupi_n_169, csa_tree_add_51_79_groupi_n_979, csa_tree_add_51_79_groupi_n_981, csa_tree_add_51_79_groupi_n_981, csa_tree_add_51_79_groupi_n_173, csa_tree_add_51_79_groupi_n_174, csa_tree_add_51_79_groupi_n_175;
  wire csa_tree_add_51_79_groupi_n_976, csa_tree_add_51_79_groupi_n_978, csa_tree_add_51_79_groupi_n_978, csa_tree_add_51_79_groupi_n_179, csa_tree_add_51_79_groupi_n_180, csa_tree_add_51_79_groupi_n_181, csa_tree_add_51_79_groupi_n_964, csa_tree_add_51_79_groupi_n_966;
  wire csa_tree_add_51_79_groupi_n_966, csa_tree_add_51_79_groupi_n_185, csa_tree_add_51_79_groupi_n_186, csa_tree_add_51_79_groupi_n_187, csa_tree_add_51_79_groupi_n_970, csa_tree_add_51_79_groupi_n_972, csa_tree_add_51_79_groupi_n_972, csa_tree_add_51_79_groupi_n_191;
  wire csa_tree_add_51_79_groupi_n_192, csa_tree_add_51_79_groupi_n_193, csa_tree_add_51_79_groupi_n_967, csa_tree_add_51_79_groupi_n_969, csa_tree_add_51_79_groupi_n_969, csa_tree_add_51_79_groupi_n_197, csa_tree_add_51_79_groupi_n_198, csa_tree_add_51_79_groupi_n_199;
  wire csa_tree_add_51_79_groupi_n_1045, csa_tree_add_51_79_groupi_n_1047, csa_tree_add_51_79_groupi_n_1047, csa_tree_add_51_79_groupi_n_203, csa_tree_add_51_79_groupi_n_204, csa_tree_add_51_79_groupi_n_205, csa_tree_add_51_79_groupi_n_955, csa_tree_add_51_79_groupi_n_957;
  wire csa_tree_add_51_79_groupi_n_957, csa_tree_add_51_79_groupi_n_209, csa_tree_add_51_79_groupi_n_210, csa_tree_add_51_79_groupi_n_211, csa_tree_add_51_79_groupi_n_961, csa_tree_add_51_79_groupi_n_963, csa_tree_add_51_79_groupi_n_963, csa_tree_add_51_79_groupi_n_215;
  wire csa_tree_add_51_79_groupi_n_216, csa_tree_add_51_79_groupi_n_217, csa_tree_add_51_79_groupi_n_958, csa_tree_add_51_79_groupi_n_960, csa_tree_add_51_79_groupi_n_960, csa_tree_add_51_79_groupi_n_221, csa_tree_add_51_79_groupi_n_222, csa_tree_add_51_79_groupi_n_223;
  wire csa_tree_add_51_79_groupi_n_946, csa_tree_add_51_79_groupi_n_948, csa_tree_add_51_79_groupi_n_948, csa_tree_add_51_79_groupi_n_227, csa_tree_add_51_79_groupi_n_228, csa_tree_add_51_79_groupi_n_229, csa_tree_add_51_79_groupi_n_952, csa_tree_add_51_79_groupi_n_954;
  wire csa_tree_add_51_79_groupi_n_954, csa_tree_add_51_79_groupi_n_233, csa_tree_add_51_79_groupi_n_234, csa_tree_add_51_79_groupi_n_235, csa_tree_add_51_79_groupi_n_949, csa_tree_add_51_79_groupi_n_951, csa_tree_add_51_79_groupi_n_951, csa_tree_add_51_79_groupi_n_239;
  wire csa_tree_add_51_79_groupi_n_240, csa_tree_add_51_79_groupi_n_241, csa_tree_add_51_79_groupi_n_1048, csa_tree_add_51_79_groupi_n_1050, csa_tree_add_51_79_groupi_n_1050, csa_tree_add_51_79_groupi_n_245, csa_tree_add_51_79_groupi_n_246, csa_tree_add_51_79_groupi_n_247;
  wire csa_tree_add_51_79_groupi_n_1042, csa_tree_add_51_79_groupi_n_1044, csa_tree_add_51_79_groupi_n_1044, csa_tree_add_51_79_groupi_n_251, csa_tree_add_51_79_groupi_n_252, csa_tree_add_51_79_groupi_n_253, csa_tree_add_51_79_groupi_n_1039, csa_tree_add_51_79_groupi_n_1041;
  wire csa_tree_add_51_79_groupi_n_1041, csa_tree_add_51_79_groupi_n_257, csa_tree_add_51_79_groupi_n_258, csa_tree_add_51_79_groupi_n_259, csa_tree_add_51_79_groupi_n_937, csa_tree_add_51_79_groupi_n_939, csa_tree_add_51_79_groupi_n_939, csa_tree_add_51_79_groupi_n_263;
  wire csa_tree_add_51_79_groupi_n_264, csa_tree_add_51_79_groupi_n_265, csa_tree_add_51_79_groupi_n_943, csa_tree_add_51_79_groupi_n_945, csa_tree_add_51_79_groupi_n_945, csa_tree_add_51_79_groupi_n_269, csa_tree_add_51_79_groupi_n_270, csa_tree_add_51_79_groupi_n_271;
  wire csa_tree_add_51_79_groupi_n_940, csa_tree_add_51_79_groupi_n_942, csa_tree_add_51_79_groupi_n_942, csa_tree_add_51_79_groupi_n_275, csa_tree_add_51_79_groupi_n_276, csa_tree_add_51_79_groupi_n_277, csa_tree_add_51_79_groupi_n_928, csa_tree_add_51_79_groupi_n_930;
  wire csa_tree_add_51_79_groupi_n_930, csa_tree_add_51_79_groupi_n_281, csa_tree_add_51_79_groupi_n_282, csa_tree_add_51_79_groupi_n_283, csa_tree_add_51_79_groupi_n_934, csa_tree_add_51_79_groupi_n_936, csa_tree_add_51_79_groupi_n_936, csa_tree_add_51_79_groupi_n_287;
  wire csa_tree_add_51_79_groupi_n_288, csa_tree_add_51_79_groupi_n_289, csa_tree_add_51_79_groupi_n_931, csa_tree_add_51_79_groupi_n_933, csa_tree_add_51_79_groupi_n_933, csa_tree_add_51_79_groupi_n_293, csa_tree_add_51_79_groupi_n_294, csa_tree_add_51_79_groupi_n_295;
  wire csa_tree_add_51_79_groupi_n_1033, csa_tree_add_51_79_groupi_n_1035, csa_tree_add_51_79_groupi_n_1035, csa_tree_add_51_79_groupi_n_299, csa_tree_add_51_79_groupi_n_300, csa_tree_add_51_79_groupi_n_301, csa_tree_add_51_79_groupi_n_919, csa_tree_add_51_79_groupi_n_921;
  wire csa_tree_add_51_79_groupi_n_921, csa_tree_add_51_79_groupi_n_305, csa_tree_add_51_79_groupi_n_306, csa_tree_add_51_79_groupi_n_307, csa_tree_add_51_79_groupi_n_925, csa_tree_add_51_79_groupi_n_927, csa_tree_add_51_79_groupi_n_927, csa_tree_add_51_79_groupi_n_311;
  wire csa_tree_add_51_79_groupi_n_312, csa_tree_add_51_79_groupi_n_313, csa_tree_add_51_79_groupi_n_922, csa_tree_add_51_79_groupi_n_924, csa_tree_add_51_79_groupi_n_924, csa_tree_add_51_79_groupi_n_317, csa_tree_add_51_79_groupi_n_318, csa_tree_add_51_79_groupi_n_319;
  wire csa_tree_add_51_79_groupi_n_910, csa_tree_add_51_79_groupi_n_912, csa_tree_add_51_79_groupi_n_912, csa_tree_add_51_79_groupi_n_323, csa_tree_add_51_79_groupi_n_324, csa_tree_add_51_79_groupi_n_325, csa_tree_add_51_79_groupi_n_916, csa_tree_add_51_79_groupi_n_918;
  wire csa_tree_add_51_79_groupi_n_918, csa_tree_add_51_79_groupi_n_329, csa_tree_add_51_79_groupi_n_330, csa_tree_add_51_79_groupi_n_331, csa_tree_add_51_79_groupi_n_913, csa_tree_add_51_79_groupi_n_915, csa_tree_add_51_79_groupi_n_915, csa_tree_add_51_79_groupi_n_335;
  wire csa_tree_add_51_79_groupi_n_336, csa_tree_add_51_79_groupi_n_337, csa_tree_add_51_79_groupi_n_1030, csa_tree_add_51_79_groupi_n_1032, csa_tree_add_51_79_groupi_n_1032, csa_tree_add_51_79_groupi_n_341, csa_tree_add_51_79_groupi_n_342, csa_tree_add_51_79_groupi_n_343;
  wire csa_tree_add_51_79_groupi_n_1027, csa_tree_add_51_79_groupi_n_1029, csa_tree_add_51_79_groupi_n_1029, csa_tree_add_51_79_groupi_n_347, csa_tree_add_51_79_groupi_n_348, csa_tree_add_51_79_groupi_n_349, csa_tree_add_51_79_groupi_n_901, csa_tree_add_51_79_groupi_n_903;
  wire csa_tree_add_51_79_groupi_n_903, csa_tree_add_51_79_groupi_n_353, csa_tree_add_51_79_groupi_n_354, csa_tree_add_51_79_groupi_n_355, csa_tree_add_51_79_groupi_n_907, csa_tree_add_51_79_groupi_n_909, csa_tree_add_51_79_groupi_n_909, csa_tree_add_51_79_groupi_n_359;
  wire csa_tree_add_51_79_groupi_n_360, csa_tree_add_51_79_groupi_n_361, csa_tree_add_51_79_groupi_n_904, csa_tree_add_51_79_groupi_n_906, csa_tree_add_51_79_groupi_n_906, csa_tree_add_51_79_groupi_n_365, csa_tree_add_51_79_groupi_n_366, csa_tree_add_51_79_groupi_n_367;
  wire csa_tree_add_51_79_groupi_n_895, csa_tree_add_51_79_groupi_n_897, csa_tree_add_51_79_groupi_n_897, csa_tree_add_51_79_groupi_n_371, csa_tree_add_51_79_groupi_n_372, csa_tree_add_51_79_groupi_n_373, csa_tree_add_51_79_groupi_n_898, csa_tree_add_51_79_groupi_n_900;
  wire csa_tree_add_51_79_groupi_n_900, csa_tree_add_51_79_groupi_n_377, csa_tree_add_51_79_groupi_n_378, csa_tree_add_51_79_groupi_n_379, csa_tree_add_51_79_groupi_n_892, csa_tree_add_51_79_groupi_n_894, csa_tree_add_51_79_groupi_n_894, csa_tree_add_51_79_groupi_n_383;
  wire csa_tree_add_51_79_groupi_n_384, csa_tree_add_51_79_groupi_n_385, csa_tree_add_51_79_groupi_n_1021, csa_tree_add_51_79_groupi_n_1023, csa_tree_add_51_79_groupi_n_1023, csa_tree_add_51_79_groupi_n_389, csa_tree_add_51_79_groupi_n_390, csa_tree_add_51_79_groupi_n_391;
  wire csa_tree_add_51_79_groupi_n_889, csa_tree_add_51_79_groupi_n_891, csa_tree_add_51_79_groupi_n_891, csa_tree_add_51_79_groupi_n_395, csa_tree_add_51_79_groupi_n_396, csa_tree_add_51_79_groupi_n_397, csa_tree_add_51_79_groupi_n_1012, csa_tree_add_51_79_groupi_n_1014;
  wire csa_tree_add_51_79_groupi_n_1014, csa_tree_add_51_79_groupi_n_401, csa_tree_add_51_79_groupi_n_402, csa_tree_add_51_79_groupi_n_403, csa_tree_add_51_79_groupi_n_404, csa_tree_add_51_79_groupi_n_405, csa_tree_add_51_79_groupi_n_406, csa_tree_add_51_79_groupi_n_407;
  wire csa_tree_add_51_79_groupi_n_408, csa_tree_add_51_79_groupi_n_409, csa_tree_add_51_79_groupi_n_410, csa_tree_add_51_79_groupi_n_411, csa_tree_add_51_79_groupi_n_412, csa_tree_add_51_79_groupi_n_413, csa_tree_add_51_79_groupi_n_414, csa_tree_add_51_79_groupi_n_415;
  wire csa_tree_add_51_79_groupi_n_416, csa_tree_add_51_79_groupi_n_417, csa_tree_add_51_79_groupi_n_418, csa_tree_add_51_79_groupi_n_419, csa_tree_add_51_79_groupi_n_420, csa_tree_add_51_79_groupi_n_421, csa_tree_add_51_79_groupi_n_422, csa_tree_add_51_79_groupi_n_423;
  wire csa_tree_add_51_79_groupi_n_424, csa_tree_add_51_79_groupi_n_425, csa_tree_add_51_79_groupi_n_426, csa_tree_add_51_79_groupi_n_427, csa_tree_add_51_79_groupi_n_428, csa_tree_add_51_79_groupi_n_429, csa_tree_add_51_79_groupi_n_430, csa_tree_add_51_79_groupi_n_431;
  wire csa_tree_add_51_79_groupi_n_432, csa_tree_add_51_79_groupi_n_433, csa_tree_add_51_79_groupi_n_434, csa_tree_add_51_79_groupi_n_435, csa_tree_add_51_79_groupi_n_436, csa_tree_add_51_79_groupi_n_437, csa_tree_add_51_79_groupi_n_438, csa_tree_add_51_79_groupi_n_439;
  wire csa_tree_add_51_79_groupi_n_440, csa_tree_add_51_79_groupi_n_441, csa_tree_add_51_79_groupi_n_442, csa_tree_add_51_79_groupi_n_443, csa_tree_add_51_79_groupi_n_444, csa_tree_add_51_79_groupi_n_445, csa_tree_add_51_79_groupi_n_446, csa_tree_add_51_79_groupi_n_447;
  wire csa_tree_add_51_79_groupi_n_448, csa_tree_add_51_79_groupi_n_449, csa_tree_add_51_79_groupi_n_450, csa_tree_add_51_79_groupi_n_451, csa_tree_add_51_79_groupi_n_452, csa_tree_add_51_79_groupi_n_453, csa_tree_add_51_79_groupi_n_454, csa_tree_add_51_79_groupi_n_455;
  wire csa_tree_add_51_79_groupi_n_456, csa_tree_add_51_79_groupi_n_457, csa_tree_add_51_79_groupi_n_458, csa_tree_add_51_79_groupi_n_459, csa_tree_add_51_79_groupi_n_460, csa_tree_add_51_79_groupi_n_461, csa_tree_add_51_79_groupi_n_462, csa_tree_add_51_79_groupi_n_463;
  wire csa_tree_add_51_79_groupi_n_464, csa_tree_add_51_79_groupi_n_465, csa_tree_add_51_79_groupi_n_466, csa_tree_add_51_79_groupi_n_467, csa_tree_add_51_79_groupi_n_468, csa_tree_add_51_79_groupi_n_469, csa_tree_add_51_79_groupi_n_470, csa_tree_add_51_79_groupi_n_471;
  wire csa_tree_add_51_79_groupi_n_472, csa_tree_add_51_79_groupi_n_473, csa_tree_add_51_79_groupi_n_474, csa_tree_add_51_79_groupi_n_475, csa_tree_add_51_79_groupi_n_476, csa_tree_add_51_79_groupi_n_477, csa_tree_add_51_79_groupi_n_478, csa_tree_add_51_79_groupi_n_479;
  wire csa_tree_add_51_79_groupi_n_480, csa_tree_add_51_79_groupi_n_481, csa_tree_add_51_79_groupi_n_482, csa_tree_add_51_79_groupi_n_483, csa_tree_add_51_79_groupi_n_484, csa_tree_add_51_79_groupi_n_485, csa_tree_add_51_79_groupi_n_486, csa_tree_add_51_79_groupi_n_487;
  wire csa_tree_add_51_79_groupi_n_488, csa_tree_add_51_79_groupi_n_489, csa_tree_add_51_79_groupi_n_490, csa_tree_add_51_79_groupi_n_491, csa_tree_add_51_79_groupi_n_492, csa_tree_add_51_79_groupi_n_493, csa_tree_add_51_79_groupi_n_494, csa_tree_add_51_79_groupi_n_495;
  wire csa_tree_add_51_79_groupi_n_496, csa_tree_add_51_79_groupi_n_497, csa_tree_add_51_79_groupi_n_498, csa_tree_add_51_79_groupi_n_499, csa_tree_add_51_79_groupi_n_500, csa_tree_add_51_79_groupi_n_501, csa_tree_add_51_79_groupi_n_502, csa_tree_add_51_79_groupi_n_503;
  wire csa_tree_add_51_79_groupi_n_504, csa_tree_add_51_79_groupi_n_505, csa_tree_add_51_79_groupi_n_506, csa_tree_add_51_79_groupi_n_507, csa_tree_add_51_79_groupi_n_508, csa_tree_add_51_79_groupi_n_509, csa_tree_add_51_79_groupi_n_510, csa_tree_add_51_79_groupi_n_511;
  wire csa_tree_add_51_79_groupi_n_512, csa_tree_add_51_79_groupi_n_513, csa_tree_add_51_79_groupi_n_514, csa_tree_add_51_79_groupi_n_515, csa_tree_add_51_79_groupi_n_516, csa_tree_add_51_79_groupi_n_517, csa_tree_add_51_79_groupi_n_518, csa_tree_add_51_79_groupi_n_519;
  wire csa_tree_add_51_79_groupi_n_520, csa_tree_add_51_79_groupi_n_521, csa_tree_add_51_79_groupi_n_522, csa_tree_add_51_79_groupi_n_523, csa_tree_add_51_79_groupi_n_524, csa_tree_add_51_79_groupi_n_525, csa_tree_add_51_79_groupi_n_526, csa_tree_add_51_79_groupi_n_527;
  wire csa_tree_add_51_79_groupi_n_528, csa_tree_add_51_79_groupi_n_529, csa_tree_add_51_79_groupi_n_530, csa_tree_add_51_79_groupi_n_531, csa_tree_add_51_79_groupi_n_532, csa_tree_add_51_79_groupi_n_533, csa_tree_add_51_79_groupi_n_534, csa_tree_add_51_79_groupi_n_535;
  wire csa_tree_add_51_79_groupi_n_536, csa_tree_add_51_79_groupi_n_537, csa_tree_add_51_79_groupi_n_538, csa_tree_add_51_79_groupi_n_539, csa_tree_add_51_79_groupi_n_540, csa_tree_add_51_79_groupi_n_541, csa_tree_add_51_79_groupi_n_542, csa_tree_add_51_79_groupi_n_543;
  wire csa_tree_add_51_79_groupi_n_544, csa_tree_add_51_79_groupi_n_545, csa_tree_add_51_79_groupi_n_546, csa_tree_add_51_79_groupi_n_547, csa_tree_add_51_79_groupi_n_548, csa_tree_add_51_79_groupi_n_549, csa_tree_add_51_79_groupi_n_550, csa_tree_add_51_79_groupi_n_551;
  wire csa_tree_add_51_79_groupi_n_552, csa_tree_add_51_79_groupi_n_553, csa_tree_add_51_79_groupi_n_554, csa_tree_add_51_79_groupi_n_555, csa_tree_add_51_79_groupi_n_556, csa_tree_add_51_79_groupi_n_557, csa_tree_add_51_79_groupi_n_558, csa_tree_add_51_79_groupi_n_559;
  wire csa_tree_add_51_79_groupi_n_560, csa_tree_add_51_79_groupi_n_561, csa_tree_add_51_79_groupi_n_562, csa_tree_add_51_79_groupi_n_563, csa_tree_add_51_79_groupi_n_564, csa_tree_add_51_79_groupi_n_565, csa_tree_add_51_79_groupi_n_566, csa_tree_add_51_79_groupi_n_567;
  wire csa_tree_add_51_79_groupi_n_568, csa_tree_add_51_79_groupi_n_569, csa_tree_add_51_79_groupi_n_570, csa_tree_add_51_79_groupi_n_571, csa_tree_add_51_79_groupi_n_572, csa_tree_add_51_79_groupi_n_573, csa_tree_add_51_79_groupi_n_574, csa_tree_add_51_79_groupi_n_575;
  wire csa_tree_add_51_79_groupi_n_576, csa_tree_add_51_79_groupi_n_577, csa_tree_add_51_79_groupi_n_578, csa_tree_add_51_79_groupi_n_579, csa_tree_add_51_79_groupi_n_580, csa_tree_add_51_79_groupi_n_581, csa_tree_add_51_79_groupi_n_582, csa_tree_add_51_79_groupi_n_583;
  wire csa_tree_add_51_79_groupi_n_584, csa_tree_add_51_79_groupi_n_585, csa_tree_add_51_79_groupi_n_586, csa_tree_add_51_79_groupi_n_587, csa_tree_add_51_79_groupi_n_588, csa_tree_add_51_79_groupi_n_589, csa_tree_add_51_79_groupi_n_590, csa_tree_add_51_79_groupi_n_591;
  wire csa_tree_add_51_79_groupi_n_592, csa_tree_add_51_79_groupi_n_593, csa_tree_add_51_79_groupi_n_594, csa_tree_add_51_79_groupi_n_595, csa_tree_add_51_79_groupi_n_596, csa_tree_add_51_79_groupi_n_597, csa_tree_add_51_79_groupi_n_598, csa_tree_add_51_79_groupi_n_599;
  wire csa_tree_add_51_79_groupi_n_600, csa_tree_add_51_79_groupi_n_601, csa_tree_add_51_79_groupi_n_602, csa_tree_add_51_79_groupi_n_603, csa_tree_add_51_79_groupi_n_604, csa_tree_add_51_79_groupi_n_605, csa_tree_add_51_79_groupi_n_606, csa_tree_add_51_79_groupi_n_607;
  wire csa_tree_add_51_79_groupi_n_1066, csa_tree_add_51_79_groupi_n_1068, csa_tree_add_51_79_groupi_n_1068, csa_tree_add_51_79_groupi_n_1468, csa_tree_add_51_79_groupi_n_1469, csa_tree_add_51_79_groupi_n_1469, csa_tree_add_51_79_groupi_n_1470, csa_tree_add_51_79_groupi_n_1471;
  wire csa_tree_add_51_79_groupi_n_1471, csa_tree_add_51_79_groupi_n_1466, csa_tree_add_51_79_groupi_n_1467, csa_tree_add_51_79_groupi_n_1467, csa_tree_add_51_79_groupi_n_683, csa_tree_add_51_79_groupi_n_685, csa_tree_add_51_79_groupi_n_685, csa_tree_add_51_79_groupi_n_695;
  wire csa_tree_add_51_79_groupi_n_697, csa_tree_add_51_79_groupi_n_697, csa_tree_add_51_79_groupi_n_698, csa_tree_add_51_79_groupi_n_700, csa_tree_add_51_79_groupi_n_700, csa_tree_add_51_79_groupi_n_668, csa_tree_add_51_79_groupi_n_670, csa_tree_add_51_79_groupi_n_670;
  wire csa_tree_add_51_79_groupi_n_737, csa_tree_add_51_79_groupi_n_739, csa_tree_add_51_79_groupi_n_739, csa_tree_add_51_79_groupi_n_674, csa_tree_add_51_79_groupi_n_676, csa_tree_add_51_79_groupi_n_676, csa_tree_add_51_79_groupi_n_749, csa_tree_add_51_79_groupi_n_751;
  wire csa_tree_add_51_79_groupi_n_751, csa_tree_add_51_79_groupi_n_728, csa_tree_add_51_79_groupi_n_730, csa_tree_add_51_79_groupi_n_730, csa_tree_add_51_79_groupi_n_692, csa_tree_add_51_79_groupi_n_694, csa_tree_add_51_79_groupi_n_694, csa_tree_add_51_79_groupi_n_656;
  wire csa_tree_add_51_79_groupi_n_658, csa_tree_add_51_79_groupi_n_658, csa_tree_add_51_79_groupi_n_671, csa_tree_add_51_79_groupi_n_673, csa_tree_add_51_79_groupi_n_673, csa_tree_add_51_79_groupi_n_725, csa_tree_add_51_79_groupi_n_727, csa_tree_add_51_79_groupi_n_727;
  wire csa_tree_add_51_79_groupi_n_656, csa_tree_add_51_79_groupi_n_658, csa_tree_add_51_79_groupi_n_658, csa_tree_add_51_79_groupi_n_710, csa_tree_add_51_79_groupi_n_712, csa_tree_add_51_79_groupi_n_712, csa_tree_add_51_79_groupi_n_680, csa_tree_add_51_79_groupi_n_682;
  wire csa_tree_add_51_79_groupi_n_682, csa_tree_add_51_79_groupi_n_707, csa_tree_add_51_79_groupi_n_709, csa_tree_add_51_79_groupi_n_709, csa_tree_add_51_79_groupi_n_668, csa_tree_add_51_79_groupi_n_670, csa_tree_add_51_79_groupi_n_670, csa_tree_add_51_79_groupi_n_671;
  wire csa_tree_add_51_79_groupi_n_673, csa_tree_add_51_79_groupi_n_673, csa_tree_add_51_79_groupi_n_674, csa_tree_add_51_79_groupi_n_676, csa_tree_add_51_79_groupi_n_676, csa_tree_add_51_79_groupi_n_722, csa_tree_add_51_79_groupi_n_724, csa_tree_add_51_79_groupi_n_724;
  wire csa_tree_add_51_79_groupi_n_680, csa_tree_add_51_79_groupi_n_682, csa_tree_add_51_79_groupi_n_682, csa_tree_add_51_79_groupi_n_683, csa_tree_add_51_79_groupi_n_685, csa_tree_add_51_79_groupi_n_685, csa_tree_add_51_79_groupi_n_704, csa_tree_add_51_79_groupi_n_706;
  wire csa_tree_add_51_79_groupi_n_706, csa_tree_add_51_79_groupi_n_740, csa_tree_add_51_79_groupi_n_742, csa_tree_add_51_79_groupi_n_742, csa_tree_add_51_79_groupi_n_692, csa_tree_add_51_79_groupi_n_694, csa_tree_add_51_79_groupi_n_694, csa_tree_add_51_79_groupi_n_695;
  wire csa_tree_add_51_79_groupi_n_697, csa_tree_add_51_79_groupi_n_697, csa_tree_add_51_79_groupi_n_698, csa_tree_add_51_79_groupi_n_700, csa_tree_add_51_79_groupi_n_700, csa_tree_add_51_79_groupi_n_716, csa_tree_add_51_79_groupi_n_718, csa_tree_add_51_79_groupi_n_718;
  wire csa_tree_add_51_79_groupi_n_704, csa_tree_add_51_79_groupi_n_706, csa_tree_add_51_79_groupi_n_706, csa_tree_add_51_79_groupi_n_707, csa_tree_add_51_79_groupi_n_709, csa_tree_add_51_79_groupi_n_709, csa_tree_add_51_79_groupi_n_710, csa_tree_add_51_79_groupi_n_712;
  wire csa_tree_add_51_79_groupi_n_712, csa_tree_add_51_79_groupi_n_734, csa_tree_add_51_79_groupi_n_736, csa_tree_add_51_79_groupi_n_736, csa_tree_add_51_79_groupi_n_716, csa_tree_add_51_79_groupi_n_718, csa_tree_add_51_79_groupi_n_718, csa_tree_add_51_79_groupi_n_746;
  wire csa_tree_add_51_79_groupi_n_748, csa_tree_add_51_79_groupi_n_748, csa_tree_add_51_79_groupi_n_722, csa_tree_add_51_79_groupi_n_724, csa_tree_add_51_79_groupi_n_724, csa_tree_add_51_79_groupi_n_725, csa_tree_add_51_79_groupi_n_727, csa_tree_add_51_79_groupi_n_727;
  wire csa_tree_add_51_79_groupi_n_728, csa_tree_add_51_79_groupi_n_730, csa_tree_add_51_79_groupi_n_730, csa_tree_add_51_79_groupi_n_743, csa_tree_add_51_79_groupi_n_745, csa_tree_add_51_79_groupi_n_745, csa_tree_add_51_79_groupi_n_734, csa_tree_add_51_79_groupi_n_736;
  wire csa_tree_add_51_79_groupi_n_736, csa_tree_add_51_79_groupi_n_737, csa_tree_add_51_79_groupi_n_739, csa_tree_add_51_79_groupi_n_739, csa_tree_add_51_79_groupi_n_740, csa_tree_add_51_79_groupi_n_742, csa_tree_add_51_79_groupi_n_742, csa_tree_add_51_79_groupi_n_743;
  wire csa_tree_add_51_79_groupi_n_745, csa_tree_add_51_79_groupi_n_745, csa_tree_add_51_79_groupi_n_746, csa_tree_add_51_79_groupi_n_748, csa_tree_add_51_79_groupi_n_748, csa_tree_add_51_79_groupi_n_749, csa_tree_add_51_79_groupi_n_751, csa_tree_add_51_79_groupi_n_751;
  wire csa_tree_add_51_79_groupi_n_1460, csa_tree_add_51_79_groupi_n_1122, csa_tree_add_51_79_groupi_n_1460, csa_tree_add_51_79_groupi_n_1454, csa_tree_add_51_79_groupi_n_1457, csa_tree_add_51_79_groupi_n_1122, csa_tree_add_51_79_groupi_n_1457, csa_tree_add_51_79_groupi_n_1448;
  wire csa_tree_add_51_79_groupi_n_764, csa_tree_add_51_79_groupi_n_765, csa_tree_add_51_79_groupi_n_4811, csa_tree_add_51_79_groupi_n_763, csa_tree_add_51_79_groupi_n_764, csa_tree_add_51_79_groupi_n_765, csa_tree_add_51_79_groupi_n_843, csa_tree_add_51_79_groupi_n_844;
  wire csa_tree_add_51_79_groupi_n_844, csa_tree_add_51_79_groupi_n_845, csa_tree_add_51_79_groupi_n_846, csa_tree_add_51_79_groupi_n_846, csa_tree_add_51_79_groupi_n_841, csa_tree_add_51_79_groupi_n_842, csa_tree_add_51_79_groupi_n_842, csa_tree_add_51_79_groupi_n_796;
  wire csa_tree_add_51_79_groupi_n_798, csa_tree_add_51_79_groupi_n_798, csa_tree_add_51_79_groupi_n_847, csa_tree_add_51_79_groupi_n_848, csa_tree_add_51_79_groupi_n_848, csa_tree_add_51_79_groupi_n_805, csa_tree_add_51_79_groupi_n_807, csa_tree_add_51_79_groupi_n_807;
  wire csa_tree_add_51_79_groupi_n_808, csa_tree_add_51_79_groupi_n_810, csa_tree_add_51_79_groupi_n_810, csa_tree_add_51_79_groupi_n_835, csa_tree_add_51_79_groupi_n_836, csa_tree_add_51_79_groupi_n_836, csa_tree_add_51_79_groupi_n_837, csa_tree_add_51_79_groupi_n_838;
  wire csa_tree_add_51_79_groupi_n_838, csa_tree_add_51_79_groupi_n_839, csa_tree_add_51_79_groupi_n_840, csa_tree_add_51_79_groupi_n_840, csa_tree_add_51_79_groupi_n_796, csa_tree_add_51_79_groupi_n_798, csa_tree_add_51_79_groupi_n_798, csa_tree_add_51_79_groupi_n_851;
  wire csa_tree_add_51_79_groupi_n_852, csa_tree_add_51_79_groupi_n_852, csa_tree_add_51_79_groupi_n_849, csa_tree_add_51_79_groupi_n_850, csa_tree_add_51_79_groupi_n_850, csa_tree_add_51_79_groupi_n_805, csa_tree_add_51_79_groupi_n_807, csa_tree_add_51_79_groupi_n_807;
  wire csa_tree_add_51_79_groupi_n_808, csa_tree_add_51_79_groupi_n_810, csa_tree_add_51_79_groupi_n_810, csa_tree_add_51_79_groupi_n_827, csa_tree_add_51_79_groupi_n_828, csa_tree_add_51_79_groupi_n_828, csa_tree_add_51_79_groupi_n_822, csa_tree_add_51_79_groupi_n_823;
  wire csa_tree_add_51_79_groupi_n_823, csa_tree_add_51_79_groupi_n_820, csa_tree_add_51_79_groupi_n_821, csa_tree_add_51_79_groupi_n_821, csa_tree_add_51_79_groupi_n_820, csa_tree_add_51_79_groupi_n_821, csa_tree_add_51_79_groupi_n_822, csa_tree_add_51_79_groupi_n_823;
  wire csa_tree_add_51_79_groupi_n_887, csa_tree_add_51_79_groupi_n_888, csa_tree_add_51_79_groupi_n_888, csa_tree_add_51_79_groupi_n_827, csa_tree_add_51_79_groupi_n_828, csa_tree_add_51_79_groupi_n_870, csa_tree_add_51_79_groupi_n_871, csa_tree_add_51_79_groupi_n_871;
  wire csa_tree_add_51_79_groupi_n_863, csa_tree_add_51_79_groupi_n_864, csa_tree_add_51_79_groupi_n_864, csa_tree_add_51_79_groupi_n_835, csa_tree_add_51_79_groupi_n_836, csa_tree_add_51_79_groupi_n_837, csa_tree_add_51_79_groupi_n_838, csa_tree_add_51_79_groupi_n_839;
  wire csa_tree_add_51_79_groupi_n_840, csa_tree_add_51_79_groupi_n_841, csa_tree_add_51_79_groupi_n_842, csa_tree_add_51_79_groupi_n_843, csa_tree_add_51_79_groupi_n_844, csa_tree_add_51_79_groupi_n_845, csa_tree_add_51_79_groupi_n_846, csa_tree_add_51_79_groupi_n_847;
  wire csa_tree_add_51_79_groupi_n_848, csa_tree_add_51_79_groupi_n_849, csa_tree_add_51_79_groupi_n_850, csa_tree_add_51_79_groupi_n_851, csa_tree_add_51_79_groupi_n_852, csa_tree_add_51_79_groupi_n_856, csa_tree_add_51_79_groupi_n_857, csa_tree_add_51_79_groupi_n_857;
  wire csa_tree_add_51_79_groupi_n_856, csa_tree_add_51_79_groupi_n_857, csa_tree_add_51_79_groupi_n_861, csa_tree_add_51_79_groupi_n_862, csa_tree_add_51_79_groupi_n_862, csa_tree_add_51_79_groupi_n_861, csa_tree_add_51_79_groupi_n_862, csa_tree_add_51_79_groupi_n_863;
  wire csa_tree_add_51_79_groupi_n_864, csa_tree_add_51_79_groupi_n_868, csa_tree_add_51_79_groupi_n_869, csa_tree_add_51_79_groupi_n_869, csa_tree_add_51_79_groupi_n_868, csa_tree_add_51_79_groupi_n_869, csa_tree_add_51_79_groupi_n_870, csa_tree_add_51_79_groupi_n_871;
  wire csa_tree_add_51_79_groupi_n_875, csa_tree_add_51_79_groupi_n_876, csa_tree_add_51_79_groupi_n_876, csa_tree_add_51_79_groupi_n_875, csa_tree_add_51_79_groupi_n_876, csa_tree_add_51_79_groupi_n_880, csa_tree_add_51_79_groupi_n_881, csa_tree_add_51_79_groupi_n_881;
  wire csa_tree_add_51_79_groupi_n_880, csa_tree_add_51_79_groupi_n_881, csa_tree_add_51_79_groupi_n_885, csa_tree_add_51_79_groupi_n_886, csa_tree_add_51_79_groupi_n_886, csa_tree_add_51_79_groupi_n_885, csa_tree_add_51_79_groupi_n_886, csa_tree_add_51_79_groupi_n_887;
  wire csa_tree_add_51_79_groupi_n_888, csa_tree_add_51_79_groupi_n_889, csa_tree_add_51_79_groupi_n_891, csa_tree_add_51_79_groupi_n_891, csa_tree_add_51_79_groupi_n_892, csa_tree_add_51_79_groupi_n_894, csa_tree_add_51_79_groupi_n_894, csa_tree_add_51_79_groupi_n_895;
  wire csa_tree_add_51_79_groupi_n_897, csa_tree_add_51_79_groupi_n_897, csa_tree_add_51_79_groupi_n_898, csa_tree_add_51_79_groupi_n_900, csa_tree_add_51_79_groupi_n_900, csa_tree_add_51_79_groupi_n_901, csa_tree_add_51_79_groupi_n_903, csa_tree_add_51_79_groupi_n_903;
  wire csa_tree_add_51_79_groupi_n_904, csa_tree_add_51_79_groupi_n_906, csa_tree_add_51_79_groupi_n_906, csa_tree_add_51_79_groupi_n_907, csa_tree_add_51_79_groupi_n_909, csa_tree_add_51_79_groupi_n_909, csa_tree_add_51_79_groupi_n_910, csa_tree_add_51_79_groupi_n_912;
  wire csa_tree_add_51_79_groupi_n_912, csa_tree_add_51_79_groupi_n_913, csa_tree_add_51_79_groupi_n_915, csa_tree_add_51_79_groupi_n_915, csa_tree_add_51_79_groupi_n_916, csa_tree_add_51_79_groupi_n_918, csa_tree_add_51_79_groupi_n_918, csa_tree_add_51_79_groupi_n_919;
  wire csa_tree_add_51_79_groupi_n_921, csa_tree_add_51_79_groupi_n_921, csa_tree_add_51_79_groupi_n_922, csa_tree_add_51_79_groupi_n_924, csa_tree_add_51_79_groupi_n_924, csa_tree_add_51_79_groupi_n_925, csa_tree_add_51_79_groupi_n_927, csa_tree_add_51_79_groupi_n_927;
  wire csa_tree_add_51_79_groupi_n_928, csa_tree_add_51_79_groupi_n_930, csa_tree_add_51_79_groupi_n_930, csa_tree_add_51_79_groupi_n_931, csa_tree_add_51_79_groupi_n_933, csa_tree_add_51_79_groupi_n_933, csa_tree_add_51_79_groupi_n_934, csa_tree_add_51_79_groupi_n_936;
  wire csa_tree_add_51_79_groupi_n_936, csa_tree_add_51_79_groupi_n_937, csa_tree_add_51_79_groupi_n_939, csa_tree_add_51_79_groupi_n_939, csa_tree_add_51_79_groupi_n_940, csa_tree_add_51_79_groupi_n_942, csa_tree_add_51_79_groupi_n_942, csa_tree_add_51_79_groupi_n_943;
  wire csa_tree_add_51_79_groupi_n_945, csa_tree_add_51_79_groupi_n_945, csa_tree_add_51_79_groupi_n_946, csa_tree_add_51_79_groupi_n_948, csa_tree_add_51_79_groupi_n_948, csa_tree_add_51_79_groupi_n_949, csa_tree_add_51_79_groupi_n_951, csa_tree_add_51_79_groupi_n_951;
  wire csa_tree_add_51_79_groupi_n_952, csa_tree_add_51_79_groupi_n_954, csa_tree_add_51_79_groupi_n_954, csa_tree_add_51_79_groupi_n_955, csa_tree_add_51_79_groupi_n_957, csa_tree_add_51_79_groupi_n_957, csa_tree_add_51_79_groupi_n_958, csa_tree_add_51_79_groupi_n_960;
  wire csa_tree_add_51_79_groupi_n_960, csa_tree_add_51_79_groupi_n_961, csa_tree_add_51_79_groupi_n_963, csa_tree_add_51_79_groupi_n_963, csa_tree_add_51_79_groupi_n_964, csa_tree_add_51_79_groupi_n_966, csa_tree_add_51_79_groupi_n_966, csa_tree_add_51_79_groupi_n_967;
  wire csa_tree_add_51_79_groupi_n_969, csa_tree_add_51_79_groupi_n_969, csa_tree_add_51_79_groupi_n_970, csa_tree_add_51_79_groupi_n_972, csa_tree_add_51_79_groupi_n_972, csa_tree_add_51_79_groupi_n_973, csa_tree_add_51_79_groupi_n_975, csa_tree_add_51_79_groupi_n_975;
  wire csa_tree_add_51_79_groupi_n_976, csa_tree_add_51_79_groupi_n_978, csa_tree_add_51_79_groupi_n_978, csa_tree_add_51_79_groupi_n_979, csa_tree_add_51_79_groupi_n_981, csa_tree_add_51_79_groupi_n_981, csa_tree_add_51_79_groupi_n_982, csa_tree_add_51_79_groupi_n_984;
  wire csa_tree_add_51_79_groupi_n_984, csa_tree_add_51_79_groupi_n_985, csa_tree_add_51_79_groupi_n_987, csa_tree_add_51_79_groupi_n_987, csa_tree_add_51_79_groupi_n_988, csa_tree_add_51_79_groupi_n_990, csa_tree_add_51_79_groupi_n_990, csa_tree_add_51_79_groupi_n_991;
  wire csa_tree_add_51_79_groupi_n_993, csa_tree_add_51_79_groupi_n_993, csa_tree_add_51_79_groupi_n_994, csa_tree_add_51_79_groupi_n_996, csa_tree_add_51_79_groupi_n_996, csa_tree_add_51_79_groupi_n_997, csa_tree_add_51_79_groupi_n_999, csa_tree_add_51_79_groupi_n_999;
  wire csa_tree_add_51_79_groupi_n_1000, csa_tree_add_51_79_groupi_n_1002, csa_tree_add_51_79_groupi_n_1002, csa_tree_add_51_79_groupi_n_1003, csa_tree_add_51_79_groupi_n_1005, csa_tree_add_51_79_groupi_n_1005, csa_tree_add_51_79_groupi_n_1006, csa_tree_add_51_79_groupi_n_1008;
  wire csa_tree_add_51_79_groupi_n_1008, csa_tree_add_51_79_groupi_n_1009, csa_tree_add_51_79_groupi_n_1011, csa_tree_add_51_79_groupi_n_1011, csa_tree_add_51_79_groupi_n_1012, csa_tree_add_51_79_groupi_n_1014, csa_tree_add_51_79_groupi_n_1014, csa_tree_add_51_79_groupi_n_1015;
  wire csa_tree_add_51_79_groupi_n_1017, csa_tree_add_51_79_groupi_n_1017, csa_tree_add_51_79_groupi_n_1018, csa_tree_add_51_79_groupi_n_1020, csa_tree_add_51_79_groupi_n_1020, csa_tree_add_51_79_groupi_n_1021, csa_tree_add_51_79_groupi_n_1023, csa_tree_add_51_79_groupi_n_1023;
  wire csa_tree_add_51_79_groupi_n_1024, csa_tree_add_51_79_groupi_n_1026, csa_tree_add_51_79_groupi_n_1026, csa_tree_add_51_79_groupi_n_1027, csa_tree_add_51_79_groupi_n_1029, csa_tree_add_51_79_groupi_n_1029, csa_tree_add_51_79_groupi_n_1030, csa_tree_add_51_79_groupi_n_1032;
  wire csa_tree_add_51_79_groupi_n_1032, csa_tree_add_51_79_groupi_n_1033, csa_tree_add_51_79_groupi_n_1035, csa_tree_add_51_79_groupi_n_1035, csa_tree_add_51_79_groupi_n_1036, csa_tree_add_51_79_groupi_n_1038, csa_tree_add_51_79_groupi_n_1038, csa_tree_add_51_79_groupi_n_1039;
  wire csa_tree_add_51_79_groupi_n_1041, csa_tree_add_51_79_groupi_n_1041, csa_tree_add_51_79_groupi_n_1042, csa_tree_add_51_79_groupi_n_1044, csa_tree_add_51_79_groupi_n_1044, csa_tree_add_51_79_groupi_n_1045, csa_tree_add_51_79_groupi_n_1047, csa_tree_add_51_79_groupi_n_1047;
  wire csa_tree_add_51_79_groupi_n_1048, csa_tree_add_51_79_groupi_n_1050, csa_tree_add_51_79_groupi_n_1050, csa_tree_add_51_79_groupi_n_1051, csa_tree_add_51_79_groupi_n_1053, csa_tree_add_51_79_groupi_n_1053, csa_tree_add_51_79_groupi_n_1054, csa_tree_add_51_79_groupi_n_1056;
  wire csa_tree_add_51_79_groupi_n_1056, csa_tree_add_51_79_groupi_n_1057, csa_tree_add_51_79_groupi_n_1059, csa_tree_add_51_79_groupi_n_1059, csa_tree_add_51_79_groupi_n_1060, csa_tree_add_51_79_groupi_n_1062, csa_tree_add_51_79_groupi_n_1062, csa_tree_add_51_79_groupi_n_1063;
  wire csa_tree_add_51_79_groupi_n_1065, csa_tree_add_51_79_groupi_n_1065, csa_tree_add_51_79_groupi_n_1066, csa_tree_add_51_79_groupi_n_1068, csa_tree_add_51_79_groupi_n_1068, csa_tree_add_51_79_groupi_n_1069, csa_tree_add_51_79_groupi_n_1070, csa_tree_add_51_79_groupi_n_1071;
  wire csa_tree_add_51_79_groupi_n_1072, csa_tree_add_51_79_groupi_n_1073, csa_tree_add_51_79_groupi_n_1074, csa_tree_add_51_79_groupi_n_1075, csa_tree_add_51_79_groupi_n_1076, csa_tree_add_51_79_groupi_n_1077, csa_tree_add_51_79_groupi_n_1078, csa_tree_add_51_79_groupi_n_1079;
  wire csa_tree_add_51_79_groupi_n_1080, csa_tree_add_51_79_groupi_n_1081, csa_tree_add_51_79_groupi_n_1082, csa_tree_add_51_79_groupi_n_1083, csa_tree_add_51_79_groupi_n_1084, csa_tree_add_51_79_groupi_n_1085, csa_tree_add_51_79_groupi_n_1086, csa_tree_add_51_79_groupi_n_1087;
  wire csa_tree_add_51_79_groupi_n_1088, csa_tree_add_51_79_groupi_n_1089, csa_tree_add_51_79_groupi_n_1090, csa_tree_add_51_79_groupi_n_1091, csa_tree_add_51_79_groupi_n_1092, csa_tree_add_51_79_groupi_n_1093, csa_tree_add_51_79_groupi_n_1094, csa_tree_add_51_79_groupi_n_1095;
  wire csa_tree_add_51_79_groupi_n_1096, csa_tree_add_51_79_groupi_n_1097, csa_tree_add_51_79_groupi_n_1098, csa_tree_add_51_79_groupi_n_1099, csa_tree_add_51_79_groupi_n_1100, csa_tree_add_51_79_groupi_n_1101, csa_tree_add_51_79_groupi_n_1102, csa_tree_add_51_79_groupi_n_1103;
  wire csa_tree_add_51_79_groupi_n_1104, csa_tree_add_51_79_groupi_n_1105, csa_tree_add_51_79_groupi_n_1106, csa_tree_add_51_79_groupi_n_1107, csa_tree_add_51_79_groupi_n_1108, csa_tree_add_51_79_groupi_n_1109, csa_tree_add_51_79_groupi_n_1110, csa_tree_add_51_79_groupi_n_1111;
  wire csa_tree_add_51_79_groupi_n_1112, csa_tree_add_51_79_groupi_n_1113, csa_tree_add_51_79_groupi_n_1114, csa_tree_add_51_79_groupi_n_1115, csa_tree_add_51_79_groupi_n_1457, csa_tree_add_51_79_groupi_n_1459, csa_tree_add_51_79_groupi_n_1459, csa_tree_add_51_79_groupi_n_1460;
  wire csa_tree_add_51_79_groupi_n_1462, csa_tree_add_51_79_groupi_n_1462, csa_tree_add_51_79_groupi_n_1122, csa_tree_add_51_79_groupi_n_1124, csa_tree_add_51_79_groupi_n_1124, csa_tree_add_51_79_groupi_n_1125, csa_tree_add_51_79_groupi_n_1126, csa_tree_add_51_79_groupi_n_1127;
  wire csa_tree_add_51_79_groupi_n_1128, csa_tree_add_51_79_groupi_n_1129, csa_tree_add_51_79_groupi_n_1130, csa_tree_add_51_79_groupi_n_1131, csa_tree_add_51_79_groupi_n_1132, csa_tree_add_51_79_groupi_n_1133, csa_tree_add_51_79_groupi_n_1134, csa_tree_add_51_79_groupi_n_1135;
  wire csa_tree_add_51_79_groupi_n_1136, csa_tree_add_51_79_groupi_n_1137, csa_tree_add_51_79_groupi_n_1138, csa_tree_add_51_79_groupi_n_1139, csa_tree_add_51_79_groupi_n_1140, csa_tree_add_51_79_groupi_n_1141, csa_tree_add_51_79_groupi_n_1142, csa_tree_add_51_79_groupi_n_1143;
  wire csa_tree_add_51_79_groupi_n_1144, csa_tree_add_51_79_groupi_n_1145, csa_tree_add_51_79_groupi_n_1146, csa_tree_add_51_79_groupi_n_1241, csa_tree_add_51_79_groupi_n_1217, csa_tree_add_51_79_groupi_n_2524, csa_tree_add_51_79_groupi_n_1082, csa_tree_add_51_79_groupi_n_2518;
  wire csa_tree_add_51_79_groupi_n_1078, csa_tree_add_51_79_groupi_n_2538, csa_tree_add_51_79_groupi_n_1084, csa_tree_add_51_79_groupi_n_1250, csa_tree_add_51_79_groupi_n_2515, csa_tree_add_51_79_groupi_n_1080, csa_tree_add_51_79_groupi_n_1232, csa_tree_add_51_79_groupi_n_1238;
  wire csa_tree_add_51_79_groupi_n_1256, csa_tree_add_51_79_groupi_n_1247, csa_tree_add_51_79_groupi_n_1229, csa_tree_add_51_79_groupi_n_1253, csa_tree_add_51_79_groupi_n_1220, csa_tree_add_51_79_groupi_n_1244, csa_tree_add_51_79_groupi_n_1262, csa_tree_add_51_79_groupi_n_1235;
  wire csa_tree_add_51_79_groupi_n_1259, csa_tree_add_51_79_groupi_n_1211, csa_tree_add_51_79_groupi_n_1214, csa_tree_add_51_79_groupi_n_1223, csa_tree_add_51_79_groupi_n_1226, csa_tree_add_51_79_groupi_n_1173, csa_tree_add_51_79_groupi_n_1174, csa_tree_add_51_79_groupi_n_1175;
  wire csa_tree_add_51_79_groupi_n_1176, csa_tree_add_51_79_groupi_n_1177, csa_tree_add_51_79_groupi_n_1178, csa_tree_add_51_79_groupi_n_1409, csa_tree_add_51_79_groupi_n_1403, csa_tree_add_51_79_groupi_n_1274, csa_tree_add_51_79_groupi_n_1292, csa_tree_add_51_79_groupi_n_1298;
  wire csa_tree_add_51_79_groupi_n_1427, csa_tree_add_51_79_groupi_n_1304, csa_tree_add_51_79_groupi_n_1316, csa_tree_add_51_79_groupi_n_1286, csa_tree_add_51_79_groupi_n_1328, csa_tree_add_51_79_groupi_n_1334, csa_tree_add_51_79_groupi_n_1442, csa_tree_add_51_79_groupi_n_1340;
  wire csa_tree_add_51_79_groupi_n_1310, csa_tree_add_51_79_groupi_n_1280, csa_tree_add_51_79_groupi_n_1352, csa_tree_add_51_79_groupi_n_1358, csa_tree_add_51_79_groupi_n_1367, csa_tree_add_51_79_groupi_n_1382, csa_tree_add_51_79_groupi_n_1391, csa_tree_add_51_79_groupi_n_1364;
  wire csa_tree_add_51_79_groupi_n_1415, csa_tree_add_51_79_groupi_n_1418, csa_tree_add_51_79_groupi_n_1322, csa_tree_add_51_79_groupi_n_1388, csa_tree_add_51_79_groupi_n_1271, csa_tree_add_51_79_groupi_n_1346, csa_tree_add_51_79_groupi_n_1373, csa_tree_add_51_79_groupi_n_1400;
  wire csa_tree_add_51_79_groupi_n_1436, csa_tree_add_51_79_groupi_n_1210, csa_tree_add_51_79_groupi_n_1210, csa_tree_add_51_79_groupi_n_1211, csa_tree_add_51_79_groupi_n_1213, csa_tree_add_51_79_groupi_n_1213, csa_tree_add_51_79_groupi_n_1214, csa_tree_add_51_79_groupi_n_1216;
  wire csa_tree_add_51_79_groupi_n_1216, csa_tree_add_51_79_groupi_n_1217, csa_tree_add_51_79_groupi_n_1219, csa_tree_add_51_79_groupi_n_1219, csa_tree_add_51_79_groupi_n_1220, csa_tree_add_51_79_groupi_n_1222, csa_tree_add_51_79_groupi_n_1222, csa_tree_add_51_79_groupi_n_1223;
  wire csa_tree_add_51_79_groupi_n_1225, csa_tree_add_51_79_groupi_n_1225, csa_tree_add_51_79_groupi_n_1226, csa_tree_add_51_79_groupi_n_1228, csa_tree_add_51_79_groupi_n_1228, csa_tree_add_51_79_groupi_n_1229, csa_tree_add_51_79_groupi_n_1231, csa_tree_add_51_79_groupi_n_1231;
  wire csa_tree_add_51_79_groupi_n_1232, csa_tree_add_51_79_groupi_n_1234, csa_tree_add_51_79_groupi_n_1234, csa_tree_add_51_79_groupi_n_1235, csa_tree_add_51_79_groupi_n_1237, csa_tree_add_51_79_groupi_n_1237, csa_tree_add_51_79_groupi_n_1238, csa_tree_add_51_79_groupi_n_1240;
  wire csa_tree_add_51_79_groupi_n_1240, csa_tree_add_51_79_groupi_n_1241, csa_tree_add_51_79_groupi_n_1243, csa_tree_add_51_79_groupi_n_1243, csa_tree_add_51_79_groupi_n_1244, csa_tree_add_51_79_groupi_n_1246, csa_tree_add_51_79_groupi_n_1246, csa_tree_add_51_79_groupi_n_1247;
  wire csa_tree_add_51_79_groupi_n_1249, csa_tree_add_51_79_groupi_n_1249, csa_tree_add_51_79_groupi_n_1250, csa_tree_add_51_79_groupi_n_1252, csa_tree_add_51_79_groupi_n_1252, csa_tree_add_51_79_groupi_n_1253, csa_tree_add_51_79_groupi_n_1255, csa_tree_add_51_79_groupi_n_1255;
  wire csa_tree_add_51_79_groupi_n_1256, csa_tree_add_51_79_groupi_n_1258, csa_tree_add_51_79_groupi_n_1258, csa_tree_add_51_79_groupi_n_1259, csa_tree_add_51_79_groupi_n_1261, csa_tree_add_51_79_groupi_n_1261, csa_tree_add_51_79_groupi_n_1262, csa_tree_add_51_79_groupi_n_1264;
  wire csa_tree_add_51_79_groupi_n_1264, csa_tree_add_51_79_groupi_n_1265, csa_tree_add_51_79_groupi_n_1267, csa_tree_add_51_79_groupi_n_1267, csa_tree_add_51_79_groupi_n_1268, csa_tree_add_51_79_groupi_n_1270, csa_tree_add_51_79_groupi_n_1270, csa_tree_add_51_79_groupi_n_1271;
  wire csa_tree_add_51_79_groupi_n_1273, csa_tree_add_51_79_groupi_n_1273, csa_tree_add_51_79_groupi_n_1274, csa_tree_add_51_79_groupi_n_1276, csa_tree_add_51_79_groupi_n_1276, csa_tree_add_51_79_groupi_n_1277, csa_tree_add_51_79_groupi_n_1279, csa_tree_add_51_79_groupi_n_1279;
  wire csa_tree_add_51_79_groupi_n_1280, csa_tree_add_51_79_groupi_n_1282, csa_tree_add_51_79_groupi_n_1282, csa_tree_add_51_79_groupi_n_1283, csa_tree_add_51_79_groupi_n_1285, csa_tree_add_51_79_groupi_n_1285, csa_tree_add_51_79_groupi_n_1286, csa_tree_add_51_79_groupi_n_1288;
  wire csa_tree_add_51_79_groupi_n_1288, csa_tree_add_51_79_groupi_n_1289, csa_tree_add_51_79_groupi_n_1291, csa_tree_add_51_79_groupi_n_1291, csa_tree_add_51_79_groupi_n_1292, csa_tree_add_51_79_groupi_n_1294, csa_tree_add_51_79_groupi_n_1294, csa_tree_add_51_79_groupi_n_1295;
  wire csa_tree_add_51_79_groupi_n_1297, csa_tree_add_51_79_groupi_n_1297, csa_tree_add_51_79_groupi_n_1298, csa_tree_add_51_79_groupi_n_1300, csa_tree_add_51_79_groupi_n_1300, csa_tree_add_51_79_groupi_n_1301, csa_tree_add_51_79_groupi_n_1303, csa_tree_add_51_79_groupi_n_1303;
  wire csa_tree_add_51_79_groupi_n_1304, csa_tree_add_51_79_groupi_n_1306, csa_tree_add_51_79_groupi_n_1306, csa_tree_add_51_79_groupi_n_1307, csa_tree_add_51_79_groupi_n_1309, csa_tree_add_51_79_groupi_n_1309, csa_tree_add_51_79_groupi_n_1310, csa_tree_add_51_79_groupi_n_1312;
  wire csa_tree_add_51_79_groupi_n_1312, csa_tree_add_51_79_groupi_n_1313, csa_tree_add_51_79_groupi_n_1315, csa_tree_add_51_79_groupi_n_1315, csa_tree_add_51_79_groupi_n_1316, csa_tree_add_51_79_groupi_n_1318, csa_tree_add_51_79_groupi_n_1318, csa_tree_add_51_79_groupi_n_1319;
  wire csa_tree_add_51_79_groupi_n_1321, csa_tree_add_51_79_groupi_n_1321, csa_tree_add_51_79_groupi_n_1322, csa_tree_add_51_79_groupi_n_1324, csa_tree_add_51_79_groupi_n_1324, csa_tree_add_51_79_groupi_n_1325, csa_tree_add_51_79_groupi_n_1327, csa_tree_add_51_79_groupi_n_1327;
  wire csa_tree_add_51_79_groupi_n_1328, csa_tree_add_51_79_groupi_n_1330, csa_tree_add_51_79_groupi_n_1330, csa_tree_add_51_79_groupi_n_1331, csa_tree_add_51_79_groupi_n_1333, csa_tree_add_51_79_groupi_n_1333, csa_tree_add_51_79_groupi_n_1334, csa_tree_add_51_79_groupi_n_1336;
  wire csa_tree_add_51_79_groupi_n_1336, csa_tree_add_51_79_groupi_n_1337, csa_tree_add_51_79_groupi_n_1339, csa_tree_add_51_79_groupi_n_1339, csa_tree_add_51_79_groupi_n_1340, csa_tree_add_51_79_groupi_n_1342, csa_tree_add_51_79_groupi_n_1342, csa_tree_add_51_79_groupi_n_1343;
  wire csa_tree_add_51_79_groupi_n_1345, csa_tree_add_51_79_groupi_n_1345, csa_tree_add_51_79_groupi_n_1346, csa_tree_add_51_79_groupi_n_1348, csa_tree_add_51_79_groupi_n_1348, csa_tree_add_51_79_groupi_n_1349, csa_tree_add_51_79_groupi_n_1351, csa_tree_add_51_79_groupi_n_1351;
  wire csa_tree_add_51_79_groupi_n_1352, csa_tree_add_51_79_groupi_n_1354, csa_tree_add_51_79_groupi_n_1354, csa_tree_add_51_79_groupi_n_1355, csa_tree_add_51_79_groupi_n_1357, csa_tree_add_51_79_groupi_n_1357, csa_tree_add_51_79_groupi_n_1358, csa_tree_add_51_79_groupi_n_1360;
  wire csa_tree_add_51_79_groupi_n_1360, csa_tree_add_51_79_groupi_n_1361, csa_tree_add_51_79_groupi_n_1363, csa_tree_add_51_79_groupi_n_1363, csa_tree_add_51_79_groupi_n_1364, csa_tree_add_51_79_groupi_n_1366, csa_tree_add_51_79_groupi_n_1366, csa_tree_add_51_79_groupi_n_1367;
  wire csa_tree_add_51_79_groupi_n_1369, csa_tree_add_51_79_groupi_n_1369, csa_tree_add_51_79_groupi_n_1370, csa_tree_add_51_79_groupi_n_1372, csa_tree_add_51_79_groupi_n_1372, csa_tree_add_51_79_groupi_n_1373, csa_tree_add_51_79_groupi_n_1375, csa_tree_add_51_79_groupi_n_1375;
  wire csa_tree_add_51_79_groupi_n_1376, csa_tree_add_51_79_groupi_n_1378, csa_tree_add_51_79_groupi_n_1378, csa_tree_add_51_79_groupi_n_1379, csa_tree_add_51_79_groupi_n_1381, csa_tree_add_51_79_groupi_n_1381, csa_tree_add_51_79_groupi_n_1382, csa_tree_add_51_79_groupi_n_1384;
  wire csa_tree_add_51_79_groupi_n_1384, csa_tree_add_51_79_groupi_n_1385, csa_tree_add_51_79_groupi_n_1387, csa_tree_add_51_79_groupi_n_1387, csa_tree_add_51_79_groupi_n_1388, csa_tree_add_51_79_groupi_n_1390, csa_tree_add_51_79_groupi_n_1390, csa_tree_add_51_79_groupi_n_1391;
  wire csa_tree_add_51_79_groupi_n_1393, csa_tree_add_51_79_groupi_n_1393, csa_tree_add_51_79_groupi_n_1394, csa_tree_add_51_79_groupi_n_1396, csa_tree_add_51_79_groupi_n_1396, csa_tree_add_51_79_groupi_n_1397, csa_tree_add_51_79_groupi_n_1399, csa_tree_add_51_79_groupi_n_1399;
  wire csa_tree_add_51_79_groupi_n_1400, csa_tree_add_51_79_groupi_n_1402, csa_tree_add_51_79_groupi_n_1402, csa_tree_add_51_79_groupi_n_1403, csa_tree_add_51_79_groupi_n_1405, csa_tree_add_51_79_groupi_n_1405, csa_tree_add_51_79_groupi_n_1406, csa_tree_add_51_79_groupi_n_1408;
  wire csa_tree_add_51_79_groupi_n_1408, csa_tree_add_51_79_groupi_n_1409, csa_tree_add_51_79_groupi_n_1411, csa_tree_add_51_79_groupi_n_1411, csa_tree_add_51_79_groupi_n_1412, csa_tree_add_51_79_groupi_n_1414, csa_tree_add_51_79_groupi_n_1414, csa_tree_add_51_79_groupi_n_1415;
  wire csa_tree_add_51_79_groupi_n_1417, csa_tree_add_51_79_groupi_n_1417, csa_tree_add_51_79_groupi_n_1418, csa_tree_add_51_79_groupi_n_1420, csa_tree_add_51_79_groupi_n_1420, csa_tree_add_51_79_groupi_n_1421, csa_tree_add_51_79_groupi_n_1423, csa_tree_add_51_79_groupi_n_1423;
  wire csa_tree_add_51_79_groupi_n_1424, csa_tree_add_51_79_groupi_n_1426, csa_tree_add_51_79_groupi_n_1426, csa_tree_add_51_79_groupi_n_1427, csa_tree_add_51_79_groupi_n_1429, csa_tree_add_51_79_groupi_n_1429, csa_tree_add_51_79_groupi_n_1430, csa_tree_add_51_79_groupi_n_1432;
  wire csa_tree_add_51_79_groupi_n_1432, csa_tree_add_51_79_groupi_n_1433, csa_tree_add_51_79_groupi_n_1435, csa_tree_add_51_79_groupi_n_1435, csa_tree_add_51_79_groupi_n_1436, csa_tree_add_51_79_groupi_n_1438, csa_tree_add_51_79_groupi_n_1438, csa_tree_add_51_79_groupi_n_1439;
  wire csa_tree_add_51_79_groupi_n_1441, csa_tree_add_51_79_groupi_n_1441, csa_tree_add_51_79_groupi_n_1442, csa_tree_add_51_79_groupi_n_1444, csa_tree_add_51_79_groupi_n_1444, csa_tree_add_51_79_groupi_n_1448, csa_tree_add_51_79_groupi_n_1450, csa_tree_add_51_79_groupi_n_1450;
  wire csa_tree_add_51_79_groupi_n_1448, csa_tree_add_51_79_groupi_n_1450, csa_tree_add_51_79_groupi_n_1450, csa_tree_add_51_79_groupi_n_1454, csa_tree_add_51_79_groupi_n_1456, csa_tree_add_51_79_groupi_n_1456, csa_tree_add_51_79_groupi_n_1454, csa_tree_add_51_79_groupi_n_1456;
  wire csa_tree_add_51_79_groupi_n_1456, csa_tree_add_51_79_groupi_n_1457, csa_tree_add_51_79_groupi_n_1459, csa_tree_add_51_79_groupi_n_1459, csa_tree_add_51_79_groupi_n_1460, csa_tree_add_51_79_groupi_n_1462, csa_tree_add_51_79_groupi_n_1462, csa_tree_add_51_79_groupi_n_1122;
  wire csa_tree_add_51_79_groupi_n_1124, csa_tree_add_51_79_groupi_n_1124, csa_tree_add_51_79_groupi_n_1466, csa_tree_add_51_79_groupi_n_1467, csa_tree_add_51_79_groupi_n_1468, csa_tree_add_51_79_groupi_n_1469, csa_tree_add_51_79_groupi_n_1470, csa_tree_add_51_79_groupi_n_1471;
  wire csa_tree_add_51_79_groupi_n_1970, csa_tree_add_51_79_groupi_n_1973, csa_tree_add_51_79_groupi_n_1976, csa_tree_add_51_79_groupi_n_1475, csa_tree_add_51_79_groupi_n_1476, csa_tree_add_51_79_groupi_n_1477, csa_tree_add_51_79_groupi_n_1478, csa_tree_add_51_79_groupi_n_1479;
  wire csa_tree_add_51_79_groupi_n_1480, csa_tree_add_51_79_groupi_n_1481, csa_tree_add_51_79_groupi_n_1482, csa_tree_add_51_79_groupi_n_1995, csa_tree_add_51_79_groupi_n_1484, csa_tree_add_51_79_groupi_n_1485, csa_tree_add_51_79_groupi_n_2002, csa_tree_add_51_79_groupi_n_2005;
  wire csa_tree_add_51_79_groupi_n_2008, csa_tree_add_51_79_groupi_n_2011, csa_tree_add_51_79_groupi_n_2014, csa_tree_add_51_79_groupi_n_1491, csa_tree_add_51_79_groupi_n_2438, csa_tree_add_51_79_groupi_n_2441, csa_tree_add_51_79_groupi_n_2444, csa_tree_add_51_79_groupi_n_1495;
  wire csa_tree_add_51_79_groupi_n_2449, csa_tree_add_51_79_groupi_n_2452, csa_tree_add_51_79_groupi_n_1498, csa_tree_add_51_79_groupi_n_2457, csa_tree_add_51_79_groupi_n_2460, csa_tree_add_51_79_groupi_n_2463, csa_tree_add_51_79_groupi_n_2466, csa_tree_add_51_79_groupi_n_2469;
  wire csa_tree_add_51_79_groupi_n_2472, csa_tree_add_51_79_groupi_n_2475, csa_tree_add_51_79_groupi_n_2478, csa_tree_add_51_79_groupi_n_1507, csa_tree_add_51_79_groupi_n_2483, csa_tree_add_51_79_groupi_n_2486, csa_tree_add_51_79_groupi_n_1510, csa_tree_add_51_79_groupi_n_2491;
  wire csa_tree_add_51_79_groupi_n_2494, csa_tree_add_51_79_groupi_n_2497, csa_tree_add_51_79_groupi_n_2500, csa_tree_add_51_79_groupi_n_1515, csa_tree_add_51_79_groupi_n_2505, csa_tree_add_51_79_groupi_n_1517, csa_tree_add_51_79_groupi_n_2510, csa_tree_add_51_79_groupi_n_1519;
  wire csa_tree_add_51_79_groupi_n_2513, csa_tree_add_51_79_groupi_n_1521, csa_tree_add_51_79_groupi_n_1521, csa_tree_add_51_79_groupi_n_2522, csa_tree_add_51_79_groupi_n_1524, csa_tree_add_51_79_groupi_n_1524, csa_tree_add_51_79_groupi_n_1527, csa_tree_add_51_79_groupi_n_1527;
  wire csa_tree_add_51_79_groupi_n_1528, csa_tree_add_51_79_groupi_n_1529, csa_tree_add_51_79_groupi_n_1530, csa_tree_add_51_79_groupi_n_1531, csa_tree_add_51_79_groupi_n_1532, csa_tree_add_51_79_groupi_n_1533, csa_tree_add_51_79_groupi_n_1534, csa_tree_add_51_79_groupi_n_1535;
  wire csa_tree_add_51_79_groupi_n_1536, csa_tree_add_51_79_groupi_n_1537, csa_tree_add_51_79_groupi_n_1538, csa_tree_add_51_79_groupi_n_1539, csa_tree_add_51_79_groupi_n_1540, csa_tree_add_51_79_groupi_n_1541, csa_tree_add_51_79_groupi_n_1542, csa_tree_add_51_79_groupi_n_1543;
  wire csa_tree_add_51_79_groupi_n_1544, csa_tree_add_51_79_groupi_n_1545, csa_tree_add_51_79_groupi_n_1546, csa_tree_add_51_79_groupi_n_1547, csa_tree_add_51_79_groupi_n_1548, csa_tree_add_51_79_groupi_n_1549, csa_tree_add_51_79_groupi_n_1550, csa_tree_add_51_79_groupi_n_1551;
  wire csa_tree_add_51_79_groupi_n_1552, csa_tree_add_51_79_groupi_n_1553, csa_tree_add_51_79_groupi_n_1554, csa_tree_add_51_79_groupi_n_1555, csa_tree_add_51_79_groupi_n_1556, csa_tree_add_51_79_groupi_n_1557, csa_tree_add_51_79_groupi_n_1558, csa_tree_add_51_79_groupi_n_1559;
  wire csa_tree_add_51_79_groupi_n_1560, csa_tree_add_51_79_groupi_n_1561, csa_tree_add_51_79_groupi_n_1562, csa_tree_add_51_79_groupi_n_1563, csa_tree_add_51_79_groupi_n_1564, csa_tree_add_51_79_groupi_n_1565, csa_tree_add_51_79_groupi_n_1566, csa_tree_add_51_79_groupi_n_1567;
  wire csa_tree_add_51_79_groupi_n_1568, csa_tree_add_51_79_groupi_n_1569, csa_tree_add_51_79_groupi_n_1570, csa_tree_add_51_79_groupi_n_1571, csa_tree_add_51_79_groupi_n_1572, csa_tree_add_51_79_groupi_n_1573, csa_tree_add_51_79_groupi_n_1574, csa_tree_add_51_79_groupi_n_1575;
  wire csa_tree_add_51_79_groupi_n_1576, csa_tree_add_51_79_groupi_n_1577, csa_tree_add_51_79_groupi_n_1578, csa_tree_add_51_79_groupi_n_1579, csa_tree_add_51_79_groupi_n_1580, csa_tree_add_51_79_groupi_n_1581, csa_tree_add_51_79_groupi_n_1582, csa_tree_add_51_79_groupi_n_1583;
  wire csa_tree_add_51_79_groupi_n_1584, csa_tree_add_51_79_groupi_n_1585, csa_tree_add_51_79_groupi_n_1586, csa_tree_add_51_79_groupi_n_1587, csa_tree_add_51_79_groupi_n_1588, csa_tree_add_51_79_groupi_n_1589, csa_tree_add_51_79_groupi_n_1590, csa_tree_add_51_79_groupi_n_1591;
  wire csa_tree_add_51_79_groupi_n_1592, csa_tree_add_51_79_groupi_n_1593, csa_tree_add_51_79_groupi_n_1594, csa_tree_add_51_79_groupi_n_1595, csa_tree_add_51_79_groupi_n_1596, csa_tree_add_51_79_groupi_n_1597, csa_tree_add_51_79_groupi_n_1598, csa_tree_add_51_79_groupi_n_1599;
  wire csa_tree_add_51_79_groupi_n_1600, csa_tree_add_51_79_groupi_n_1601, csa_tree_add_51_79_groupi_n_1602, csa_tree_add_51_79_groupi_n_1603, csa_tree_add_51_79_groupi_n_1604, csa_tree_add_51_79_groupi_n_1605, csa_tree_add_51_79_groupi_n_1606, csa_tree_add_51_79_groupi_n_1607;
  wire csa_tree_add_51_79_groupi_n_1608, csa_tree_add_51_79_groupi_n_1609, csa_tree_add_51_79_groupi_n_1610, csa_tree_add_51_79_groupi_n_1611, csa_tree_add_51_79_groupi_n_1612, csa_tree_add_51_79_groupi_n_1613, csa_tree_add_51_79_groupi_n_1614, csa_tree_add_51_79_groupi_n_1615;
  wire csa_tree_add_51_79_groupi_n_1616, csa_tree_add_51_79_groupi_n_1617, csa_tree_add_51_79_groupi_n_1618, csa_tree_add_51_79_groupi_n_1619, csa_tree_add_51_79_groupi_n_1620, csa_tree_add_51_79_groupi_n_1621, csa_tree_add_51_79_groupi_n_1622, csa_tree_add_51_79_groupi_n_1623;
  wire csa_tree_add_51_79_groupi_n_1624, csa_tree_add_51_79_groupi_n_1625, csa_tree_add_51_79_groupi_n_1626, csa_tree_add_51_79_groupi_n_1627, csa_tree_add_51_79_groupi_n_1628, csa_tree_add_51_79_groupi_n_1629, csa_tree_add_51_79_groupi_n_1630, csa_tree_add_51_79_groupi_n_1631;
  wire csa_tree_add_51_79_groupi_n_1632, csa_tree_add_51_79_groupi_n_1633, csa_tree_add_51_79_groupi_n_1634, csa_tree_add_51_79_groupi_n_1635, csa_tree_add_51_79_groupi_n_1636, csa_tree_add_51_79_groupi_n_1637, csa_tree_add_51_79_groupi_n_1638, csa_tree_add_51_79_groupi_n_1639;
  wire csa_tree_add_51_79_groupi_n_1640, csa_tree_add_51_79_groupi_n_1641, csa_tree_add_51_79_groupi_n_1642, csa_tree_add_51_79_groupi_n_1643, csa_tree_add_51_79_groupi_n_1644, csa_tree_add_51_79_groupi_n_1645, csa_tree_add_51_79_groupi_n_1646, csa_tree_add_51_79_groupi_n_1647;
  wire csa_tree_add_51_79_groupi_n_1648, csa_tree_add_51_79_groupi_n_1649, csa_tree_add_51_79_groupi_n_1650, csa_tree_add_51_79_groupi_n_1651, csa_tree_add_51_79_groupi_n_1652, csa_tree_add_51_79_groupi_n_1653, csa_tree_add_51_79_groupi_n_1654, csa_tree_add_51_79_groupi_n_1655;
  wire csa_tree_add_51_79_groupi_n_1656, csa_tree_add_51_79_groupi_n_1657, csa_tree_add_51_79_groupi_n_1658, csa_tree_add_51_79_groupi_n_1659, csa_tree_add_51_79_groupi_n_1660, csa_tree_add_51_79_groupi_n_1661, csa_tree_add_51_79_groupi_n_1662, csa_tree_add_51_79_groupi_n_1663;
  wire csa_tree_add_51_79_groupi_n_1664, csa_tree_add_51_79_groupi_n_1665, csa_tree_add_51_79_groupi_n_1666, csa_tree_add_51_79_groupi_n_1667, csa_tree_add_51_79_groupi_n_1668, csa_tree_add_51_79_groupi_n_1669, csa_tree_add_51_79_groupi_n_1670, csa_tree_add_51_79_groupi_n_1671;
  wire csa_tree_add_51_79_groupi_n_1672, csa_tree_add_51_79_groupi_n_1673, csa_tree_add_51_79_groupi_n_1674, csa_tree_add_51_79_groupi_n_1675, csa_tree_add_51_79_groupi_n_1676, csa_tree_add_51_79_groupi_n_1677, csa_tree_add_51_79_groupi_n_1678, csa_tree_add_51_79_groupi_n_1679;
  wire csa_tree_add_51_79_groupi_n_1680, csa_tree_add_51_79_groupi_n_1681, csa_tree_add_51_79_groupi_n_1682, csa_tree_add_51_79_groupi_n_1683, csa_tree_add_51_79_groupi_n_1684, csa_tree_add_51_79_groupi_n_1685, csa_tree_add_51_79_groupi_n_1686, csa_tree_add_51_79_groupi_n_1687;
  wire csa_tree_add_51_79_groupi_n_1688, csa_tree_add_51_79_groupi_n_1689, csa_tree_add_51_79_groupi_n_1690, csa_tree_add_51_79_groupi_n_1691, csa_tree_add_51_79_groupi_n_1692, csa_tree_add_51_79_groupi_n_1693, csa_tree_add_51_79_groupi_n_1694, csa_tree_add_51_79_groupi_n_1695;
  wire csa_tree_add_51_79_groupi_n_1696, csa_tree_add_51_79_groupi_n_1697, csa_tree_add_51_79_groupi_n_1698, csa_tree_add_51_79_groupi_n_1699, csa_tree_add_51_79_groupi_n_1700, csa_tree_add_51_79_groupi_n_1701, csa_tree_add_51_79_groupi_n_1702, csa_tree_add_51_79_groupi_n_1703;
  wire csa_tree_add_51_79_groupi_n_1704, csa_tree_add_51_79_groupi_n_1705, csa_tree_add_51_79_groupi_n_1706, csa_tree_add_51_79_groupi_n_1707, csa_tree_add_51_79_groupi_n_1708, csa_tree_add_51_79_groupi_n_1709, csa_tree_add_51_79_groupi_n_1710, csa_tree_add_51_79_groupi_n_1711;
  wire csa_tree_add_51_79_groupi_n_1712, csa_tree_add_51_79_groupi_n_1713, csa_tree_add_51_79_groupi_n_1714, csa_tree_add_51_79_groupi_n_1715, csa_tree_add_51_79_groupi_n_1716, csa_tree_add_51_79_groupi_n_1717, csa_tree_add_51_79_groupi_n_1718, csa_tree_add_51_79_groupi_n_1719;
  wire csa_tree_add_51_79_groupi_n_1720, csa_tree_add_51_79_groupi_n_1721, csa_tree_add_51_79_groupi_n_1722, csa_tree_add_51_79_groupi_n_1723, csa_tree_add_51_79_groupi_n_1724, csa_tree_add_51_79_groupi_n_1725, csa_tree_add_51_79_groupi_n_1726, csa_tree_add_51_79_groupi_n_1727;
  wire csa_tree_add_51_79_groupi_n_1728, csa_tree_add_51_79_groupi_n_1729, csa_tree_add_51_79_groupi_n_1730, csa_tree_add_51_79_groupi_n_1731, csa_tree_add_51_79_groupi_n_1732, csa_tree_add_51_79_groupi_n_1733, csa_tree_add_51_79_groupi_n_1734, csa_tree_add_51_79_groupi_n_1735;
  wire csa_tree_add_51_79_groupi_n_1736, csa_tree_add_51_79_groupi_n_1737, csa_tree_add_51_79_groupi_n_1738, csa_tree_add_51_79_groupi_n_1739, csa_tree_add_51_79_groupi_n_1740, csa_tree_add_51_79_groupi_n_1741, csa_tree_add_51_79_groupi_n_1742, csa_tree_add_51_79_groupi_n_1743;
  wire csa_tree_add_51_79_groupi_n_1744, csa_tree_add_51_79_groupi_n_1745, csa_tree_add_51_79_groupi_n_1746, csa_tree_add_51_79_groupi_n_1747, csa_tree_add_51_79_groupi_n_1748, csa_tree_add_51_79_groupi_n_1749, csa_tree_add_51_79_groupi_n_1750, csa_tree_add_51_79_groupi_n_1751;
  wire csa_tree_add_51_79_groupi_n_1752, csa_tree_add_51_79_groupi_n_1753, csa_tree_add_51_79_groupi_n_1754, csa_tree_add_51_79_groupi_n_1755, csa_tree_add_51_79_groupi_n_1756, csa_tree_add_51_79_groupi_n_1757, csa_tree_add_51_79_groupi_n_1758, csa_tree_add_51_79_groupi_n_1759;
  wire csa_tree_add_51_79_groupi_n_1760, csa_tree_add_51_79_groupi_n_1761, csa_tree_add_51_79_groupi_n_1762, csa_tree_add_51_79_groupi_n_1763, csa_tree_add_51_79_groupi_n_1764, csa_tree_add_51_79_groupi_n_1765, csa_tree_add_51_79_groupi_n_1766, csa_tree_add_51_79_groupi_n_1767;
  wire csa_tree_add_51_79_groupi_n_1768, csa_tree_add_51_79_groupi_n_1769, csa_tree_add_51_79_groupi_n_1770, csa_tree_add_51_79_groupi_n_1771, csa_tree_add_51_79_groupi_n_1772, csa_tree_add_51_79_groupi_n_1773, csa_tree_add_51_79_groupi_n_1774, csa_tree_add_51_79_groupi_n_1775;
  wire csa_tree_add_51_79_groupi_n_1776, csa_tree_add_51_79_groupi_n_1777, csa_tree_add_51_79_groupi_n_1778, csa_tree_add_51_79_groupi_n_1779, csa_tree_add_51_79_groupi_n_1780, csa_tree_add_51_79_groupi_n_1781, csa_tree_add_51_79_groupi_n_1782, csa_tree_add_51_79_groupi_n_1783;
  wire csa_tree_add_51_79_groupi_n_1784, csa_tree_add_51_79_groupi_n_1785, csa_tree_add_51_79_groupi_n_1786, csa_tree_add_51_79_groupi_n_1787, csa_tree_add_51_79_groupi_n_1788, csa_tree_add_51_79_groupi_n_1789, csa_tree_add_51_79_groupi_n_1790, csa_tree_add_51_79_groupi_n_1791;
  wire csa_tree_add_51_79_groupi_n_1792, csa_tree_add_51_79_groupi_n_1793, csa_tree_add_51_79_groupi_n_1794, csa_tree_add_51_79_groupi_n_1795, csa_tree_add_51_79_groupi_n_1796, csa_tree_add_51_79_groupi_n_1797, csa_tree_add_51_79_groupi_n_1798, csa_tree_add_51_79_groupi_n_1799;
  wire csa_tree_add_51_79_groupi_n_1800, csa_tree_add_51_79_groupi_n_1801, csa_tree_add_51_79_groupi_n_1802, csa_tree_add_51_79_groupi_n_1803, csa_tree_add_51_79_groupi_n_1804, csa_tree_add_51_79_groupi_n_1805, csa_tree_add_51_79_groupi_n_1806, csa_tree_add_51_79_groupi_n_1807;
  wire csa_tree_add_51_79_groupi_n_1808, csa_tree_add_51_79_groupi_n_1809, csa_tree_add_51_79_groupi_n_1810, csa_tree_add_51_79_groupi_n_1811, csa_tree_add_51_79_groupi_n_1812, csa_tree_add_51_79_groupi_n_1813, csa_tree_add_51_79_groupi_n_1814, csa_tree_add_51_79_groupi_n_1815;
  wire csa_tree_add_51_79_groupi_n_1816, csa_tree_add_51_79_groupi_n_1817, csa_tree_add_51_79_groupi_n_1818, csa_tree_add_51_79_groupi_n_1540, csa_tree_add_51_79_groupi_n_1820, csa_tree_add_51_79_groupi_n_1821, csa_tree_add_51_79_groupi_n_1822, csa_tree_add_51_79_groupi_n_1823;
  wire csa_tree_add_51_79_groupi_n_1824, csa_tree_add_51_79_groupi_n_1825, csa_tree_add_51_79_groupi_n_1826, csa_tree_add_51_79_groupi_n_1827, csa_tree_add_51_79_groupi_n_1828, csa_tree_add_51_79_groupi_n_1829, csa_tree_add_51_79_groupi_n_1830, csa_tree_add_51_79_groupi_n_1831;
  wire csa_tree_add_51_79_groupi_n_1832, csa_tree_add_51_79_groupi_n_1833, csa_tree_add_51_79_groupi_n_1834, csa_tree_add_51_79_groupi_n_1835, csa_tree_add_51_79_groupi_n_1836, csa_tree_add_51_79_groupi_n_1837, csa_tree_add_51_79_groupi_n_1838, csa_tree_add_51_79_groupi_n_1839;
  wire csa_tree_add_51_79_groupi_n_1840, csa_tree_add_51_79_groupi_n_1841, csa_tree_add_51_79_groupi_n_1842, csa_tree_add_51_79_groupi_n_1843, csa_tree_add_51_79_groupi_n_1844, csa_tree_add_51_79_groupi_n_1845, csa_tree_add_51_79_groupi_n_1846, csa_tree_add_51_79_groupi_n_1847;
  wire csa_tree_add_51_79_groupi_n_1848, csa_tree_add_51_79_groupi_n_1849, csa_tree_add_51_79_groupi_n_1850, csa_tree_add_51_79_groupi_n_1851, csa_tree_add_51_79_groupi_n_1852, csa_tree_add_51_79_groupi_n_1853, csa_tree_add_51_79_groupi_n_1854, csa_tree_add_51_79_groupi_n_1855;
  wire csa_tree_add_51_79_groupi_n_1856, csa_tree_add_51_79_groupi_n_1857, csa_tree_add_51_79_groupi_n_1858, csa_tree_add_51_79_groupi_n_1859, csa_tree_add_51_79_groupi_n_1860, csa_tree_add_51_79_groupi_n_1861, csa_tree_add_51_79_groupi_n_1862, csa_tree_add_51_79_groupi_n_1863;
  wire csa_tree_add_51_79_groupi_n_1864, csa_tree_add_51_79_groupi_n_1865, csa_tree_add_51_79_groupi_n_1866, csa_tree_add_51_79_groupi_n_1867, csa_tree_add_51_79_groupi_n_1868, csa_tree_add_51_79_groupi_n_1869, csa_tree_add_51_79_groupi_n_1870, csa_tree_add_51_79_groupi_n_1871;
  wire csa_tree_add_51_79_groupi_n_1872, csa_tree_add_51_79_groupi_n_1873, csa_tree_add_51_79_groupi_n_1874, csa_tree_add_51_79_groupi_n_1875, csa_tree_add_51_79_groupi_n_1876, csa_tree_add_51_79_groupi_n_1877, csa_tree_add_51_79_groupi_n_1878, csa_tree_add_51_79_groupi_n_1879;
  wire csa_tree_add_51_79_groupi_n_1880, csa_tree_add_51_79_groupi_n_1881, csa_tree_add_51_79_groupi_n_1882, csa_tree_add_51_79_groupi_n_1883, csa_tree_add_51_79_groupi_n_1884, csa_tree_add_51_79_groupi_n_1885, csa_tree_add_51_79_groupi_n_1886, csa_tree_add_51_79_groupi_n_1887;
  wire csa_tree_add_51_79_groupi_n_1888, csa_tree_add_51_79_groupi_n_1889, csa_tree_add_51_79_groupi_n_1890, csa_tree_add_51_79_groupi_n_1891, csa_tree_add_51_79_groupi_n_1892, csa_tree_add_51_79_groupi_n_1893, csa_tree_add_51_79_groupi_n_1894, csa_tree_add_51_79_groupi_n_1895;
  wire csa_tree_add_51_79_groupi_n_1896, csa_tree_add_51_79_groupi_n_1897, csa_tree_add_51_79_groupi_n_1898, csa_tree_add_51_79_groupi_n_1899, csa_tree_add_51_79_groupi_n_1900, csa_tree_add_51_79_groupi_n_1901, csa_tree_add_51_79_groupi_n_1902, csa_tree_add_51_79_groupi_n_1903;
  wire csa_tree_add_51_79_groupi_n_1904, csa_tree_add_51_79_groupi_n_1905, csa_tree_add_51_79_groupi_n_1906, csa_tree_add_51_79_groupi_n_1907, csa_tree_add_51_79_groupi_n_1908, csa_tree_add_51_79_groupi_n_1909, csa_tree_add_51_79_groupi_n_1910, csa_tree_add_51_79_groupi_n_1911;
  wire csa_tree_add_51_79_groupi_n_1912, csa_tree_add_51_79_groupi_n_1913, csa_tree_add_51_79_groupi_n_1914, csa_tree_add_51_79_groupi_n_1915, csa_tree_add_51_79_groupi_n_1916, csa_tree_add_51_79_groupi_n_1612, csa_tree_add_51_79_groupi_n_1918, csa_tree_add_51_79_groupi_n_1919;
  wire csa_tree_add_51_79_groupi_n_1920, csa_tree_add_51_79_groupi_n_1921, csa_tree_add_51_79_groupi_n_1922, csa_tree_add_51_79_groupi_n_1923, csa_tree_add_51_79_groupi_n_1924, csa_tree_add_51_79_groupi_n_1925, csa_tree_add_51_79_groupi_n_1926, csa_tree_add_51_79_groupi_n_1927;
  wire csa_tree_add_51_79_groupi_n_1928, csa_tree_add_51_79_groupi_n_1929, csa_tree_add_51_79_groupi_n_1930, csa_tree_add_51_79_groupi_n_1931, csa_tree_add_51_79_groupi_n_1932, csa_tree_add_51_79_groupi_n_1933, csa_tree_add_51_79_groupi_n_1934, csa_tree_add_51_79_groupi_n_1935;
  wire csa_tree_add_51_79_groupi_n_1936, csa_tree_add_51_79_groupi_n_1937, csa_tree_add_51_79_groupi_n_1938, csa_tree_add_51_79_groupi_n_1939, csa_tree_add_51_79_groupi_n_1940, csa_tree_add_51_79_groupi_n_1941, csa_tree_add_51_79_groupi_n_1942, csa_tree_add_51_79_groupi_n_1943;
  wire csa_tree_add_51_79_groupi_n_1944, csa_tree_add_51_79_groupi_n_1945, csa_tree_add_51_79_groupi_n_1946, csa_tree_add_51_79_groupi_n_1947, csa_tree_add_51_79_groupi_n_1948, csa_tree_add_51_79_groupi_n_1949, csa_tree_add_51_79_groupi_n_1950, csa_tree_add_51_79_groupi_n_1951;
  wire csa_tree_add_51_79_groupi_n_1952, csa_tree_add_51_79_groupi_n_1953, csa_tree_add_51_79_groupi_n_1954, csa_tree_add_51_79_groupi_n_1955, csa_tree_add_51_79_groupi_n_1956, csa_tree_add_51_79_groupi_n_1957, csa_tree_add_51_79_groupi_n_1958, csa_tree_add_51_79_groupi_n_1959;
  wire csa_tree_add_51_79_groupi_n_1960, csa_tree_add_51_79_groupi_n_1961, csa_tree_add_51_79_groupi_n_1962, csa_tree_add_51_79_groupi_n_1963, csa_tree_add_51_79_groupi_n_1964, csa_tree_add_51_79_groupi_n_1965, csa_tree_add_51_79_groupi_n_1966, csa_tree_add_51_79_groupi_n_1967;
  wire csa_tree_add_51_79_groupi_n_1968, csa_tree_add_51_79_groupi_n_1405, csa_tree_add_51_79_groupi_n_1970, csa_tree_add_51_79_groupi_n_1971, csa_tree_add_51_79_groupi_n_1411, csa_tree_add_51_79_groupi_n_1973, csa_tree_add_51_79_groupi_n_1974, csa_tree_add_51_79_groupi_n_1420;
  wire csa_tree_add_51_79_groupi_n_1976, csa_tree_add_51_79_groupi_n_1977, csa_tree_add_51_79_groupi_n_1240, csa_tree_add_51_79_groupi_n_1979, csa_tree_add_51_79_groupi_n_1243, csa_tree_add_51_79_groupi_n_1981, csa_tree_add_51_79_groupi_n_1246, csa_tree_add_51_79_groupi_n_1983;
  wire csa_tree_add_51_79_groupi_n_1231, csa_tree_add_51_79_groupi_n_1985, csa_tree_add_51_79_groupi_n_1252, csa_tree_add_51_79_groupi_n_1987, csa_tree_add_51_79_groupi_n_1255, csa_tree_add_51_79_groupi_n_1989, csa_tree_add_51_79_groupi_n_1237, csa_tree_add_51_79_groupi_n_1991;
  wire csa_tree_add_51_79_groupi_n_1258, csa_tree_add_51_79_groupi_n_1993, csa_tree_add_51_79_groupi_n_1444, csa_tree_add_51_79_groupi_n_1995, csa_tree_add_51_79_groupi_n_1996, csa_tree_add_51_79_groupi_n_1264, csa_tree_add_51_79_groupi_n_1998, csa_tree_add_51_79_groupi_n_1213;
  wire csa_tree_add_51_79_groupi_n_2000, csa_tree_add_51_79_groupi_n_1276, csa_tree_add_51_79_groupi_n_2002, csa_tree_add_51_79_groupi_n_2003, csa_tree_add_51_79_groupi_n_1282, csa_tree_add_51_79_groupi_n_2005, csa_tree_add_51_79_groupi_n_2006, csa_tree_add_51_79_groupi_n_1288;
  wire csa_tree_add_51_79_groupi_n_2008, csa_tree_add_51_79_groupi_n_2009, csa_tree_add_51_79_groupi_n_1294, csa_tree_add_51_79_groupi_n_2011, csa_tree_add_51_79_groupi_n_2012, csa_tree_add_51_79_groupi_n_1300, csa_tree_add_51_79_groupi_n_2014, csa_tree_add_51_79_groupi_n_2015;
  wire csa_tree_add_51_79_groupi_n_2016, csa_tree_add_51_79_groupi_n_2017, csa_tree_add_51_79_groupi_n_2018, csa_tree_add_51_79_groupi_n_2019, csa_tree_add_51_79_groupi_n_2020, csa_tree_add_51_79_groupi_n_2021, csa_tree_add_51_79_groupi_n_2022, csa_tree_add_51_79_groupi_n_2023;
  wire csa_tree_add_51_79_groupi_n_2024, csa_tree_add_51_79_groupi_n_2025, csa_tree_add_51_79_groupi_n_2026, csa_tree_add_51_79_groupi_n_2027, csa_tree_add_51_79_groupi_n_2028, csa_tree_add_51_79_groupi_n_2029, csa_tree_add_51_79_groupi_n_2030, csa_tree_add_51_79_groupi_n_2031;
  wire csa_tree_add_51_79_groupi_n_2032, csa_tree_add_51_79_groupi_n_2033, csa_tree_add_51_79_groupi_n_2034, csa_tree_add_51_79_groupi_n_2035, csa_tree_add_51_79_groupi_n_2036, csa_tree_add_51_79_groupi_n_2037, csa_tree_add_51_79_groupi_n_2038, csa_tree_add_51_79_groupi_n_2039;
  wire csa_tree_add_51_79_groupi_n_2040, csa_tree_add_51_79_groupi_n_2041, csa_tree_add_51_79_groupi_n_2042, csa_tree_add_51_79_groupi_n_2043, csa_tree_add_51_79_groupi_n_2044, csa_tree_add_51_79_groupi_n_2045, csa_tree_add_51_79_groupi_n_2046, csa_tree_add_51_79_groupi_n_2047;
  wire csa_tree_add_51_79_groupi_n_2048, csa_tree_add_51_79_groupi_n_2049, csa_tree_add_51_79_groupi_n_2050, csa_tree_add_51_79_groupi_n_2051, csa_tree_add_51_79_groupi_n_2052, csa_tree_add_51_79_groupi_n_2053, csa_tree_add_51_79_groupi_n_2054, csa_tree_add_51_79_groupi_n_2055;
  wire csa_tree_add_51_79_groupi_n_2056, csa_tree_add_51_79_groupi_n_2057, csa_tree_add_51_79_groupi_n_2058, csa_tree_add_51_79_groupi_n_2059, csa_tree_add_51_79_groupi_n_2060, csa_tree_add_51_79_groupi_n_2061, csa_tree_add_51_79_groupi_n_2062, csa_tree_add_51_79_groupi_n_2063;
  wire csa_tree_add_51_79_groupi_n_2064, csa_tree_add_51_79_groupi_n_2065, csa_tree_add_51_79_groupi_n_2066, csa_tree_add_51_79_groupi_n_2067, csa_tree_add_51_79_groupi_n_2068, csa_tree_add_51_79_groupi_n_2069, csa_tree_add_51_79_groupi_n_2070, csa_tree_add_51_79_groupi_n_2071;
  wire csa_tree_add_51_79_groupi_n_2072, csa_tree_add_51_79_groupi_n_2073, csa_tree_add_51_79_groupi_n_2074, csa_tree_add_51_79_groupi_n_2075, csa_tree_add_51_79_groupi_n_2076, csa_tree_add_51_79_groupi_n_2077, csa_tree_add_51_79_groupi_n_2078, csa_tree_add_51_79_groupi_n_2079;
  wire csa_tree_add_51_79_groupi_n_2080, csa_tree_add_51_79_groupi_n_2081, csa_tree_add_51_79_groupi_n_2082, csa_tree_add_51_79_groupi_n_2083, csa_tree_add_51_79_groupi_n_2084, csa_tree_add_51_79_groupi_n_2085, csa_tree_add_51_79_groupi_n_2086, csa_tree_add_51_79_groupi_n_2087;
  wire csa_tree_add_51_79_groupi_n_2088, csa_tree_add_51_79_groupi_n_2089, csa_tree_add_51_79_groupi_n_2090, csa_tree_add_51_79_groupi_n_2091, csa_tree_add_51_79_groupi_n_2092, csa_tree_add_51_79_groupi_n_2093, csa_tree_add_51_79_groupi_n_2094, csa_tree_add_51_79_groupi_n_2095;
  wire csa_tree_add_51_79_groupi_n_2096, csa_tree_add_51_79_groupi_n_2097, csa_tree_add_51_79_groupi_n_2098, csa_tree_add_51_79_groupi_n_2099, csa_tree_add_51_79_groupi_n_2100, csa_tree_add_51_79_groupi_n_2101, csa_tree_add_51_79_groupi_n_2102, csa_tree_add_51_79_groupi_n_2103;
  wire csa_tree_add_51_79_groupi_n_2104, csa_tree_add_51_79_groupi_n_2105, csa_tree_add_51_79_groupi_n_2106, csa_tree_add_51_79_groupi_n_2107, csa_tree_add_51_79_groupi_n_2108, csa_tree_add_51_79_groupi_n_2109, csa_tree_add_51_79_groupi_n_2110, csa_tree_add_51_79_groupi_n_2111;
  wire csa_tree_add_51_79_groupi_n_2112, csa_tree_add_51_79_groupi_n_2113, csa_tree_add_51_79_groupi_n_2114, csa_tree_add_51_79_groupi_n_2115, csa_tree_add_51_79_groupi_n_2116, csa_tree_add_51_79_groupi_n_2117, csa_tree_add_51_79_groupi_n_2118, csa_tree_add_51_79_groupi_n_2119;
  wire csa_tree_add_51_79_groupi_n_2120, csa_tree_add_51_79_groupi_n_2121, csa_tree_add_51_79_groupi_n_2122, csa_tree_add_51_79_groupi_n_2123, csa_tree_add_51_79_groupi_n_2124, csa_tree_add_51_79_groupi_n_2125, csa_tree_add_51_79_groupi_n_2126, csa_tree_add_51_79_groupi_n_2127;
  wire csa_tree_add_51_79_groupi_n_2128, csa_tree_add_51_79_groupi_n_2129, csa_tree_add_51_79_groupi_n_2130, csa_tree_add_51_79_groupi_n_2131, csa_tree_add_51_79_groupi_n_2132, csa_tree_add_51_79_groupi_n_2133, csa_tree_add_51_79_groupi_n_2134, csa_tree_add_51_79_groupi_n_2135;
  wire csa_tree_add_51_79_groupi_n_2136, csa_tree_add_51_79_groupi_n_2137, csa_tree_add_51_79_groupi_n_2138, csa_tree_add_51_79_groupi_n_2139, csa_tree_add_51_79_groupi_n_2140, csa_tree_add_51_79_groupi_n_2141, csa_tree_add_51_79_groupi_n_2142, csa_tree_add_51_79_groupi_n_2143;
  wire csa_tree_add_51_79_groupi_n_2144, csa_tree_add_51_79_groupi_n_2145, csa_tree_add_51_79_groupi_n_2146, csa_tree_add_51_79_groupi_n_2147, csa_tree_add_51_79_groupi_n_2148, csa_tree_add_51_79_groupi_n_2149, csa_tree_add_51_79_groupi_n_2150, csa_tree_add_51_79_groupi_n_2151;
  wire csa_tree_add_51_79_groupi_n_2152, csa_tree_add_51_79_groupi_n_2153, csa_tree_add_51_79_groupi_n_2154, csa_tree_add_51_79_groupi_n_2155, csa_tree_add_51_79_groupi_n_2156, csa_tree_add_51_79_groupi_n_2157, csa_tree_add_51_79_groupi_n_2158, csa_tree_add_51_79_groupi_n_2159;
  wire csa_tree_add_51_79_groupi_n_2160, csa_tree_add_51_79_groupi_n_2161, csa_tree_add_51_79_groupi_n_2162, csa_tree_add_51_79_groupi_n_2163, csa_tree_add_51_79_groupi_n_2164, csa_tree_add_51_79_groupi_n_2165, csa_tree_add_51_79_groupi_n_2166, csa_tree_add_51_79_groupi_n_2167;
  wire csa_tree_add_51_79_groupi_n_2168, csa_tree_add_51_79_groupi_n_2169, csa_tree_add_51_79_groupi_n_2170, csa_tree_add_51_79_groupi_n_2171, csa_tree_add_51_79_groupi_n_2172, csa_tree_add_51_79_groupi_n_2173, csa_tree_add_51_79_groupi_n_2174, csa_tree_add_51_79_groupi_n_2175;
  wire csa_tree_add_51_79_groupi_n_2176, csa_tree_add_51_79_groupi_n_2177, csa_tree_add_51_79_groupi_n_2178, csa_tree_add_51_79_groupi_n_2179, csa_tree_add_51_79_groupi_n_2180, csa_tree_add_51_79_groupi_n_2181, csa_tree_add_51_79_groupi_n_2182, csa_tree_add_51_79_groupi_n_2183;
  wire csa_tree_add_51_79_groupi_n_2184, csa_tree_add_51_79_groupi_n_2185, csa_tree_add_51_79_groupi_n_2186, csa_tree_add_51_79_groupi_n_2187, csa_tree_add_51_79_groupi_n_2188, csa_tree_add_51_79_groupi_n_2189, csa_tree_add_51_79_groupi_n_2190, csa_tree_add_51_79_groupi_n_2191;
  wire csa_tree_add_51_79_groupi_n_2192, csa_tree_add_51_79_groupi_n_2193, csa_tree_add_51_79_groupi_n_2194, csa_tree_add_51_79_groupi_n_2195, csa_tree_add_51_79_groupi_n_2196, csa_tree_add_51_79_groupi_n_2197, csa_tree_add_51_79_groupi_n_2198, csa_tree_add_51_79_groupi_n_2199;
  wire csa_tree_add_51_79_groupi_n_2200, csa_tree_add_51_79_groupi_n_2201, csa_tree_add_51_79_groupi_n_2202, csa_tree_add_51_79_groupi_n_2203, csa_tree_add_51_79_groupi_n_2204, csa_tree_add_51_79_groupi_n_2205, csa_tree_add_51_79_groupi_n_2206, csa_tree_add_51_79_groupi_n_2207;
  wire csa_tree_add_51_79_groupi_n_2208, csa_tree_add_51_79_groupi_n_2209, csa_tree_add_51_79_groupi_n_2210, csa_tree_add_51_79_groupi_n_2211, csa_tree_add_51_79_groupi_n_2212, csa_tree_add_51_79_groupi_n_2213, csa_tree_add_51_79_groupi_n_2214, csa_tree_add_51_79_groupi_n_2215;
  wire csa_tree_add_51_79_groupi_n_2216, csa_tree_add_51_79_groupi_n_2217, csa_tree_add_51_79_groupi_n_2218, csa_tree_add_51_79_groupi_n_2219, csa_tree_add_51_79_groupi_n_2220, csa_tree_add_51_79_groupi_n_2221, csa_tree_add_51_79_groupi_n_2222, csa_tree_add_51_79_groupi_n_2223;
  wire csa_tree_add_51_79_groupi_n_2224, csa_tree_add_51_79_groupi_n_2225, csa_tree_add_51_79_groupi_n_2226, csa_tree_add_51_79_groupi_n_2227, csa_tree_add_51_79_groupi_n_2228, csa_tree_add_51_79_groupi_n_2229, csa_tree_add_51_79_groupi_n_2230, csa_tree_add_51_79_groupi_n_2231;
  wire csa_tree_add_51_79_groupi_n_2232, csa_tree_add_51_79_groupi_n_2233, csa_tree_add_51_79_groupi_n_2234, csa_tree_add_51_79_groupi_n_2235, csa_tree_add_51_79_groupi_n_2236, csa_tree_add_51_79_groupi_n_2237, csa_tree_add_51_79_groupi_n_2238, csa_tree_add_51_79_groupi_n_2239;
  wire csa_tree_add_51_79_groupi_n_2240, csa_tree_add_51_79_groupi_n_2241, csa_tree_add_51_79_groupi_n_2242, csa_tree_add_51_79_groupi_n_2243, csa_tree_add_51_79_groupi_n_2244, csa_tree_add_51_79_groupi_n_2245, csa_tree_add_51_79_groupi_n_2246, csa_tree_add_51_79_groupi_n_2247;
  wire csa_tree_add_51_79_groupi_n_2248, csa_tree_add_51_79_groupi_n_2249, csa_tree_add_51_79_groupi_n_2250, csa_tree_add_51_79_groupi_n_2251, csa_tree_add_51_79_groupi_n_2252, csa_tree_add_51_79_groupi_n_2253, csa_tree_add_51_79_groupi_n_2254, csa_tree_add_51_79_groupi_n_2255;
  wire csa_tree_add_51_79_groupi_n_2256, csa_tree_add_51_79_groupi_n_2257, csa_tree_add_51_79_groupi_n_2258, csa_tree_add_51_79_groupi_n_2259, csa_tree_add_51_79_groupi_n_2260, csa_tree_add_51_79_groupi_n_2261, csa_tree_add_51_79_groupi_n_2262, csa_tree_add_51_79_groupi_n_2263;
  wire csa_tree_add_51_79_groupi_n_2264, csa_tree_add_51_79_groupi_n_2265, csa_tree_add_51_79_groupi_n_2266, csa_tree_add_51_79_groupi_n_2267, csa_tree_add_51_79_groupi_n_2268, csa_tree_add_51_79_groupi_n_2269, csa_tree_add_51_79_groupi_n_2270, csa_tree_add_51_79_groupi_n_2271;
  wire csa_tree_add_51_79_groupi_n_2272, csa_tree_add_51_79_groupi_n_2273, csa_tree_add_51_79_groupi_n_2274, csa_tree_add_51_79_groupi_n_2275, csa_tree_add_51_79_groupi_n_2276, csa_tree_add_51_79_groupi_n_2277, csa_tree_add_51_79_groupi_n_2278, csa_tree_add_51_79_groupi_n_2279;
  wire csa_tree_add_51_79_groupi_n_2280, csa_tree_add_51_79_groupi_n_2281, csa_tree_add_51_79_groupi_n_2282, csa_tree_add_51_79_groupi_n_2283, csa_tree_add_51_79_groupi_n_2284, csa_tree_add_51_79_groupi_n_2285, csa_tree_add_51_79_groupi_n_2286, csa_tree_add_51_79_groupi_n_2287;
  wire csa_tree_add_51_79_groupi_n_2288, csa_tree_add_51_79_groupi_n_2289, csa_tree_add_51_79_groupi_n_2290, csa_tree_add_51_79_groupi_n_2291, csa_tree_add_51_79_groupi_n_2292, csa_tree_add_51_79_groupi_n_2293, csa_tree_add_51_79_groupi_n_2294, csa_tree_add_51_79_groupi_n_2295;
  wire csa_tree_add_51_79_groupi_n_2296, csa_tree_add_51_79_groupi_n_2297, csa_tree_add_51_79_groupi_n_2298, csa_tree_add_51_79_groupi_n_2299, csa_tree_add_51_79_groupi_n_2300, csa_tree_add_51_79_groupi_n_2301, csa_tree_add_51_79_groupi_n_2302, csa_tree_add_51_79_groupi_n_2303;
  wire csa_tree_add_51_79_groupi_n_2304, csa_tree_add_51_79_groupi_n_2305, csa_tree_add_51_79_groupi_n_2306, csa_tree_add_51_79_groupi_n_2307, csa_tree_add_51_79_groupi_n_2308, csa_tree_add_51_79_groupi_n_2309, csa_tree_add_51_79_groupi_n_2310, csa_tree_add_51_79_groupi_n_2311;
  wire csa_tree_add_51_79_groupi_n_2312, csa_tree_add_51_79_groupi_n_2313, csa_tree_add_51_79_groupi_n_2314, csa_tree_add_51_79_groupi_n_2315, csa_tree_add_51_79_groupi_n_2316, csa_tree_add_51_79_groupi_n_2317, csa_tree_add_51_79_groupi_n_2318, csa_tree_add_51_79_groupi_n_2319;
  wire csa_tree_add_51_79_groupi_n_2320, csa_tree_add_51_79_groupi_n_2321, csa_tree_add_51_79_groupi_n_1542, csa_tree_add_51_79_groupi_n_2323, csa_tree_add_51_79_groupi_n_2324, csa_tree_add_51_79_groupi_n_2325, csa_tree_add_51_79_groupi_n_2326, csa_tree_add_51_79_groupi_n_2327;
  wire csa_tree_add_51_79_groupi_n_2328, csa_tree_add_51_79_groupi_n_2329, csa_tree_add_51_79_groupi_n_1601, csa_tree_add_51_79_groupi_n_2331, csa_tree_add_51_79_groupi_n_2332, csa_tree_add_51_79_groupi_n_2333, csa_tree_add_51_79_groupi_n_2334, csa_tree_add_51_79_groupi_n_2335;
  wire csa_tree_add_51_79_groupi_n_2336, csa_tree_add_51_79_groupi_n_2337, csa_tree_add_51_79_groupi_n_2338, csa_tree_add_51_79_groupi_n_2339, csa_tree_add_51_79_groupi_n_2340, csa_tree_add_51_79_groupi_n_1539, csa_tree_add_51_79_groupi_n_2342, csa_tree_add_51_79_groupi_n_1550;
  wire csa_tree_add_51_79_groupi_n_2344, csa_tree_add_51_79_groupi_n_2345, csa_tree_add_51_79_groupi_n_2346, csa_tree_add_51_79_groupi_n_2347, csa_tree_add_51_79_groupi_n_2348, csa_tree_add_51_79_groupi_n_2349, csa_tree_add_51_79_groupi_n_2350, csa_tree_add_51_79_groupi_n_1537;
  wire csa_tree_add_51_79_groupi_n_2352, csa_tree_add_51_79_groupi_n_2353, csa_tree_add_51_79_groupi_n_2354, csa_tree_add_51_79_groupi_n_2355, csa_tree_add_51_79_groupi_n_2356, csa_tree_add_51_79_groupi_n_1599, csa_tree_add_51_79_groupi_n_2358, csa_tree_add_51_79_groupi_n_2359;
  wire csa_tree_add_51_79_groupi_n_2360, csa_tree_add_51_79_groupi_n_1617, csa_tree_add_51_79_groupi_n_2362, csa_tree_add_51_79_groupi_n_2363, csa_tree_add_51_79_groupi_n_2364, csa_tree_add_51_79_groupi_n_2365, csa_tree_add_51_79_groupi_n_2366, csa_tree_add_51_79_groupi_n_2367;
  wire csa_tree_add_51_79_groupi_n_2368, csa_tree_add_51_79_groupi_n_2369, csa_tree_add_51_79_groupi_n_2370, csa_tree_add_51_79_groupi_n_2371, csa_tree_add_51_79_groupi_n_2372, csa_tree_add_51_79_groupi_n_2373, csa_tree_add_51_79_groupi_n_2374, csa_tree_add_51_79_groupi_n_2375;
  wire csa_tree_add_51_79_groupi_n_2376, csa_tree_add_51_79_groupi_n_2377, csa_tree_add_51_79_groupi_n_2378, csa_tree_add_51_79_groupi_n_2379, csa_tree_add_51_79_groupi_n_2380, csa_tree_add_51_79_groupi_n_2381, csa_tree_add_51_79_groupi_n_2382, csa_tree_add_51_79_groupi_n_2383;
  wire csa_tree_add_51_79_groupi_n_2384, csa_tree_add_51_79_groupi_n_2385, csa_tree_add_51_79_groupi_n_2386, csa_tree_add_51_79_groupi_n_2387, csa_tree_add_51_79_groupi_n_2388, csa_tree_add_51_79_groupi_n_2389, csa_tree_add_51_79_groupi_n_2390, csa_tree_add_51_79_groupi_n_2391;
  wire csa_tree_add_51_79_groupi_n_2392, csa_tree_add_51_79_groupi_n_2393, csa_tree_add_51_79_groupi_n_2394, csa_tree_add_51_79_groupi_n_2395, csa_tree_add_51_79_groupi_n_2396, csa_tree_add_51_79_groupi_n_2397, csa_tree_add_51_79_groupi_n_2398, csa_tree_add_51_79_groupi_n_1607;
  wire csa_tree_add_51_79_groupi_n_2400, csa_tree_add_51_79_groupi_n_2401, csa_tree_add_51_79_groupi_n_2402, csa_tree_add_51_79_groupi_n_2403, csa_tree_add_51_79_groupi_n_2404, csa_tree_add_51_79_groupi_n_2405, csa_tree_add_51_79_groupi_n_1610, csa_tree_add_51_79_groupi_n_2407;
  wire csa_tree_add_51_79_groupi_n_2408, csa_tree_add_51_79_groupi_n_2409, csa_tree_add_51_79_groupi_n_2410, csa_tree_add_51_79_groupi_n_2411, csa_tree_add_51_79_groupi_n_2412, csa_tree_add_51_79_groupi_n_2413, csa_tree_add_51_79_groupi_n_2414, csa_tree_add_51_79_groupi_n_2415;
  wire csa_tree_add_51_79_groupi_n_2416, csa_tree_add_51_79_groupi_n_2417, csa_tree_add_51_79_groupi_n_2418, csa_tree_add_51_79_groupi_n_1606, csa_tree_add_51_79_groupi_n_2420, csa_tree_add_51_79_groupi_n_2421, csa_tree_add_51_79_groupi_n_2422, csa_tree_add_51_79_groupi_n_2423;
  wire csa_tree_add_51_79_groupi_n_2424, csa_tree_add_51_79_groupi_n_2425, csa_tree_add_51_79_groupi_n_2426, csa_tree_add_51_79_groupi_n_2427, csa_tree_add_51_79_groupi_n_2428, csa_tree_add_51_79_groupi_n_2429, csa_tree_add_51_79_groupi_n_2430, csa_tree_add_51_79_groupi_n_2431;
  wire csa_tree_add_51_79_groupi_n_2432, csa_tree_add_51_79_groupi_n_2433, csa_tree_add_51_79_groupi_n_2434, csa_tree_add_51_79_groupi_n_1219, csa_tree_add_51_79_groupi_n_2436, csa_tree_add_51_79_groupi_n_1306, csa_tree_add_51_79_groupi_n_2438, csa_tree_add_51_79_groupi_n_2439;
  wire csa_tree_add_51_79_groupi_n_1312, csa_tree_add_51_79_groupi_n_2441, csa_tree_add_51_79_groupi_n_2442, csa_tree_add_51_79_groupi_n_1318, csa_tree_add_51_79_groupi_n_2444, csa_tree_add_51_79_groupi_n_2445, csa_tree_add_51_79_groupi_n_1222, csa_tree_add_51_79_groupi_n_2447;
  wire csa_tree_add_51_79_groupi_n_1324, csa_tree_add_51_79_groupi_n_2449, csa_tree_add_51_79_groupi_n_2450, csa_tree_add_51_79_groupi_n_1330, csa_tree_add_51_79_groupi_n_2452, csa_tree_add_51_79_groupi_n_2453, csa_tree_add_51_79_groupi_n_1225, csa_tree_add_51_79_groupi_n_2455;
  wire csa_tree_add_51_79_groupi_n_1336, csa_tree_add_51_79_groupi_n_2457, csa_tree_add_51_79_groupi_n_2458, csa_tree_add_51_79_groupi_n_1342, csa_tree_add_51_79_groupi_n_2460, csa_tree_add_51_79_groupi_n_2461, csa_tree_add_51_79_groupi_n_1348, csa_tree_add_51_79_groupi_n_2463;
  wire csa_tree_add_51_79_groupi_n_2464, csa_tree_add_51_79_groupi_n_1354, csa_tree_add_51_79_groupi_n_2466, csa_tree_add_51_79_groupi_n_2467, csa_tree_add_51_79_groupi_n_1360, csa_tree_add_51_79_groupi_n_2469, csa_tree_add_51_79_groupi_n_2470, csa_tree_add_51_79_groupi_n_1369;
  wire csa_tree_add_51_79_groupi_n_2472, csa_tree_add_51_79_groupi_n_2473, csa_tree_add_51_79_groupi_n_1375, csa_tree_add_51_79_groupi_n_2475, csa_tree_add_51_79_groupi_n_2476, csa_tree_add_51_79_groupi_n_1384, csa_tree_add_51_79_groupi_n_2478, csa_tree_add_51_79_groupi_n_2479;
  wire csa_tree_add_51_79_groupi_n_1228, csa_tree_add_51_79_groupi_n_2481, csa_tree_add_51_79_groupi_n_1390, csa_tree_add_51_79_groupi_n_2483, csa_tree_add_51_79_groupi_n_2484, csa_tree_add_51_79_groupi_n_1438, csa_tree_add_51_79_groupi_n_2486, csa_tree_add_51_79_groupi_n_2487;
  wire csa_tree_add_51_79_groupi_n_1234, csa_tree_add_51_79_groupi_n_2489, csa_tree_add_51_79_groupi_n_1366, csa_tree_add_51_79_groupi_n_2491, csa_tree_add_51_79_groupi_n_2492, csa_tree_add_51_79_groupi_n_1402, csa_tree_add_51_79_groupi_n_2494, csa_tree_add_51_79_groupi_n_2495;
  wire csa_tree_add_51_79_groupi_n_1417, csa_tree_add_51_79_groupi_n_2497, csa_tree_add_51_79_groupi_n_2498, csa_tree_add_51_79_groupi_n_1429, csa_tree_add_51_79_groupi_n_2500, csa_tree_add_51_79_groupi_n_2501, csa_tree_add_51_79_groupi_n_1249, csa_tree_add_51_79_groupi_n_2503;
  wire csa_tree_add_51_79_groupi_n_1393, csa_tree_add_51_79_groupi_n_2505, csa_tree_add_51_79_groupi_n_2506, csa_tree_add_51_79_groupi_n_1261, csa_tree_add_51_79_groupi_n_2508, csa_tree_add_51_79_groupi_n_1273, csa_tree_add_51_79_groupi_n_2510, csa_tree_add_51_79_groupi_n_2511;
  wire csa_tree_add_51_79_groupi_n_1216, csa_tree_add_51_79_groupi_n_2513, csa_tree_add_51_79_groupi_n_2514, csa_tree_add_51_79_groupi_n_2515, csa_tree_add_51_79_groupi_n_2516, csa_tree_add_51_79_groupi_n_1081, csa_tree_add_51_79_groupi_n_2518, csa_tree_add_51_79_groupi_n_2519;
  wire csa_tree_add_51_79_groupi_n_1079, csa_tree_add_51_79_groupi_n_2521, csa_tree_add_51_79_groupi_n_2522, csa_tree_add_51_79_groupi_n_2523, csa_tree_add_51_79_groupi_n_2524, csa_tree_add_51_79_groupi_n_2525, csa_tree_add_51_79_groupi_n_1083, csa_tree_add_51_79_groupi_n_2527;
  wire csa_tree_add_51_79_groupi_n_2528, csa_tree_add_51_79_groupi_n_2529, csa_tree_add_51_79_groupi_n_2530, csa_tree_add_51_79_groupi_n_2531, csa_tree_add_51_79_groupi_n_2532, csa_tree_add_51_79_groupi_n_2533, csa_tree_add_51_79_groupi_n_2534, csa_tree_add_51_79_groupi_n_2535;
  wire csa_tree_add_51_79_groupi_n_2536, csa_tree_add_51_79_groupi_n_2537, csa_tree_add_51_79_groupi_n_2538, csa_tree_add_51_79_groupi_n_2539, csa_tree_add_51_79_groupi_n_1085, csa_tree_add_51_79_groupi_n_2541, csa_tree_add_51_79_groupi_n_2542, csa_tree_add_51_79_groupi_n_2543;
  wire csa_tree_add_51_79_groupi_n_2544, csa_tree_add_51_79_groupi_n_2545, csa_tree_add_51_79_groupi_n_2546, csa_tree_add_51_79_groupi_n_2547, csa_tree_add_51_79_groupi_n_2548, csa_tree_add_51_79_groupi_n_2549, csa_tree_add_51_79_groupi_n_2550, csa_tree_add_51_79_groupi_n_2551;
  wire csa_tree_add_51_79_groupi_n_2552, csa_tree_add_51_79_groupi_n_2553, csa_tree_add_51_79_groupi_n_2554, csa_tree_add_51_79_groupi_n_2555, csa_tree_add_51_79_groupi_n_2556, csa_tree_add_51_79_groupi_n_2557, csa_tree_add_51_79_groupi_n_2558, csa_tree_add_51_79_groupi_n_2559;
  wire csa_tree_add_51_79_groupi_n_2560, csa_tree_add_51_79_groupi_n_2561, csa_tree_add_51_79_groupi_n_2562, csa_tree_add_51_79_groupi_n_2563, csa_tree_add_51_79_groupi_n_2564, csa_tree_add_51_79_groupi_n_2565, csa_tree_add_51_79_groupi_n_2566, csa_tree_add_51_79_groupi_n_2567;
  wire csa_tree_add_51_79_groupi_n_2568, csa_tree_add_51_79_groupi_n_2569, csa_tree_add_51_79_groupi_n_2570, csa_tree_add_51_79_groupi_n_2571, csa_tree_add_51_79_groupi_n_2572, csa_tree_add_51_79_groupi_n_2573, csa_tree_add_51_79_groupi_n_2574, csa_tree_add_51_79_groupi_n_2575;
  wire csa_tree_add_51_79_groupi_n_2576, csa_tree_add_51_79_groupi_n_2577, csa_tree_add_51_79_groupi_n_2578, csa_tree_add_51_79_groupi_n_2579, csa_tree_add_51_79_groupi_n_2580, csa_tree_add_51_79_groupi_n_2581, csa_tree_add_51_79_groupi_n_2582, csa_tree_add_51_79_groupi_n_2583;
  wire csa_tree_add_51_79_groupi_n_2584, csa_tree_add_51_79_groupi_n_2585, csa_tree_add_51_79_groupi_n_2586, csa_tree_add_51_79_groupi_n_2587, csa_tree_add_51_79_groupi_n_2588, csa_tree_add_51_79_groupi_n_2589, csa_tree_add_51_79_groupi_n_2590, csa_tree_add_51_79_groupi_n_2591;
  wire csa_tree_add_51_79_groupi_n_2592, csa_tree_add_51_79_groupi_n_2593, csa_tree_add_51_79_groupi_n_2594, csa_tree_add_51_79_groupi_n_2595, csa_tree_add_51_79_groupi_n_2596, csa_tree_add_51_79_groupi_n_2597, csa_tree_add_51_79_groupi_n_2598, csa_tree_add_51_79_groupi_n_2599;
  wire csa_tree_add_51_79_groupi_n_2600, csa_tree_add_51_79_groupi_n_2601, csa_tree_add_51_79_groupi_n_2602, csa_tree_add_51_79_groupi_n_2603, csa_tree_add_51_79_groupi_n_2604, csa_tree_add_51_79_groupi_n_2605, csa_tree_add_51_79_groupi_n_2606, csa_tree_add_51_79_groupi_n_2607;
  wire csa_tree_add_51_79_groupi_n_2608, csa_tree_add_51_79_groupi_n_2609, csa_tree_add_51_79_groupi_n_2610, csa_tree_add_51_79_groupi_n_2611, csa_tree_add_51_79_groupi_n_2612, csa_tree_add_51_79_groupi_n_2613, csa_tree_add_51_79_groupi_n_2614, csa_tree_add_51_79_groupi_n_2615;
  wire csa_tree_add_51_79_groupi_n_2616, csa_tree_add_51_79_groupi_n_2617, csa_tree_add_51_79_groupi_n_2618, csa_tree_add_51_79_groupi_n_2619, csa_tree_add_51_79_groupi_n_2620, csa_tree_add_51_79_groupi_n_2621, csa_tree_add_51_79_groupi_n_2622, csa_tree_add_51_79_groupi_n_2623;
  wire csa_tree_add_51_79_groupi_n_2624, csa_tree_add_51_79_groupi_n_2625, csa_tree_add_51_79_groupi_n_2626, csa_tree_add_51_79_groupi_n_2627, csa_tree_add_51_79_groupi_n_2628, csa_tree_add_51_79_groupi_n_2629, csa_tree_add_51_79_groupi_n_2630, csa_tree_add_51_79_groupi_n_2631;
  wire csa_tree_add_51_79_groupi_n_2632, csa_tree_add_51_79_groupi_n_2633, csa_tree_add_51_79_groupi_n_2634, csa_tree_add_51_79_groupi_n_2635, csa_tree_add_51_79_groupi_n_2636, csa_tree_add_51_79_groupi_n_2637, csa_tree_add_51_79_groupi_n_2638, csa_tree_add_51_79_groupi_n_2639;
  wire csa_tree_add_51_79_groupi_n_2640, csa_tree_add_51_79_groupi_n_2641, csa_tree_add_51_79_groupi_n_2642, csa_tree_add_51_79_groupi_n_2643, csa_tree_add_51_79_groupi_n_2644, csa_tree_add_51_79_groupi_n_2645, csa_tree_add_51_79_groupi_n_2646, csa_tree_add_51_79_groupi_n_2647;
  wire csa_tree_add_51_79_groupi_n_2648, csa_tree_add_51_79_groupi_n_2649, csa_tree_add_51_79_groupi_n_2650, csa_tree_add_51_79_groupi_n_2651, csa_tree_add_51_79_groupi_n_2652, csa_tree_add_51_79_groupi_n_2653, csa_tree_add_51_79_groupi_n_2654, csa_tree_add_51_79_groupi_n_2655;
  wire csa_tree_add_51_79_groupi_n_2656, csa_tree_add_51_79_groupi_n_2657, csa_tree_add_51_79_groupi_n_2658, csa_tree_add_51_79_groupi_n_2659, csa_tree_add_51_79_groupi_n_2660, csa_tree_add_51_79_groupi_n_2661, csa_tree_add_51_79_groupi_n_2662, csa_tree_add_51_79_groupi_n_2663;
  wire csa_tree_add_51_79_groupi_n_2664, csa_tree_add_51_79_groupi_n_2665, csa_tree_add_51_79_groupi_n_2666, csa_tree_add_51_79_groupi_n_2667, csa_tree_add_51_79_groupi_n_2668, csa_tree_add_51_79_groupi_n_2669, csa_tree_add_51_79_groupi_n_2670, csa_tree_add_51_79_groupi_n_2671;
  wire csa_tree_add_51_79_groupi_n_2672, csa_tree_add_51_79_groupi_n_2673, csa_tree_add_51_79_groupi_n_2674, csa_tree_add_51_79_groupi_n_2675, csa_tree_add_51_79_groupi_n_2676, csa_tree_add_51_79_groupi_n_2677, csa_tree_add_51_79_groupi_n_2678, csa_tree_add_51_79_groupi_n_2679;
  wire csa_tree_add_51_79_groupi_n_2680, csa_tree_add_51_79_groupi_n_2681, csa_tree_add_51_79_groupi_n_2682, csa_tree_add_51_79_groupi_n_2683, csa_tree_add_51_79_groupi_n_2684, csa_tree_add_51_79_groupi_n_2685, csa_tree_add_51_79_groupi_n_2686, csa_tree_add_51_79_groupi_n_2687;
  wire csa_tree_add_51_79_groupi_n_2688, csa_tree_add_51_79_groupi_n_2689, csa_tree_add_51_79_groupi_n_2690, csa_tree_add_51_79_groupi_n_2691, csa_tree_add_51_79_groupi_n_2692, csa_tree_add_51_79_groupi_n_2693, csa_tree_add_51_79_groupi_n_2694, csa_tree_add_51_79_groupi_n_2695;
  wire csa_tree_add_51_79_groupi_n_2696, csa_tree_add_51_79_groupi_n_2697, csa_tree_add_51_79_groupi_n_2698, csa_tree_add_51_79_groupi_n_2699, csa_tree_add_51_79_groupi_n_2700, csa_tree_add_51_79_groupi_n_2701, csa_tree_add_51_79_groupi_n_2702, csa_tree_add_51_79_groupi_n_2703;
  wire csa_tree_add_51_79_groupi_n_2704, csa_tree_add_51_79_groupi_n_2705, csa_tree_add_51_79_groupi_n_2706, csa_tree_add_51_79_groupi_n_2707, csa_tree_add_51_79_groupi_n_2708, csa_tree_add_51_79_groupi_n_2709, csa_tree_add_51_79_groupi_n_2710, csa_tree_add_51_79_groupi_n_2711;
  wire csa_tree_add_51_79_groupi_n_2712, csa_tree_add_51_79_groupi_n_2713, csa_tree_add_51_79_groupi_n_2714, csa_tree_add_51_79_groupi_n_2715, csa_tree_add_51_79_groupi_n_2716, csa_tree_add_51_79_groupi_n_2717, csa_tree_add_51_79_groupi_n_2718, csa_tree_add_51_79_groupi_n_2719;
  wire csa_tree_add_51_79_groupi_n_2720, csa_tree_add_51_79_groupi_n_2721, csa_tree_add_51_79_groupi_n_2722, csa_tree_add_51_79_groupi_n_2723, csa_tree_add_51_79_groupi_n_2724, csa_tree_add_51_79_groupi_n_2725, csa_tree_add_51_79_groupi_n_2726, csa_tree_add_51_79_groupi_n_2727;
  wire csa_tree_add_51_79_groupi_n_2728, csa_tree_add_51_79_groupi_n_2729, csa_tree_add_51_79_groupi_n_2730, csa_tree_add_51_79_groupi_n_2731, csa_tree_add_51_79_groupi_n_2732, csa_tree_add_51_79_groupi_n_2733, csa_tree_add_51_79_groupi_n_2734, csa_tree_add_51_79_groupi_n_2735;
  wire csa_tree_add_51_79_groupi_n_2736, csa_tree_add_51_79_groupi_n_2737, csa_tree_add_51_79_groupi_n_2738, csa_tree_add_51_79_groupi_n_2739, csa_tree_add_51_79_groupi_n_2740, csa_tree_add_51_79_groupi_n_2741, csa_tree_add_51_79_groupi_n_2742, csa_tree_add_51_79_groupi_n_2743;
  wire csa_tree_add_51_79_groupi_n_2744, csa_tree_add_51_79_groupi_n_2745, csa_tree_add_51_79_groupi_n_2746, csa_tree_add_51_79_groupi_n_2747, csa_tree_add_51_79_groupi_n_2748, csa_tree_add_51_79_groupi_n_2749, csa_tree_add_51_79_groupi_n_2750, csa_tree_add_51_79_groupi_n_2751;
  wire csa_tree_add_51_79_groupi_n_2752, csa_tree_add_51_79_groupi_n_2753, csa_tree_add_51_79_groupi_n_2754, csa_tree_add_51_79_groupi_n_2755, csa_tree_add_51_79_groupi_n_2756, csa_tree_add_51_79_groupi_n_2757, csa_tree_add_51_79_groupi_n_2758, csa_tree_add_51_79_groupi_n_2759;
  wire csa_tree_add_51_79_groupi_n_2760, csa_tree_add_51_79_groupi_n_2761, csa_tree_add_51_79_groupi_n_2762, csa_tree_add_51_79_groupi_n_2763, csa_tree_add_51_79_groupi_n_2764, csa_tree_add_51_79_groupi_n_2765, csa_tree_add_51_79_groupi_n_2766, csa_tree_add_51_79_groupi_n_2767;
  wire csa_tree_add_51_79_groupi_n_2768, csa_tree_add_51_79_groupi_n_2769, csa_tree_add_51_79_groupi_n_2770, csa_tree_add_51_79_groupi_n_2771, csa_tree_add_51_79_groupi_n_2772, csa_tree_add_51_79_groupi_n_2773, csa_tree_add_51_79_groupi_n_2774, csa_tree_add_51_79_groupi_n_2775;
  wire csa_tree_add_51_79_groupi_n_2776, csa_tree_add_51_79_groupi_n_2777, csa_tree_add_51_79_groupi_n_2778, csa_tree_add_51_79_groupi_n_2779, csa_tree_add_51_79_groupi_n_2780, csa_tree_add_51_79_groupi_n_2781, csa_tree_add_51_79_groupi_n_2782, csa_tree_add_51_79_groupi_n_2783;
  wire csa_tree_add_51_79_groupi_n_2784, csa_tree_add_51_79_groupi_n_2785, csa_tree_add_51_79_groupi_n_2786, csa_tree_add_51_79_groupi_n_2787, csa_tree_add_51_79_groupi_n_2788, csa_tree_add_51_79_groupi_n_2789, csa_tree_add_51_79_groupi_n_2790, csa_tree_add_51_79_groupi_n_2791;
  wire csa_tree_add_51_79_groupi_n_2792, csa_tree_add_51_79_groupi_n_2793, csa_tree_add_51_79_groupi_n_2794, csa_tree_add_51_79_groupi_n_2795, csa_tree_add_51_79_groupi_n_2796, csa_tree_add_51_79_groupi_n_2797, csa_tree_add_51_79_groupi_n_2798, csa_tree_add_51_79_groupi_n_2799;
  wire csa_tree_add_51_79_groupi_n_2800, csa_tree_add_51_79_groupi_n_2801, csa_tree_add_51_79_groupi_n_2802, csa_tree_add_51_79_groupi_n_2803, csa_tree_add_51_79_groupi_n_2804, csa_tree_add_51_79_groupi_n_2805, csa_tree_add_51_79_groupi_n_2806, csa_tree_add_51_79_groupi_n_2807;
  wire csa_tree_add_51_79_groupi_n_2808, csa_tree_add_51_79_groupi_n_2809, csa_tree_add_51_79_groupi_n_2810, csa_tree_add_51_79_groupi_n_2811, csa_tree_add_51_79_groupi_n_2812, csa_tree_add_51_79_groupi_n_2813, csa_tree_add_51_79_groupi_n_2814, csa_tree_add_51_79_groupi_n_2815;
  wire csa_tree_add_51_79_groupi_n_2816, csa_tree_add_51_79_groupi_n_2817, csa_tree_add_51_79_groupi_n_2818, csa_tree_add_51_79_groupi_n_2819, csa_tree_add_51_79_groupi_n_2820, csa_tree_add_51_79_groupi_n_2821, csa_tree_add_51_79_groupi_n_2822, csa_tree_add_51_79_groupi_n_2823;
  wire csa_tree_add_51_79_groupi_n_2824, csa_tree_add_51_79_groupi_n_2825, csa_tree_add_51_79_groupi_n_2826, csa_tree_add_51_79_groupi_n_2827, csa_tree_add_51_79_groupi_n_2828, csa_tree_add_51_79_groupi_n_2829, csa_tree_add_51_79_groupi_n_2830, csa_tree_add_51_79_groupi_n_2831;
  wire csa_tree_add_51_79_groupi_n_2832, csa_tree_add_51_79_groupi_n_2833, csa_tree_add_51_79_groupi_n_2834, csa_tree_add_51_79_groupi_n_2835, csa_tree_add_51_79_groupi_n_2836, csa_tree_add_51_79_groupi_n_2837, csa_tree_add_51_79_groupi_n_2838, csa_tree_add_51_79_groupi_n_2839;
  wire csa_tree_add_51_79_groupi_n_2840, csa_tree_add_51_79_groupi_n_2841, csa_tree_add_51_79_groupi_n_2842, csa_tree_add_51_79_groupi_n_2843, csa_tree_add_51_79_groupi_n_2844, csa_tree_add_51_79_groupi_n_2845, csa_tree_add_51_79_groupi_n_2846, csa_tree_add_51_79_groupi_n_2847;
  wire csa_tree_add_51_79_groupi_n_2848, csa_tree_add_51_79_groupi_n_2849, csa_tree_add_51_79_groupi_n_2850, csa_tree_add_51_79_groupi_n_2851, csa_tree_add_51_79_groupi_n_2852, csa_tree_add_51_79_groupi_n_2853, csa_tree_add_51_79_groupi_n_2854, csa_tree_add_51_79_groupi_n_2855;
  wire csa_tree_add_51_79_groupi_n_2856, csa_tree_add_51_79_groupi_n_2857, csa_tree_add_51_79_groupi_n_2858, csa_tree_add_51_79_groupi_n_2859, csa_tree_add_51_79_groupi_n_2860, csa_tree_add_51_79_groupi_n_2861, csa_tree_add_51_79_groupi_n_2862, csa_tree_add_51_79_groupi_n_2863;
  wire csa_tree_add_51_79_groupi_n_2864, csa_tree_add_51_79_groupi_n_2865, csa_tree_add_51_79_groupi_n_2866, csa_tree_add_51_79_groupi_n_2867, csa_tree_add_51_79_groupi_n_2868, csa_tree_add_51_79_groupi_n_2869, csa_tree_add_51_79_groupi_n_2870, csa_tree_add_51_79_groupi_n_2871;
  wire csa_tree_add_51_79_groupi_n_2872, csa_tree_add_51_79_groupi_n_2873, csa_tree_add_51_79_groupi_n_2874, csa_tree_add_51_79_groupi_n_2875, csa_tree_add_51_79_groupi_n_2876, csa_tree_add_51_79_groupi_n_2877, csa_tree_add_51_79_groupi_n_2878, csa_tree_add_51_79_groupi_n_2879;
  wire csa_tree_add_51_79_groupi_n_2880, csa_tree_add_51_79_groupi_n_2881, csa_tree_add_51_79_groupi_n_2882, csa_tree_add_51_79_groupi_n_2883, csa_tree_add_51_79_groupi_n_2884, csa_tree_add_51_79_groupi_n_2885, csa_tree_add_51_79_groupi_n_2886, csa_tree_add_51_79_groupi_n_2887;
  wire csa_tree_add_51_79_groupi_n_2888, csa_tree_add_51_79_groupi_n_2889, csa_tree_add_51_79_groupi_n_2890, csa_tree_add_51_79_groupi_n_2891, csa_tree_add_51_79_groupi_n_2892, csa_tree_add_51_79_groupi_n_2893, csa_tree_add_51_79_groupi_n_2894, csa_tree_add_51_79_groupi_n_2895;
  wire csa_tree_add_51_79_groupi_n_2896, csa_tree_add_51_79_groupi_n_2897, csa_tree_add_51_79_groupi_n_2898, csa_tree_add_51_79_groupi_n_2899, csa_tree_add_51_79_groupi_n_2900, csa_tree_add_51_79_groupi_n_2901, csa_tree_add_51_79_groupi_n_2902, csa_tree_add_51_79_groupi_n_2903;
  wire csa_tree_add_51_79_groupi_n_2904, csa_tree_add_51_79_groupi_n_2905, csa_tree_add_51_79_groupi_n_2906, csa_tree_add_51_79_groupi_n_2907, csa_tree_add_51_79_groupi_n_2908, csa_tree_add_51_79_groupi_n_2909, csa_tree_add_51_79_groupi_n_2910, csa_tree_add_51_79_groupi_n_2911;
  wire csa_tree_add_51_79_groupi_n_2912, csa_tree_add_51_79_groupi_n_2913, csa_tree_add_51_79_groupi_n_2914, csa_tree_add_51_79_groupi_n_2915, csa_tree_add_51_79_groupi_n_2916, csa_tree_add_51_79_groupi_n_2917, csa_tree_add_51_79_groupi_n_2918, csa_tree_add_51_79_groupi_n_2919;
  wire csa_tree_add_51_79_groupi_n_2920, csa_tree_add_51_79_groupi_n_2921, csa_tree_add_51_79_groupi_n_2922, csa_tree_add_51_79_groupi_n_2923, csa_tree_add_51_79_groupi_n_2924, csa_tree_add_51_79_groupi_n_2925, csa_tree_add_51_79_groupi_n_2926, csa_tree_add_51_79_groupi_n_2927;
  wire csa_tree_add_51_79_groupi_n_2928, csa_tree_add_51_79_groupi_n_2929, csa_tree_add_51_79_groupi_n_2930, csa_tree_add_51_79_groupi_n_2931, csa_tree_add_51_79_groupi_n_2932, csa_tree_add_51_79_groupi_n_2933, csa_tree_add_51_79_groupi_n_2934, csa_tree_add_51_79_groupi_n_2935;
  wire csa_tree_add_51_79_groupi_n_2936, csa_tree_add_51_79_groupi_n_2937, csa_tree_add_51_79_groupi_n_2938, csa_tree_add_51_79_groupi_n_2939, csa_tree_add_51_79_groupi_n_2940, csa_tree_add_51_79_groupi_n_2941, csa_tree_add_51_79_groupi_n_2942, csa_tree_add_51_79_groupi_n_2943;
  wire csa_tree_add_51_79_groupi_n_2944, csa_tree_add_51_79_groupi_n_2945, csa_tree_add_51_79_groupi_n_2946, csa_tree_add_51_79_groupi_n_2947, csa_tree_add_51_79_groupi_n_2948, csa_tree_add_51_79_groupi_n_2949, csa_tree_add_51_79_groupi_n_2950, csa_tree_add_51_79_groupi_n_2951;
  wire csa_tree_add_51_79_groupi_n_2952, csa_tree_add_51_79_groupi_n_2953, csa_tree_add_51_79_groupi_n_2954, csa_tree_add_51_79_groupi_n_2955, csa_tree_add_51_79_groupi_n_2956, csa_tree_add_51_79_groupi_n_2957, csa_tree_add_51_79_groupi_n_2958, csa_tree_add_51_79_groupi_n_2959;
  wire csa_tree_add_51_79_groupi_n_2960, csa_tree_add_51_79_groupi_n_2961, csa_tree_add_51_79_groupi_n_2962, csa_tree_add_51_79_groupi_n_2963, csa_tree_add_51_79_groupi_n_2964, csa_tree_add_51_79_groupi_n_2965, csa_tree_add_51_79_groupi_n_2966, csa_tree_add_51_79_groupi_n_2967;
  wire csa_tree_add_51_79_groupi_n_2968, csa_tree_add_51_79_groupi_n_2969, csa_tree_add_51_79_groupi_n_2970, csa_tree_add_51_79_groupi_n_2971, csa_tree_add_51_79_groupi_n_2972, csa_tree_add_51_79_groupi_n_2973, csa_tree_add_51_79_groupi_n_2974, csa_tree_add_51_79_groupi_n_2975;
  wire csa_tree_add_51_79_groupi_n_2976, csa_tree_add_51_79_groupi_n_2977, csa_tree_add_51_79_groupi_n_2978, csa_tree_add_51_79_groupi_n_2979, csa_tree_add_51_79_groupi_n_2980, csa_tree_add_51_79_groupi_n_2981, csa_tree_add_51_79_groupi_n_2982, csa_tree_add_51_79_groupi_n_2983;
  wire csa_tree_add_51_79_groupi_n_2984, csa_tree_add_51_79_groupi_n_2985, csa_tree_add_51_79_groupi_n_2986, csa_tree_add_51_79_groupi_n_2987, csa_tree_add_51_79_groupi_n_2988, csa_tree_add_51_79_groupi_n_2989, csa_tree_add_51_79_groupi_n_2990, csa_tree_add_51_79_groupi_n_2991;
  wire csa_tree_add_51_79_groupi_n_2992, csa_tree_add_51_79_groupi_n_2993, csa_tree_add_51_79_groupi_n_2994, csa_tree_add_51_79_groupi_n_2995, csa_tree_add_51_79_groupi_n_2996, csa_tree_add_51_79_groupi_n_2997, csa_tree_add_51_79_groupi_n_2998, csa_tree_add_51_79_groupi_n_2999;
  wire csa_tree_add_51_79_groupi_n_3000, csa_tree_add_51_79_groupi_n_3001, csa_tree_add_51_79_groupi_n_3002, csa_tree_add_51_79_groupi_n_3003, csa_tree_add_51_79_groupi_n_3004, csa_tree_add_51_79_groupi_n_3005, csa_tree_add_51_79_groupi_n_3006, csa_tree_add_51_79_groupi_n_3007;
  wire csa_tree_add_51_79_groupi_n_3008, csa_tree_add_51_79_groupi_n_3009, csa_tree_add_51_79_groupi_n_3010, csa_tree_add_51_79_groupi_n_3011, csa_tree_add_51_79_groupi_n_3012, csa_tree_add_51_79_groupi_n_3013, csa_tree_add_51_79_groupi_n_3014, csa_tree_add_51_79_groupi_n_3015;
  wire csa_tree_add_51_79_groupi_n_3016, csa_tree_add_51_79_groupi_n_3017, csa_tree_add_51_79_groupi_n_3018, csa_tree_add_51_79_groupi_n_3019, csa_tree_add_51_79_groupi_n_3020, csa_tree_add_51_79_groupi_n_3021, csa_tree_add_51_79_groupi_n_3022, csa_tree_add_51_79_groupi_n_3023;
  wire csa_tree_add_51_79_groupi_n_3024, csa_tree_add_51_79_groupi_n_3025, csa_tree_add_51_79_groupi_n_3026, csa_tree_add_51_79_groupi_n_3027, csa_tree_add_51_79_groupi_n_3028, csa_tree_add_51_79_groupi_n_3029, csa_tree_add_51_79_groupi_n_3030, csa_tree_add_51_79_groupi_n_3031;
  wire csa_tree_add_51_79_groupi_n_3032, csa_tree_add_51_79_groupi_n_3033, csa_tree_add_51_79_groupi_n_3034, csa_tree_add_51_79_groupi_n_3035, csa_tree_add_51_79_groupi_n_3036, csa_tree_add_51_79_groupi_n_3037, csa_tree_add_51_79_groupi_n_3038, csa_tree_add_51_79_groupi_n_3039;
  wire csa_tree_add_51_79_groupi_n_3040, csa_tree_add_51_79_groupi_n_3041, csa_tree_add_51_79_groupi_n_3042, csa_tree_add_51_79_groupi_n_3043, csa_tree_add_51_79_groupi_n_3044, csa_tree_add_51_79_groupi_n_3045, csa_tree_add_51_79_groupi_n_3046, csa_tree_add_51_79_groupi_n_3047;
  wire csa_tree_add_51_79_groupi_n_3048, csa_tree_add_51_79_groupi_n_3049, csa_tree_add_51_79_groupi_n_3050, csa_tree_add_51_79_groupi_n_3051, csa_tree_add_51_79_groupi_n_3052, csa_tree_add_51_79_groupi_n_3053, csa_tree_add_51_79_groupi_n_3054, csa_tree_add_51_79_groupi_n_3055;
  wire csa_tree_add_51_79_groupi_n_3056, csa_tree_add_51_79_groupi_n_3057, csa_tree_add_51_79_groupi_n_3058, csa_tree_add_51_79_groupi_n_3059, csa_tree_add_51_79_groupi_n_3060, csa_tree_add_51_79_groupi_n_3061, csa_tree_add_51_79_groupi_n_3062, csa_tree_add_51_79_groupi_n_3063;
  wire csa_tree_add_51_79_groupi_n_3064, csa_tree_add_51_79_groupi_n_3065, csa_tree_add_51_79_groupi_n_3066, csa_tree_add_51_79_groupi_n_3067, csa_tree_add_51_79_groupi_n_3068, csa_tree_add_51_79_groupi_n_3069, csa_tree_add_51_79_groupi_n_3070, csa_tree_add_51_79_groupi_n_3071;
  wire csa_tree_add_51_79_groupi_n_3072, csa_tree_add_51_79_groupi_n_3073, csa_tree_add_51_79_groupi_n_3074, csa_tree_add_51_79_groupi_n_3075, csa_tree_add_51_79_groupi_n_3076, csa_tree_add_51_79_groupi_n_3077, csa_tree_add_51_79_groupi_n_3078, csa_tree_add_51_79_groupi_n_3079;
  wire csa_tree_add_51_79_groupi_n_3080, csa_tree_add_51_79_groupi_n_3081, csa_tree_add_51_79_groupi_n_3082, csa_tree_add_51_79_groupi_n_3083, csa_tree_add_51_79_groupi_n_3084, csa_tree_add_51_79_groupi_n_3085, csa_tree_add_51_79_groupi_n_3086, csa_tree_add_51_79_groupi_n_3087;
  wire csa_tree_add_51_79_groupi_n_3088, csa_tree_add_51_79_groupi_n_3089, csa_tree_add_51_79_groupi_n_3090, csa_tree_add_51_79_groupi_n_3091, csa_tree_add_51_79_groupi_n_3092, csa_tree_add_51_79_groupi_n_3093, csa_tree_add_51_79_groupi_n_3094, csa_tree_add_51_79_groupi_n_3095;
  wire csa_tree_add_51_79_groupi_n_3096, csa_tree_add_51_79_groupi_n_3097, csa_tree_add_51_79_groupi_n_3098, csa_tree_add_51_79_groupi_n_3099, csa_tree_add_51_79_groupi_n_3100, csa_tree_add_51_79_groupi_n_3101, csa_tree_add_51_79_groupi_n_3102, csa_tree_add_51_79_groupi_n_3103;
  wire csa_tree_add_51_79_groupi_n_3104, csa_tree_add_51_79_groupi_n_3105, csa_tree_add_51_79_groupi_n_3106, csa_tree_add_51_79_groupi_n_3107, csa_tree_add_51_79_groupi_n_3108, csa_tree_add_51_79_groupi_n_3109, csa_tree_add_51_79_groupi_n_3110, csa_tree_add_51_79_groupi_n_3111;
  wire csa_tree_add_51_79_groupi_n_3112, csa_tree_add_51_79_groupi_n_3113, csa_tree_add_51_79_groupi_n_3114, csa_tree_add_51_79_groupi_n_3115, csa_tree_add_51_79_groupi_n_3116, csa_tree_add_51_79_groupi_n_3117, csa_tree_add_51_79_groupi_n_3118, csa_tree_add_51_79_groupi_n_3119;
  wire csa_tree_add_51_79_groupi_n_3120, csa_tree_add_51_79_groupi_n_3121, csa_tree_add_51_79_groupi_n_3122, csa_tree_add_51_79_groupi_n_3123, csa_tree_add_51_79_groupi_n_3124, csa_tree_add_51_79_groupi_n_3125, csa_tree_add_51_79_groupi_n_3126, csa_tree_add_51_79_groupi_n_3127;
  wire csa_tree_add_51_79_groupi_n_3128, csa_tree_add_51_79_groupi_n_3129, csa_tree_add_51_79_groupi_n_3130, csa_tree_add_51_79_groupi_n_3131, csa_tree_add_51_79_groupi_n_3132, csa_tree_add_51_79_groupi_n_3133, csa_tree_add_51_79_groupi_n_3134, csa_tree_add_51_79_groupi_n_3135;
  wire csa_tree_add_51_79_groupi_n_3136, csa_tree_add_51_79_groupi_n_3137, csa_tree_add_51_79_groupi_n_3138, csa_tree_add_51_79_groupi_n_3139, csa_tree_add_51_79_groupi_n_3140, csa_tree_add_51_79_groupi_n_3141, csa_tree_add_51_79_groupi_n_3142, csa_tree_add_51_79_groupi_n_3143;
  wire csa_tree_add_51_79_groupi_n_3144, csa_tree_add_51_79_groupi_n_3145, csa_tree_add_51_79_groupi_n_3146, csa_tree_add_51_79_groupi_n_3147, csa_tree_add_51_79_groupi_n_3148, csa_tree_add_51_79_groupi_n_3149, csa_tree_add_51_79_groupi_n_3150, csa_tree_add_51_79_groupi_n_3151;
  wire csa_tree_add_51_79_groupi_n_3152, csa_tree_add_51_79_groupi_n_3153, csa_tree_add_51_79_groupi_n_3154, csa_tree_add_51_79_groupi_n_3155, csa_tree_add_51_79_groupi_n_3156, csa_tree_add_51_79_groupi_n_3157, csa_tree_add_51_79_groupi_n_3158, csa_tree_add_51_79_groupi_n_3159;
  wire csa_tree_add_51_79_groupi_n_3160, csa_tree_add_51_79_groupi_n_3161, csa_tree_add_51_79_groupi_n_3162, csa_tree_add_51_79_groupi_n_3163, csa_tree_add_51_79_groupi_n_3164, csa_tree_add_51_79_groupi_n_3165, csa_tree_add_51_79_groupi_n_3166, csa_tree_add_51_79_groupi_n_3167;
  wire csa_tree_add_51_79_groupi_n_3168, csa_tree_add_51_79_groupi_n_3169, csa_tree_add_51_79_groupi_n_3170, csa_tree_add_51_79_groupi_n_3171, csa_tree_add_51_79_groupi_n_3172, csa_tree_add_51_79_groupi_n_3173, csa_tree_add_51_79_groupi_n_3174, csa_tree_add_51_79_groupi_n_3175;
  wire csa_tree_add_51_79_groupi_n_3176, csa_tree_add_51_79_groupi_n_3177, csa_tree_add_51_79_groupi_n_3178, csa_tree_add_51_79_groupi_n_3179, csa_tree_add_51_79_groupi_n_3180, csa_tree_add_51_79_groupi_n_3181, csa_tree_add_51_79_groupi_n_3182, csa_tree_add_51_79_groupi_n_3183;
  wire csa_tree_add_51_79_groupi_n_3184, csa_tree_add_51_79_groupi_n_3185, csa_tree_add_51_79_groupi_n_3186, csa_tree_add_51_79_groupi_n_3187, csa_tree_add_51_79_groupi_n_3188, csa_tree_add_51_79_groupi_n_3189, csa_tree_add_51_79_groupi_n_3190, csa_tree_add_51_79_groupi_n_3191;
  wire csa_tree_add_51_79_groupi_n_3192, csa_tree_add_51_79_groupi_n_3193, csa_tree_add_51_79_groupi_n_3194, csa_tree_add_51_79_groupi_n_3195, csa_tree_add_51_79_groupi_n_3196, csa_tree_add_51_79_groupi_n_3197, csa_tree_add_51_79_groupi_n_3198, csa_tree_add_51_79_groupi_n_3199;
  wire csa_tree_add_51_79_groupi_n_3200, csa_tree_add_51_79_groupi_n_3201, csa_tree_add_51_79_groupi_n_3202, csa_tree_add_51_79_groupi_n_3203, csa_tree_add_51_79_groupi_n_3204, csa_tree_add_51_79_groupi_n_3205, csa_tree_add_51_79_groupi_n_3206, csa_tree_add_51_79_groupi_n_3207;
  wire csa_tree_add_51_79_groupi_n_3208, csa_tree_add_51_79_groupi_n_3209, csa_tree_add_51_79_groupi_n_3210, csa_tree_add_51_79_groupi_n_3211, csa_tree_add_51_79_groupi_n_3212, csa_tree_add_51_79_groupi_n_3213, csa_tree_add_51_79_groupi_n_3214, csa_tree_add_51_79_groupi_n_3215;
  wire csa_tree_add_51_79_groupi_n_3216, csa_tree_add_51_79_groupi_n_3217, csa_tree_add_51_79_groupi_n_3218, csa_tree_add_51_79_groupi_n_3219, csa_tree_add_51_79_groupi_n_3220, csa_tree_add_51_79_groupi_n_3221, csa_tree_add_51_79_groupi_n_3222, csa_tree_add_51_79_groupi_n_3223;
  wire csa_tree_add_51_79_groupi_n_3224, csa_tree_add_51_79_groupi_n_3225, csa_tree_add_51_79_groupi_n_3226, csa_tree_add_51_79_groupi_n_3227, csa_tree_add_51_79_groupi_n_3228, csa_tree_add_51_79_groupi_n_3229, csa_tree_add_51_79_groupi_n_3230, csa_tree_add_51_79_groupi_n_3231;
  wire csa_tree_add_51_79_groupi_n_3232, csa_tree_add_51_79_groupi_n_3233, csa_tree_add_51_79_groupi_n_3234, csa_tree_add_51_79_groupi_n_3235, csa_tree_add_51_79_groupi_n_3236, csa_tree_add_51_79_groupi_n_3237, csa_tree_add_51_79_groupi_n_3238, csa_tree_add_51_79_groupi_n_3239;
  wire csa_tree_add_51_79_groupi_n_3240, csa_tree_add_51_79_groupi_n_3241, csa_tree_add_51_79_groupi_n_3242, csa_tree_add_51_79_groupi_n_3243, csa_tree_add_51_79_groupi_n_3244, csa_tree_add_51_79_groupi_n_3245, csa_tree_add_51_79_groupi_n_3246, csa_tree_add_51_79_groupi_n_3247;
  wire csa_tree_add_51_79_groupi_n_3248, csa_tree_add_51_79_groupi_n_3249, csa_tree_add_51_79_groupi_n_3250, csa_tree_add_51_79_groupi_n_3251, csa_tree_add_51_79_groupi_n_3252, csa_tree_add_51_79_groupi_n_3253, csa_tree_add_51_79_groupi_n_3254, csa_tree_add_51_79_groupi_n_3255;
  wire csa_tree_add_51_79_groupi_n_3256, csa_tree_add_51_79_groupi_n_3257, csa_tree_add_51_79_groupi_n_3258, csa_tree_add_51_79_groupi_n_3259, csa_tree_add_51_79_groupi_n_3260, csa_tree_add_51_79_groupi_n_3261, csa_tree_add_51_79_groupi_n_3262, csa_tree_add_51_79_groupi_n_3263;
  wire csa_tree_add_51_79_groupi_n_3264, csa_tree_add_51_79_groupi_n_3265, csa_tree_add_51_79_groupi_n_3266, csa_tree_add_51_79_groupi_n_3267, csa_tree_add_51_79_groupi_n_3268, csa_tree_add_51_79_groupi_n_3269, csa_tree_add_51_79_groupi_n_3270, csa_tree_add_51_79_groupi_n_3271;
  wire csa_tree_add_51_79_groupi_n_3272, csa_tree_add_51_79_groupi_n_3273, csa_tree_add_51_79_groupi_n_3274, csa_tree_add_51_79_groupi_n_3275, csa_tree_add_51_79_groupi_n_3276, csa_tree_add_51_79_groupi_n_3277, csa_tree_add_51_79_groupi_n_3278, csa_tree_add_51_79_groupi_n_3279;
  wire csa_tree_add_51_79_groupi_n_3280, csa_tree_add_51_79_groupi_n_3281, csa_tree_add_51_79_groupi_n_3282, csa_tree_add_51_79_groupi_n_3283, csa_tree_add_51_79_groupi_n_3284, csa_tree_add_51_79_groupi_n_3285, csa_tree_add_51_79_groupi_n_3286, csa_tree_add_51_79_groupi_n_3287;
  wire csa_tree_add_51_79_groupi_n_3288, csa_tree_add_51_79_groupi_n_3289, csa_tree_add_51_79_groupi_n_3290, csa_tree_add_51_79_groupi_n_3291, csa_tree_add_51_79_groupi_n_3292, csa_tree_add_51_79_groupi_n_3293, csa_tree_add_51_79_groupi_n_3294, csa_tree_add_51_79_groupi_n_3295;
  wire csa_tree_add_51_79_groupi_n_3296, csa_tree_add_51_79_groupi_n_3297, csa_tree_add_51_79_groupi_n_3298, csa_tree_add_51_79_groupi_n_3299, csa_tree_add_51_79_groupi_n_3300, csa_tree_add_51_79_groupi_n_3301, csa_tree_add_51_79_groupi_n_3302, csa_tree_add_51_79_groupi_n_3303;
  wire csa_tree_add_51_79_groupi_n_3304, csa_tree_add_51_79_groupi_n_3305, csa_tree_add_51_79_groupi_n_3306, csa_tree_add_51_79_groupi_n_3307, csa_tree_add_51_79_groupi_n_3308, csa_tree_add_51_79_groupi_n_3309, csa_tree_add_51_79_groupi_n_3310, csa_tree_add_51_79_groupi_n_3311;
  wire csa_tree_add_51_79_groupi_n_3312, csa_tree_add_51_79_groupi_n_3313, csa_tree_add_51_79_groupi_n_3314, csa_tree_add_51_79_groupi_n_3315, csa_tree_add_51_79_groupi_n_3316, csa_tree_add_51_79_groupi_n_3317, csa_tree_add_51_79_groupi_n_3318, csa_tree_add_51_79_groupi_n_3319;
  wire csa_tree_add_51_79_groupi_n_3320, csa_tree_add_51_79_groupi_n_3321, csa_tree_add_51_79_groupi_n_3322, csa_tree_add_51_79_groupi_n_3323, csa_tree_add_51_79_groupi_n_3324, csa_tree_add_51_79_groupi_n_3325, csa_tree_add_51_79_groupi_n_3326, csa_tree_add_51_79_groupi_n_3327;
  wire csa_tree_add_51_79_groupi_n_3328, csa_tree_add_51_79_groupi_n_3329, csa_tree_add_51_79_groupi_n_3330, csa_tree_add_51_79_groupi_n_3331, csa_tree_add_51_79_groupi_n_3332, csa_tree_add_51_79_groupi_n_3333, csa_tree_add_51_79_groupi_n_3334, csa_tree_add_51_79_groupi_n_3335;
  wire csa_tree_add_51_79_groupi_n_3336, csa_tree_add_51_79_groupi_n_3337, csa_tree_add_51_79_groupi_n_3338, csa_tree_add_51_79_groupi_n_3339, csa_tree_add_51_79_groupi_n_3340, csa_tree_add_51_79_groupi_n_3341, csa_tree_add_51_79_groupi_n_3342, csa_tree_add_51_79_groupi_n_3343;
  wire csa_tree_add_51_79_groupi_n_3344, csa_tree_add_51_79_groupi_n_3345, csa_tree_add_51_79_groupi_n_3346, csa_tree_add_51_79_groupi_n_3347, csa_tree_add_51_79_groupi_n_3348, csa_tree_add_51_79_groupi_n_3349, csa_tree_add_51_79_groupi_n_3350, csa_tree_add_51_79_groupi_n_3351;
  wire csa_tree_add_51_79_groupi_n_3352, csa_tree_add_51_79_groupi_n_3353, csa_tree_add_51_79_groupi_n_3354, csa_tree_add_51_79_groupi_n_3355, csa_tree_add_51_79_groupi_n_3356, csa_tree_add_51_79_groupi_n_3357, csa_tree_add_51_79_groupi_n_3358, csa_tree_add_51_79_groupi_n_3359;
  wire csa_tree_add_51_79_groupi_n_3360, csa_tree_add_51_79_groupi_n_3361, csa_tree_add_51_79_groupi_n_3362, csa_tree_add_51_79_groupi_n_3363, csa_tree_add_51_79_groupi_n_3364, csa_tree_add_51_79_groupi_n_3365, csa_tree_add_51_79_groupi_n_3366, csa_tree_add_51_79_groupi_n_3367;
  wire csa_tree_add_51_79_groupi_n_3368, csa_tree_add_51_79_groupi_n_3369, csa_tree_add_51_79_groupi_n_3370, csa_tree_add_51_79_groupi_n_3371, csa_tree_add_51_79_groupi_n_3372, csa_tree_add_51_79_groupi_n_3373, csa_tree_add_51_79_groupi_n_3374, csa_tree_add_51_79_groupi_n_3375;
  wire csa_tree_add_51_79_groupi_n_3376, csa_tree_add_51_79_groupi_n_3377, csa_tree_add_51_79_groupi_n_3378, csa_tree_add_51_79_groupi_n_3379, csa_tree_add_51_79_groupi_n_3380, csa_tree_add_51_79_groupi_n_3381, csa_tree_add_51_79_groupi_n_3382, csa_tree_add_51_79_groupi_n_3383;
  wire csa_tree_add_51_79_groupi_n_3384, csa_tree_add_51_79_groupi_n_3385, csa_tree_add_51_79_groupi_n_3386, csa_tree_add_51_79_groupi_n_3387, csa_tree_add_51_79_groupi_n_3388, csa_tree_add_51_79_groupi_n_3389, csa_tree_add_51_79_groupi_n_3390, csa_tree_add_51_79_groupi_n_3391;
  wire csa_tree_add_51_79_groupi_n_3392, csa_tree_add_51_79_groupi_n_3393, csa_tree_add_51_79_groupi_n_3394, csa_tree_add_51_79_groupi_n_3395, csa_tree_add_51_79_groupi_n_3396, csa_tree_add_51_79_groupi_n_3397, csa_tree_add_51_79_groupi_n_3398, csa_tree_add_51_79_groupi_n_3399;
  wire csa_tree_add_51_79_groupi_n_3400, csa_tree_add_51_79_groupi_n_3401, csa_tree_add_51_79_groupi_n_3402, csa_tree_add_51_79_groupi_n_3403, csa_tree_add_51_79_groupi_n_3404, csa_tree_add_51_79_groupi_n_3405, csa_tree_add_51_79_groupi_n_3406, csa_tree_add_51_79_groupi_n_3407;
  wire csa_tree_add_51_79_groupi_n_3408, csa_tree_add_51_79_groupi_n_3409, csa_tree_add_51_79_groupi_n_3410, csa_tree_add_51_79_groupi_n_3411, csa_tree_add_51_79_groupi_n_3412, csa_tree_add_51_79_groupi_n_3413, csa_tree_add_51_79_groupi_n_3414, csa_tree_add_51_79_groupi_n_3415;
  wire csa_tree_add_51_79_groupi_n_3416, csa_tree_add_51_79_groupi_n_3417, csa_tree_add_51_79_groupi_n_3418, csa_tree_add_51_79_groupi_n_3419, csa_tree_add_51_79_groupi_n_3420, csa_tree_add_51_79_groupi_n_3421, csa_tree_add_51_79_groupi_n_3422, csa_tree_add_51_79_groupi_n_3423;
  wire csa_tree_add_51_79_groupi_n_3424, csa_tree_add_51_79_groupi_n_3425, csa_tree_add_51_79_groupi_n_3426, csa_tree_add_51_79_groupi_n_3427, csa_tree_add_51_79_groupi_n_3428, csa_tree_add_51_79_groupi_n_3429, csa_tree_add_51_79_groupi_n_3430, csa_tree_add_51_79_groupi_n_3431;
  wire csa_tree_add_51_79_groupi_n_3432, csa_tree_add_51_79_groupi_n_3433, csa_tree_add_51_79_groupi_n_3434, csa_tree_add_51_79_groupi_n_3435, csa_tree_add_51_79_groupi_n_3436, csa_tree_add_51_79_groupi_n_3437, csa_tree_add_51_79_groupi_n_3438, csa_tree_add_51_79_groupi_n_3439;
  wire csa_tree_add_51_79_groupi_n_3440, csa_tree_add_51_79_groupi_n_3441, csa_tree_add_51_79_groupi_n_3442, csa_tree_add_51_79_groupi_n_3443, csa_tree_add_51_79_groupi_n_3444, csa_tree_add_51_79_groupi_n_3445, csa_tree_add_51_79_groupi_n_3446, csa_tree_add_51_79_groupi_n_3447;
  wire csa_tree_add_51_79_groupi_n_3448, csa_tree_add_51_79_groupi_n_3449, csa_tree_add_51_79_groupi_n_3450, csa_tree_add_51_79_groupi_n_3451, csa_tree_add_51_79_groupi_n_3452, csa_tree_add_51_79_groupi_n_3453, csa_tree_add_51_79_groupi_n_3454, csa_tree_add_51_79_groupi_n_3455;
  wire csa_tree_add_51_79_groupi_n_3456, csa_tree_add_51_79_groupi_n_3457, csa_tree_add_51_79_groupi_n_3458, csa_tree_add_51_79_groupi_n_3459, csa_tree_add_51_79_groupi_n_3460, csa_tree_add_51_79_groupi_n_3461, csa_tree_add_51_79_groupi_n_3462, csa_tree_add_51_79_groupi_n_3463;
  wire csa_tree_add_51_79_groupi_n_3464, csa_tree_add_51_79_groupi_n_3465, csa_tree_add_51_79_groupi_n_3466, csa_tree_add_51_79_groupi_n_3467, csa_tree_add_51_79_groupi_n_3468, csa_tree_add_51_79_groupi_n_3469, csa_tree_add_51_79_groupi_n_3470, csa_tree_add_51_79_groupi_n_3471;
  wire csa_tree_add_51_79_groupi_n_3472, csa_tree_add_51_79_groupi_n_3473, csa_tree_add_51_79_groupi_n_3474, csa_tree_add_51_79_groupi_n_3475, csa_tree_add_51_79_groupi_n_3476, csa_tree_add_51_79_groupi_n_3477, csa_tree_add_51_79_groupi_n_3478, csa_tree_add_51_79_groupi_n_3479;
  wire csa_tree_add_51_79_groupi_n_3480, csa_tree_add_51_79_groupi_n_3481, csa_tree_add_51_79_groupi_n_3482, csa_tree_add_51_79_groupi_n_3483, csa_tree_add_51_79_groupi_n_3484, csa_tree_add_51_79_groupi_n_3485, csa_tree_add_51_79_groupi_n_3486, csa_tree_add_51_79_groupi_n_3487;
  wire csa_tree_add_51_79_groupi_n_3488, csa_tree_add_51_79_groupi_n_3489, csa_tree_add_51_79_groupi_n_3490, csa_tree_add_51_79_groupi_n_3491, csa_tree_add_51_79_groupi_n_3492, csa_tree_add_51_79_groupi_n_3493, csa_tree_add_51_79_groupi_n_3494, csa_tree_add_51_79_groupi_n_3495;
  wire csa_tree_add_51_79_groupi_n_3496, csa_tree_add_51_79_groupi_n_3497, csa_tree_add_51_79_groupi_n_3498, csa_tree_add_51_79_groupi_n_3499, csa_tree_add_51_79_groupi_n_3500, csa_tree_add_51_79_groupi_n_3501, csa_tree_add_51_79_groupi_n_3502, csa_tree_add_51_79_groupi_n_3503;
  wire csa_tree_add_51_79_groupi_n_3504, csa_tree_add_51_79_groupi_n_3505, csa_tree_add_51_79_groupi_n_3506, csa_tree_add_51_79_groupi_n_3507, csa_tree_add_51_79_groupi_n_3508, csa_tree_add_51_79_groupi_n_3509, csa_tree_add_51_79_groupi_n_3510, csa_tree_add_51_79_groupi_n_3511;
  wire csa_tree_add_51_79_groupi_n_3512, csa_tree_add_51_79_groupi_n_3513, csa_tree_add_51_79_groupi_n_3514, csa_tree_add_51_79_groupi_n_3515, csa_tree_add_51_79_groupi_n_3516, csa_tree_add_51_79_groupi_n_3517, csa_tree_add_51_79_groupi_n_3518, csa_tree_add_51_79_groupi_n_3519;
  wire csa_tree_add_51_79_groupi_n_3520, csa_tree_add_51_79_groupi_n_3521, csa_tree_add_51_79_groupi_n_3522, csa_tree_add_51_79_groupi_n_3523, csa_tree_add_51_79_groupi_n_3524, csa_tree_add_51_79_groupi_n_3525, csa_tree_add_51_79_groupi_n_3526, csa_tree_add_51_79_groupi_n_3527;
  wire csa_tree_add_51_79_groupi_n_3528, csa_tree_add_51_79_groupi_n_3529, csa_tree_add_51_79_groupi_n_3530, csa_tree_add_51_79_groupi_n_3531, csa_tree_add_51_79_groupi_n_3532, csa_tree_add_51_79_groupi_n_3533, csa_tree_add_51_79_groupi_n_3534, csa_tree_add_51_79_groupi_n_3535;
  wire csa_tree_add_51_79_groupi_n_3536, csa_tree_add_51_79_groupi_n_3537, csa_tree_add_51_79_groupi_n_3538, csa_tree_add_51_79_groupi_n_3539, csa_tree_add_51_79_groupi_n_3540, csa_tree_add_51_79_groupi_n_3541, csa_tree_add_51_79_groupi_n_3542, csa_tree_add_51_79_groupi_n_3543;
  wire csa_tree_add_51_79_groupi_n_3544, csa_tree_add_51_79_groupi_n_3545, csa_tree_add_51_79_groupi_n_3546, csa_tree_add_51_79_groupi_n_3547, csa_tree_add_51_79_groupi_n_3548, csa_tree_add_51_79_groupi_n_3549, csa_tree_add_51_79_groupi_n_3550, csa_tree_add_51_79_groupi_n_3551;
  wire csa_tree_add_51_79_groupi_n_3552, csa_tree_add_51_79_groupi_n_3553, csa_tree_add_51_79_groupi_n_3554, csa_tree_add_51_79_groupi_n_3555, csa_tree_add_51_79_groupi_n_3556, csa_tree_add_51_79_groupi_n_3557, csa_tree_add_51_79_groupi_n_3558, csa_tree_add_51_79_groupi_n_3559;
  wire csa_tree_add_51_79_groupi_n_3560, csa_tree_add_51_79_groupi_n_3561, csa_tree_add_51_79_groupi_n_3562, csa_tree_add_51_79_groupi_n_3563, csa_tree_add_51_79_groupi_n_3564, csa_tree_add_51_79_groupi_n_3565, csa_tree_add_51_79_groupi_n_3566, csa_tree_add_51_79_groupi_n_3567;
  wire csa_tree_add_51_79_groupi_n_3568, csa_tree_add_51_79_groupi_n_3569, csa_tree_add_51_79_groupi_n_3570, csa_tree_add_51_79_groupi_n_3571, csa_tree_add_51_79_groupi_n_3572, csa_tree_add_51_79_groupi_n_3573, csa_tree_add_51_79_groupi_n_3574, csa_tree_add_51_79_groupi_n_3575;
  wire csa_tree_add_51_79_groupi_n_3576, csa_tree_add_51_79_groupi_n_3577, csa_tree_add_51_79_groupi_n_3578, csa_tree_add_51_79_groupi_n_3579, csa_tree_add_51_79_groupi_n_3580, csa_tree_add_51_79_groupi_n_3581, csa_tree_add_51_79_groupi_n_3582, csa_tree_add_51_79_groupi_n_3583;
  wire csa_tree_add_51_79_groupi_n_3584, csa_tree_add_51_79_groupi_n_3585, csa_tree_add_51_79_groupi_n_3586, csa_tree_add_51_79_groupi_n_3587, csa_tree_add_51_79_groupi_n_3588, csa_tree_add_51_79_groupi_n_3589, csa_tree_add_51_79_groupi_n_3590, csa_tree_add_51_79_groupi_n_3591;
  wire csa_tree_add_51_79_groupi_n_3592, csa_tree_add_51_79_groupi_n_3593, csa_tree_add_51_79_groupi_n_3594, csa_tree_add_51_79_groupi_n_3595, csa_tree_add_51_79_groupi_n_3596, csa_tree_add_51_79_groupi_n_3597, csa_tree_add_51_79_groupi_n_3598, csa_tree_add_51_79_groupi_n_3599;
  wire csa_tree_add_51_79_groupi_n_3600, csa_tree_add_51_79_groupi_n_3601, csa_tree_add_51_79_groupi_n_3602, csa_tree_add_51_79_groupi_n_3603, csa_tree_add_51_79_groupi_n_3604, csa_tree_add_51_79_groupi_n_3605, csa_tree_add_51_79_groupi_n_3606, csa_tree_add_51_79_groupi_n_3607;
  wire csa_tree_add_51_79_groupi_n_3608, csa_tree_add_51_79_groupi_n_3609, csa_tree_add_51_79_groupi_n_3610, csa_tree_add_51_79_groupi_n_3611, csa_tree_add_51_79_groupi_n_3612, csa_tree_add_51_79_groupi_n_3613, csa_tree_add_51_79_groupi_n_3614, csa_tree_add_51_79_groupi_n_3615;
  wire csa_tree_add_51_79_groupi_n_3616, csa_tree_add_51_79_groupi_n_3617, csa_tree_add_51_79_groupi_n_3618, csa_tree_add_51_79_groupi_n_3619, csa_tree_add_51_79_groupi_n_3620, csa_tree_add_51_79_groupi_n_3621, csa_tree_add_51_79_groupi_n_3622, csa_tree_add_51_79_groupi_n_3623;
  wire csa_tree_add_51_79_groupi_n_3624, csa_tree_add_51_79_groupi_n_3625, csa_tree_add_51_79_groupi_n_3626, csa_tree_add_51_79_groupi_n_3627, csa_tree_add_51_79_groupi_n_3628, csa_tree_add_51_79_groupi_n_3629, csa_tree_add_51_79_groupi_n_3630, csa_tree_add_51_79_groupi_n_3631;
  wire csa_tree_add_51_79_groupi_n_3632, csa_tree_add_51_79_groupi_n_3633, csa_tree_add_51_79_groupi_n_3634, csa_tree_add_51_79_groupi_n_3635, csa_tree_add_51_79_groupi_n_3636, csa_tree_add_51_79_groupi_n_3637, csa_tree_add_51_79_groupi_n_3638, csa_tree_add_51_79_groupi_n_3639;
  wire csa_tree_add_51_79_groupi_n_3640, csa_tree_add_51_79_groupi_n_3641, csa_tree_add_51_79_groupi_n_3642, csa_tree_add_51_79_groupi_n_3643, csa_tree_add_51_79_groupi_n_3644, csa_tree_add_51_79_groupi_n_3645, csa_tree_add_51_79_groupi_n_3646, csa_tree_add_51_79_groupi_n_3647;
  wire csa_tree_add_51_79_groupi_n_3648, csa_tree_add_51_79_groupi_n_3649, csa_tree_add_51_79_groupi_n_3650, csa_tree_add_51_79_groupi_n_3651, csa_tree_add_51_79_groupi_n_3652, csa_tree_add_51_79_groupi_n_3653, csa_tree_add_51_79_groupi_n_3654, csa_tree_add_51_79_groupi_n_3655;
  wire csa_tree_add_51_79_groupi_n_3656, csa_tree_add_51_79_groupi_n_3657, csa_tree_add_51_79_groupi_n_3658, csa_tree_add_51_79_groupi_n_3659, csa_tree_add_51_79_groupi_n_3660, csa_tree_add_51_79_groupi_n_3661, csa_tree_add_51_79_groupi_n_3662, csa_tree_add_51_79_groupi_n_3663;
  wire csa_tree_add_51_79_groupi_n_3664, csa_tree_add_51_79_groupi_n_3665, csa_tree_add_51_79_groupi_n_3666, csa_tree_add_51_79_groupi_n_3667, csa_tree_add_51_79_groupi_n_3668, csa_tree_add_51_79_groupi_n_3669, csa_tree_add_51_79_groupi_n_3670, csa_tree_add_51_79_groupi_n_3671;
  wire csa_tree_add_51_79_groupi_n_3672, csa_tree_add_51_79_groupi_n_3673, csa_tree_add_51_79_groupi_n_3674, csa_tree_add_51_79_groupi_n_3675, csa_tree_add_51_79_groupi_n_3676, csa_tree_add_51_79_groupi_n_3677, csa_tree_add_51_79_groupi_n_3678, csa_tree_add_51_79_groupi_n_3679;
  wire csa_tree_add_51_79_groupi_n_3680, csa_tree_add_51_79_groupi_n_3681, csa_tree_add_51_79_groupi_n_3682, csa_tree_add_51_79_groupi_n_3683, csa_tree_add_51_79_groupi_n_3684, csa_tree_add_51_79_groupi_n_3685, csa_tree_add_51_79_groupi_n_3686, csa_tree_add_51_79_groupi_n_3687;
  wire csa_tree_add_51_79_groupi_n_3688, csa_tree_add_51_79_groupi_n_3689, csa_tree_add_51_79_groupi_n_3690, csa_tree_add_51_79_groupi_n_3691, csa_tree_add_51_79_groupi_n_3692, csa_tree_add_51_79_groupi_n_3693, csa_tree_add_51_79_groupi_n_3694, csa_tree_add_51_79_groupi_n_3695;
  wire csa_tree_add_51_79_groupi_n_3696, csa_tree_add_51_79_groupi_n_3697, csa_tree_add_51_79_groupi_n_3698, csa_tree_add_51_79_groupi_n_3699, csa_tree_add_51_79_groupi_n_3700, csa_tree_add_51_79_groupi_n_3701, csa_tree_add_51_79_groupi_n_3702, csa_tree_add_51_79_groupi_n_3703;
  wire csa_tree_add_51_79_groupi_n_3704, csa_tree_add_51_79_groupi_n_3705, csa_tree_add_51_79_groupi_n_3706, csa_tree_add_51_79_groupi_n_3707, csa_tree_add_51_79_groupi_n_3708, csa_tree_add_51_79_groupi_n_3709, csa_tree_add_51_79_groupi_n_3710, csa_tree_add_51_79_groupi_n_3711;
  wire csa_tree_add_51_79_groupi_n_3712, csa_tree_add_51_79_groupi_n_3713, csa_tree_add_51_79_groupi_n_3714, csa_tree_add_51_79_groupi_n_3715, csa_tree_add_51_79_groupi_n_3716, csa_tree_add_51_79_groupi_n_3717, csa_tree_add_51_79_groupi_n_3718, csa_tree_add_51_79_groupi_n_3719;
  wire csa_tree_add_51_79_groupi_n_3720, csa_tree_add_51_79_groupi_n_3721, csa_tree_add_51_79_groupi_n_3722, csa_tree_add_51_79_groupi_n_3723, csa_tree_add_51_79_groupi_n_3724, csa_tree_add_51_79_groupi_n_3725, csa_tree_add_51_79_groupi_n_3726, csa_tree_add_51_79_groupi_n_3727;
  wire csa_tree_add_51_79_groupi_n_3728, csa_tree_add_51_79_groupi_n_3729, csa_tree_add_51_79_groupi_n_3730, csa_tree_add_51_79_groupi_n_3731, csa_tree_add_51_79_groupi_n_3732, csa_tree_add_51_79_groupi_n_3733, csa_tree_add_51_79_groupi_n_3734, csa_tree_add_51_79_groupi_n_3735;
  wire csa_tree_add_51_79_groupi_n_3736, csa_tree_add_51_79_groupi_n_3737, csa_tree_add_51_79_groupi_n_3738, csa_tree_add_51_79_groupi_n_3739, csa_tree_add_51_79_groupi_n_3740, csa_tree_add_51_79_groupi_n_3741, csa_tree_add_51_79_groupi_n_3742, csa_tree_add_51_79_groupi_n_3743;
  wire csa_tree_add_51_79_groupi_n_3744, csa_tree_add_51_79_groupi_n_3745, csa_tree_add_51_79_groupi_n_3746, csa_tree_add_51_79_groupi_n_3747, csa_tree_add_51_79_groupi_n_3748, csa_tree_add_51_79_groupi_n_3749, csa_tree_add_51_79_groupi_n_3750, csa_tree_add_51_79_groupi_n_3751;
  wire csa_tree_add_51_79_groupi_n_3752, csa_tree_add_51_79_groupi_n_3753, csa_tree_add_51_79_groupi_n_3754, csa_tree_add_51_79_groupi_n_3755, csa_tree_add_51_79_groupi_n_3756, csa_tree_add_51_79_groupi_n_3757, csa_tree_add_51_79_groupi_n_3758, csa_tree_add_51_79_groupi_n_3759;
  wire csa_tree_add_51_79_groupi_n_3760, csa_tree_add_51_79_groupi_n_3761, csa_tree_add_51_79_groupi_n_3762, csa_tree_add_51_79_groupi_n_3763, csa_tree_add_51_79_groupi_n_3764, csa_tree_add_51_79_groupi_n_3765, csa_tree_add_51_79_groupi_n_3766, csa_tree_add_51_79_groupi_n_3767;
  wire csa_tree_add_51_79_groupi_n_3768, csa_tree_add_51_79_groupi_n_3769, csa_tree_add_51_79_groupi_n_3770, csa_tree_add_51_79_groupi_n_3771, csa_tree_add_51_79_groupi_n_3772, csa_tree_add_51_79_groupi_n_3773, csa_tree_add_51_79_groupi_n_3774, csa_tree_add_51_79_groupi_n_3775;
  wire csa_tree_add_51_79_groupi_n_3776, csa_tree_add_51_79_groupi_n_3777, csa_tree_add_51_79_groupi_n_3778, csa_tree_add_51_79_groupi_n_3779, csa_tree_add_51_79_groupi_n_3780, csa_tree_add_51_79_groupi_n_3781, csa_tree_add_51_79_groupi_n_3782, csa_tree_add_51_79_groupi_n_3783;
  wire csa_tree_add_51_79_groupi_n_3784, csa_tree_add_51_79_groupi_n_3785, csa_tree_add_51_79_groupi_n_3786, csa_tree_add_51_79_groupi_n_3787, csa_tree_add_51_79_groupi_n_3788, csa_tree_add_51_79_groupi_n_3789, csa_tree_add_51_79_groupi_n_3790, csa_tree_add_51_79_groupi_n_3791;
  wire csa_tree_add_51_79_groupi_n_3792, csa_tree_add_51_79_groupi_n_3793, csa_tree_add_51_79_groupi_n_3794, csa_tree_add_51_79_groupi_n_3795, csa_tree_add_51_79_groupi_n_3796, csa_tree_add_51_79_groupi_n_3797, csa_tree_add_51_79_groupi_n_3798, csa_tree_add_51_79_groupi_n_3799;
  wire csa_tree_add_51_79_groupi_n_3800, csa_tree_add_51_79_groupi_n_3801, csa_tree_add_51_79_groupi_n_3802, csa_tree_add_51_79_groupi_n_3803, csa_tree_add_51_79_groupi_n_3804, csa_tree_add_51_79_groupi_n_3805, csa_tree_add_51_79_groupi_n_3806, csa_tree_add_51_79_groupi_n_3807;
  wire csa_tree_add_51_79_groupi_n_3808, csa_tree_add_51_79_groupi_n_3809, csa_tree_add_51_79_groupi_n_3810, csa_tree_add_51_79_groupi_n_3811, csa_tree_add_51_79_groupi_n_3812, csa_tree_add_51_79_groupi_n_3813, csa_tree_add_51_79_groupi_n_3814, csa_tree_add_51_79_groupi_n_3815;
  wire csa_tree_add_51_79_groupi_n_3816, csa_tree_add_51_79_groupi_n_3817, csa_tree_add_51_79_groupi_n_3818, csa_tree_add_51_79_groupi_n_3819, csa_tree_add_51_79_groupi_n_3820, csa_tree_add_51_79_groupi_n_3821, csa_tree_add_51_79_groupi_n_3822, csa_tree_add_51_79_groupi_n_3823;
  wire csa_tree_add_51_79_groupi_n_3824, csa_tree_add_51_79_groupi_n_3825, csa_tree_add_51_79_groupi_n_3826, csa_tree_add_51_79_groupi_n_3827, csa_tree_add_51_79_groupi_n_3828, csa_tree_add_51_79_groupi_n_3829, csa_tree_add_51_79_groupi_n_3830, csa_tree_add_51_79_groupi_n_3831;
  wire csa_tree_add_51_79_groupi_n_3832, csa_tree_add_51_79_groupi_n_3833, csa_tree_add_51_79_groupi_n_3834, csa_tree_add_51_79_groupi_n_3835, csa_tree_add_51_79_groupi_n_3836, csa_tree_add_51_79_groupi_n_3837, csa_tree_add_51_79_groupi_n_3838, csa_tree_add_51_79_groupi_n_3839;
  wire csa_tree_add_51_79_groupi_n_3840, csa_tree_add_51_79_groupi_n_3841, csa_tree_add_51_79_groupi_n_3842, csa_tree_add_51_79_groupi_n_3843, csa_tree_add_51_79_groupi_n_3844, csa_tree_add_51_79_groupi_n_3845, csa_tree_add_51_79_groupi_n_3846, csa_tree_add_51_79_groupi_n_3847;
  wire csa_tree_add_51_79_groupi_n_3848, csa_tree_add_51_79_groupi_n_3849, csa_tree_add_51_79_groupi_n_3850, csa_tree_add_51_79_groupi_n_3851, csa_tree_add_51_79_groupi_n_3852, csa_tree_add_51_79_groupi_n_3853, csa_tree_add_51_79_groupi_n_3854, csa_tree_add_51_79_groupi_n_3855;
  wire csa_tree_add_51_79_groupi_n_3856, csa_tree_add_51_79_groupi_n_3857, csa_tree_add_51_79_groupi_n_3858, csa_tree_add_51_79_groupi_n_3859, csa_tree_add_51_79_groupi_n_3860, csa_tree_add_51_79_groupi_n_3861, csa_tree_add_51_79_groupi_n_3862, csa_tree_add_51_79_groupi_n_3863;
  wire csa_tree_add_51_79_groupi_n_3864, csa_tree_add_51_79_groupi_n_3865, csa_tree_add_51_79_groupi_n_3866, csa_tree_add_51_79_groupi_n_3867, csa_tree_add_51_79_groupi_n_3868, csa_tree_add_51_79_groupi_n_3869, csa_tree_add_51_79_groupi_n_3870, csa_tree_add_51_79_groupi_n_3871;
  wire csa_tree_add_51_79_groupi_n_3872, csa_tree_add_51_79_groupi_n_3873, csa_tree_add_51_79_groupi_n_3874, csa_tree_add_51_79_groupi_n_3875, csa_tree_add_51_79_groupi_n_3876, csa_tree_add_51_79_groupi_n_3877, csa_tree_add_51_79_groupi_n_3878, csa_tree_add_51_79_groupi_n_3879;
  wire csa_tree_add_51_79_groupi_n_3880, csa_tree_add_51_79_groupi_n_3881, csa_tree_add_51_79_groupi_n_3882, csa_tree_add_51_79_groupi_n_3883, csa_tree_add_51_79_groupi_n_3884, csa_tree_add_51_79_groupi_n_3885, csa_tree_add_51_79_groupi_n_3886, csa_tree_add_51_79_groupi_n_3887;
  wire csa_tree_add_51_79_groupi_n_3888, csa_tree_add_51_79_groupi_n_3889, csa_tree_add_51_79_groupi_n_3890, csa_tree_add_51_79_groupi_n_3891, csa_tree_add_51_79_groupi_n_3892, csa_tree_add_51_79_groupi_n_3893, csa_tree_add_51_79_groupi_n_3894, csa_tree_add_51_79_groupi_n_3895;
  wire csa_tree_add_51_79_groupi_n_3896, csa_tree_add_51_79_groupi_n_3897, csa_tree_add_51_79_groupi_n_3898, csa_tree_add_51_79_groupi_n_3899, csa_tree_add_51_79_groupi_n_3900, csa_tree_add_51_79_groupi_n_3901, csa_tree_add_51_79_groupi_n_3902, csa_tree_add_51_79_groupi_n_3903;
  wire csa_tree_add_51_79_groupi_n_3904, csa_tree_add_51_79_groupi_n_3905, csa_tree_add_51_79_groupi_n_3906, csa_tree_add_51_79_groupi_n_3907, csa_tree_add_51_79_groupi_n_3908, csa_tree_add_51_79_groupi_n_3909, csa_tree_add_51_79_groupi_n_3910, csa_tree_add_51_79_groupi_n_3911;
  wire csa_tree_add_51_79_groupi_n_3912, csa_tree_add_51_79_groupi_n_3913, csa_tree_add_51_79_groupi_n_3914, csa_tree_add_51_79_groupi_n_3915, csa_tree_add_51_79_groupi_n_3916, csa_tree_add_51_79_groupi_n_3917, csa_tree_add_51_79_groupi_n_3918, csa_tree_add_51_79_groupi_n_3919;
  wire csa_tree_add_51_79_groupi_n_3920, csa_tree_add_51_79_groupi_n_3921, csa_tree_add_51_79_groupi_n_3922, csa_tree_add_51_79_groupi_n_3923, csa_tree_add_51_79_groupi_n_3924, csa_tree_add_51_79_groupi_n_3925, csa_tree_add_51_79_groupi_n_3926, csa_tree_add_51_79_groupi_n_3927;
  wire csa_tree_add_51_79_groupi_n_3928, csa_tree_add_51_79_groupi_n_3929, csa_tree_add_51_79_groupi_n_3930, csa_tree_add_51_79_groupi_n_3931, csa_tree_add_51_79_groupi_n_3932, csa_tree_add_51_79_groupi_n_3933, csa_tree_add_51_79_groupi_n_3934, csa_tree_add_51_79_groupi_n_3935;
  wire csa_tree_add_51_79_groupi_n_3936, csa_tree_add_51_79_groupi_n_3937, csa_tree_add_51_79_groupi_n_3938, csa_tree_add_51_79_groupi_n_3939, csa_tree_add_51_79_groupi_n_3940, csa_tree_add_51_79_groupi_n_3941, csa_tree_add_51_79_groupi_n_3942, csa_tree_add_51_79_groupi_n_3943;
  wire csa_tree_add_51_79_groupi_n_3944, csa_tree_add_51_79_groupi_n_3945, csa_tree_add_51_79_groupi_n_3946, csa_tree_add_51_79_groupi_n_3947, csa_tree_add_51_79_groupi_n_3948, csa_tree_add_51_79_groupi_n_3949, csa_tree_add_51_79_groupi_n_3950, csa_tree_add_51_79_groupi_n_3951;
  wire csa_tree_add_51_79_groupi_n_3952, csa_tree_add_51_79_groupi_n_3953, csa_tree_add_51_79_groupi_n_3954, csa_tree_add_51_79_groupi_n_3955, csa_tree_add_51_79_groupi_n_3956, csa_tree_add_51_79_groupi_n_3957, csa_tree_add_51_79_groupi_n_3958, csa_tree_add_51_79_groupi_n_3959;
  wire csa_tree_add_51_79_groupi_n_3960, csa_tree_add_51_79_groupi_n_3961, csa_tree_add_51_79_groupi_n_3962, csa_tree_add_51_79_groupi_n_3963, csa_tree_add_51_79_groupi_n_3964, csa_tree_add_51_79_groupi_n_3965, csa_tree_add_51_79_groupi_n_3966, csa_tree_add_51_79_groupi_n_3967;
  wire csa_tree_add_51_79_groupi_n_3968, csa_tree_add_51_79_groupi_n_3969, csa_tree_add_51_79_groupi_n_3970, csa_tree_add_51_79_groupi_n_3971, csa_tree_add_51_79_groupi_n_3972, csa_tree_add_51_79_groupi_n_3973, csa_tree_add_51_79_groupi_n_3974, csa_tree_add_51_79_groupi_n_3975;
  wire csa_tree_add_51_79_groupi_n_3976, csa_tree_add_51_79_groupi_n_3977, csa_tree_add_51_79_groupi_n_3978, csa_tree_add_51_79_groupi_n_3979, csa_tree_add_51_79_groupi_n_3980, csa_tree_add_51_79_groupi_n_3981, csa_tree_add_51_79_groupi_n_3982, csa_tree_add_51_79_groupi_n_3983;
  wire csa_tree_add_51_79_groupi_n_3984, csa_tree_add_51_79_groupi_n_3985, csa_tree_add_51_79_groupi_n_3986, csa_tree_add_51_79_groupi_n_3987, csa_tree_add_51_79_groupi_n_3988, csa_tree_add_51_79_groupi_n_3989, csa_tree_add_51_79_groupi_n_3990, csa_tree_add_51_79_groupi_n_3991;
  wire csa_tree_add_51_79_groupi_n_3992, csa_tree_add_51_79_groupi_n_3993, csa_tree_add_51_79_groupi_n_3994, csa_tree_add_51_79_groupi_n_3995, csa_tree_add_51_79_groupi_n_3996, csa_tree_add_51_79_groupi_n_3997, csa_tree_add_51_79_groupi_n_3998, csa_tree_add_51_79_groupi_n_3999;
  wire csa_tree_add_51_79_groupi_n_4000, csa_tree_add_51_79_groupi_n_4001, csa_tree_add_51_79_groupi_n_4002, csa_tree_add_51_79_groupi_n_4003, csa_tree_add_51_79_groupi_n_4004, csa_tree_add_51_79_groupi_n_4005, csa_tree_add_51_79_groupi_n_4006, csa_tree_add_51_79_groupi_n_4007;
  wire csa_tree_add_51_79_groupi_n_4008, csa_tree_add_51_79_groupi_n_4009, csa_tree_add_51_79_groupi_n_4010, csa_tree_add_51_79_groupi_n_4011, csa_tree_add_51_79_groupi_n_4012, csa_tree_add_51_79_groupi_n_4013, csa_tree_add_51_79_groupi_n_4014, csa_tree_add_51_79_groupi_n_4015;
  wire csa_tree_add_51_79_groupi_n_4016, csa_tree_add_51_79_groupi_n_4017, csa_tree_add_51_79_groupi_n_4018, csa_tree_add_51_79_groupi_n_4019, csa_tree_add_51_79_groupi_n_4020, csa_tree_add_51_79_groupi_n_4021, csa_tree_add_51_79_groupi_n_4022, csa_tree_add_51_79_groupi_n_4023;
  wire csa_tree_add_51_79_groupi_n_4024, csa_tree_add_51_79_groupi_n_4025, csa_tree_add_51_79_groupi_n_4026, csa_tree_add_51_79_groupi_n_4027, csa_tree_add_51_79_groupi_n_4028, csa_tree_add_51_79_groupi_n_4029, csa_tree_add_51_79_groupi_n_4030, csa_tree_add_51_79_groupi_n_4031;
  wire csa_tree_add_51_79_groupi_n_4032, csa_tree_add_51_79_groupi_n_4033, csa_tree_add_51_79_groupi_n_4034, csa_tree_add_51_79_groupi_n_4035, csa_tree_add_51_79_groupi_n_4036, csa_tree_add_51_79_groupi_n_4037, csa_tree_add_51_79_groupi_n_4038, csa_tree_add_51_79_groupi_n_4039;
  wire csa_tree_add_51_79_groupi_n_4040, csa_tree_add_51_79_groupi_n_4041, csa_tree_add_51_79_groupi_n_4042, csa_tree_add_51_79_groupi_n_4043, csa_tree_add_51_79_groupi_n_4044, csa_tree_add_51_79_groupi_n_4045, csa_tree_add_51_79_groupi_n_4046, csa_tree_add_51_79_groupi_n_4047;
  wire csa_tree_add_51_79_groupi_n_4048, csa_tree_add_51_79_groupi_n_4049, csa_tree_add_51_79_groupi_n_4050, csa_tree_add_51_79_groupi_n_4051, csa_tree_add_51_79_groupi_n_4052, csa_tree_add_51_79_groupi_n_4053, csa_tree_add_51_79_groupi_n_4054, csa_tree_add_51_79_groupi_n_4055;
  wire csa_tree_add_51_79_groupi_n_4056, csa_tree_add_51_79_groupi_n_4057, csa_tree_add_51_79_groupi_n_4058, csa_tree_add_51_79_groupi_n_4059, csa_tree_add_51_79_groupi_n_4060, csa_tree_add_51_79_groupi_n_4061, csa_tree_add_51_79_groupi_n_4062, csa_tree_add_51_79_groupi_n_4063;
  wire csa_tree_add_51_79_groupi_n_4064, csa_tree_add_51_79_groupi_n_4065, csa_tree_add_51_79_groupi_n_4066, csa_tree_add_51_79_groupi_n_4067, csa_tree_add_51_79_groupi_n_4068, csa_tree_add_51_79_groupi_n_4069, csa_tree_add_51_79_groupi_n_4070, csa_tree_add_51_79_groupi_n_4071;
  wire csa_tree_add_51_79_groupi_n_4072, csa_tree_add_51_79_groupi_n_4073, csa_tree_add_51_79_groupi_n_4074, csa_tree_add_51_79_groupi_n_4075, csa_tree_add_51_79_groupi_n_4076, csa_tree_add_51_79_groupi_n_4077, csa_tree_add_51_79_groupi_n_4078, csa_tree_add_51_79_groupi_n_4079;
  wire csa_tree_add_51_79_groupi_n_4080, csa_tree_add_51_79_groupi_n_4081, csa_tree_add_51_79_groupi_n_4082, csa_tree_add_51_79_groupi_n_4083, csa_tree_add_51_79_groupi_n_4084, csa_tree_add_51_79_groupi_n_4085, csa_tree_add_51_79_groupi_n_4086, csa_tree_add_51_79_groupi_n_4087;
  wire csa_tree_add_51_79_groupi_n_4088, csa_tree_add_51_79_groupi_n_4089, csa_tree_add_51_79_groupi_n_4090, csa_tree_add_51_79_groupi_n_4091, csa_tree_add_51_79_groupi_n_4092, csa_tree_add_51_79_groupi_n_4093, csa_tree_add_51_79_groupi_n_4094, csa_tree_add_51_79_groupi_n_4095;
  wire csa_tree_add_51_79_groupi_n_4096, csa_tree_add_51_79_groupi_n_4097, csa_tree_add_51_79_groupi_n_4098, csa_tree_add_51_79_groupi_n_4099, csa_tree_add_51_79_groupi_n_4100, csa_tree_add_51_79_groupi_n_4101, csa_tree_add_51_79_groupi_n_4102, csa_tree_add_51_79_groupi_n_4103;
  wire csa_tree_add_51_79_groupi_n_4104, csa_tree_add_51_79_groupi_n_4105, csa_tree_add_51_79_groupi_n_4106, csa_tree_add_51_79_groupi_n_4107, csa_tree_add_51_79_groupi_n_4108, csa_tree_add_51_79_groupi_n_4109, csa_tree_add_51_79_groupi_n_4110, csa_tree_add_51_79_groupi_n_4111;
  wire csa_tree_add_51_79_groupi_n_4112, csa_tree_add_51_79_groupi_n_4113, csa_tree_add_51_79_groupi_n_4114, csa_tree_add_51_79_groupi_n_4115, csa_tree_add_51_79_groupi_n_4116, csa_tree_add_51_79_groupi_n_4117, csa_tree_add_51_79_groupi_n_4118, csa_tree_add_51_79_groupi_n_4119;
  wire csa_tree_add_51_79_groupi_n_4120, csa_tree_add_51_79_groupi_n_4121, csa_tree_add_51_79_groupi_n_4122, csa_tree_add_51_79_groupi_n_4123, csa_tree_add_51_79_groupi_n_4124, csa_tree_add_51_79_groupi_n_4125, csa_tree_add_51_79_groupi_n_4126, csa_tree_add_51_79_groupi_n_4127;
  wire csa_tree_add_51_79_groupi_n_4128, csa_tree_add_51_79_groupi_n_4129, csa_tree_add_51_79_groupi_n_4130, csa_tree_add_51_79_groupi_n_4131, csa_tree_add_51_79_groupi_n_4132, csa_tree_add_51_79_groupi_n_4133, csa_tree_add_51_79_groupi_n_4134, csa_tree_add_51_79_groupi_n_4135;
  wire csa_tree_add_51_79_groupi_n_4136, csa_tree_add_51_79_groupi_n_4137, csa_tree_add_51_79_groupi_n_4138, csa_tree_add_51_79_groupi_n_4139, csa_tree_add_51_79_groupi_n_4140, csa_tree_add_51_79_groupi_n_4141, csa_tree_add_51_79_groupi_n_4142, csa_tree_add_51_79_groupi_n_4143;
  wire csa_tree_add_51_79_groupi_n_4144, csa_tree_add_51_79_groupi_n_4145, csa_tree_add_51_79_groupi_n_4146, csa_tree_add_51_79_groupi_n_4147, csa_tree_add_51_79_groupi_n_4148, csa_tree_add_51_79_groupi_n_4149, csa_tree_add_51_79_groupi_n_4150, csa_tree_add_51_79_groupi_n_4151;
  wire csa_tree_add_51_79_groupi_n_4152, csa_tree_add_51_79_groupi_n_4153, csa_tree_add_51_79_groupi_n_4154, csa_tree_add_51_79_groupi_n_4155, csa_tree_add_51_79_groupi_n_4156, csa_tree_add_51_79_groupi_n_4157, csa_tree_add_51_79_groupi_n_4158, csa_tree_add_51_79_groupi_n_4159;
  wire csa_tree_add_51_79_groupi_n_4160, csa_tree_add_51_79_groupi_n_4161, csa_tree_add_51_79_groupi_n_4162, csa_tree_add_51_79_groupi_n_4163, csa_tree_add_51_79_groupi_n_4164, csa_tree_add_51_79_groupi_n_4165, csa_tree_add_51_79_groupi_n_4166, csa_tree_add_51_79_groupi_n_4167;
  wire csa_tree_add_51_79_groupi_n_4168, csa_tree_add_51_79_groupi_n_4169, csa_tree_add_51_79_groupi_n_4170, csa_tree_add_51_79_groupi_n_4171, csa_tree_add_51_79_groupi_n_4172, csa_tree_add_51_79_groupi_n_4173, csa_tree_add_51_79_groupi_n_4174, csa_tree_add_51_79_groupi_n_4175;
  wire csa_tree_add_51_79_groupi_n_4176, csa_tree_add_51_79_groupi_n_4177, csa_tree_add_51_79_groupi_n_4178, csa_tree_add_51_79_groupi_n_4179, csa_tree_add_51_79_groupi_n_4180, csa_tree_add_51_79_groupi_n_4181, csa_tree_add_51_79_groupi_n_4182, csa_tree_add_51_79_groupi_n_4183;
  wire csa_tree_add_51_79_groupi_n_4184, csa_tree_add_51_79_groupi_n_4185, csa_tree_add_51_79_groupi_n_4186, csa_tree_add_51_79_groupi_n_4187, csa_tree_add_51_79_groupi_n_4188, csa_tree_add_51_79_groupi_n_4189, csa_tree_add_51_79_groupi_n_4190, csa_tree_add_51_79_groupi_n_4191;
  wire csa_tree_add_51_79_groupi_n_4192, csa_tree_add_51_79_groupi_n_4193, csa_tree_add_51_79_groupi_n_4194, csa_tree_add_51_79_groupi_n_4195, csa_tree_add_51_79_groupi_n_4196, csa_tree_add_51_79_groupi_n_4197, csa_tree_add_51_79_groupi_n_4198, csa_tree_add_51_79_groupi_n_4199;
  wire csa_tree_add_51_79_groupi_n_4200, csa_tree_add_51_79_groupi_n_4201, csa_tree_add_51_79_groupi_n_4202, csa_tree_add_51_79_groupi_n_4203, csa_tree_add_51_79_groupi_n_4204, csa_tree_add_51_79_groupi_n_4205, csa_tree_add_51_79_groupi_n_4206, csa_tree_add_51_79_groupi_n_4207;
  wire csa_tree_add_51_79_groupi_n_4208, csa_tree_add_51_79_groupi_n_4209, csa_tree_add_51_79_groupi_n_4210, csa_tree_add_51_79_groupi_n_4211, csa_tree_add_51_79_groupi_n_4212, csa_tree_add_51_79_groupi_n_4213, csa_tree_add_51_79_groupi_n_4214, csa_tree_add_51_79_groupi_n_4215;
  wire csa_tree_add_51_79_groupi_n_4216, csa_tree_add_51_79_groupi_n_4217, csa_tree_add_51_79_groupi_n_4218, csa_tree_add_51_79_groupi_n_4219, csa_tree_add_51_79_groupi_n_4220, csa_tree_add_51_79_groupi_n_4221, csa_tree_add_51_79_groupi_n_4222, csa_tree_add_51_79_groupi_n_4223;
  wire csa_tree_add_51_79_groupi_n_4224, csa_tree_add_51_79_groupi_n_4225, csa_tree_add_51_79_groupi_n_4226, csa_tree_add_51_79_groupi_n_4227, csa_tree_add_51_79_groupi_n_4228, csa_tree_add_51_79_groupi_n_4229, csa_tree_add_51_79_groupi_n_4230, csa_tree_add_51_79_groupi_n_4231;
  wire csa_tree_add_51_79_groupi_n_4232, csa_tree_add_51_79_groupi_n_4233, csa_tree_add_51_79_groupi_n_4234, csa_tree_add_51_79_groupi_n_4235, csa_tree_add_51_79_groupi_n_4236, csa_tree_add_51_79_groupi_n_4237, csa_tree_add_51_79_groupi_n_4238, csa_tree_add_51_79_groupi_n_4239;
  wire csa_tree_add_51_79_groupi_n_4240, csa_tree_add_51_79_groupi_n_4241, csa_tree_add_51_79_groupi_n_4242, csa_tree_add_51_79_groupi_n_4243, csa_tree_add_51_79_groupi_n_4244, csa_tree_add_51_79_groupi_n_4245, csa_tree_add_51_79_groupi_n_4246, csa_tree_add_51_79_groupi_n_4247;
  wire csa_tree_add_51_79_groupi_n_4248, csa_tree_add_51_79_groupi_n_4249, csa_tree_add_51_79_groupi_n_4250, csa_tree_add_51_79_groupi_n_4251, csa_tree_add_51_79_groupi_n_4252, csa_tree_add_51_79_groupi_n_4253, csa_tree_add_51_79_groupi_n_4254, csa_tree_add_51_79_groupi_n_4255;
  wire csa_tree_add_51_79_groupi_n_4256, csa_tree_add_51_79_groupi_n_4257, csa_tree_add_51_79_groupi_n_4258, csa_tree_add_51_79_groupi_n_4259, csa_tree_add_51_79_groupi_n_4260, csa_tree_add_51_79_groupi_n_4261, csa_tree_add_51_79_groupi_n_4262, csa_tree_add_51_79_groupi_n_4263;
  wire csa_tree_add_51_79_groupi_n_4264, csa_tree_add_51_79_groupi_n_4265, csa_tree_add_51_79_groupi_n_4266, csa_tree_add_51_79_groupi_n_4267, csa_tree_add_51_79_groupi_n_4268, csa_tree_add_51_79_groupi_n_4269, csa_tree_add_51_79_groupi_n_4270, csa_tree_add_51_79_groupi_n_4271;
  wire csa_tree_add_51_79_groupi_n_4272, csa_tree_add_51_79_groupi_n_4273, csa_tree_add_51_79_groupi_n_4274, csa_tree_add_51_79_groupi_n_4275, csa_tree_add_51_79_groupi_n_4276, csa_tree_add_51_79_groupi_n_4277, csa_tree_add_51_79_groupi_n_4278, csa_tree_add_51_79_groupi_n_4279;
  wire csa_tree_add_51_79_groupi_n_4280, csa_tree_add_51_79_groupi_n_4281, csa_tree_add_51_79_groupi_n_4282, csa_tree_add_51_79_groupi_n_4283, csa_tree_add_51_79_groupi_n_4284, csa_tree_add_51_79_groupi_n_4285, csa_tree_add_51_79_groupi_n_4286, csa_tree_add_51_79_groupi_n_4287;
  wire csa_tree_add_51_79_groupi_n_4288, csa_tree_add_51_79_groupi_n_4289, csa_tree_add_51_79_groupi_n_4290, csa_tree_add_51_79_groupi_n_4291, csa_tree_add_51_79_groupi_n_4292, csa_tree_add_51_79_groupi_n_4293, csa_tree_add_51_79_groupi_n_4294, csa_tree_add_51_79_groupi_n_4295;
  wire csa_tree_add_51_79_groupi_n_4296, csa_tree_add_51_79_groupi_n_4297, csa_tree_add_51_79_groupi_n_4298, csa_tree_add_51_79_groupi_n_4299, csa_tree_add_51_79_groupi_n_4300, csa_tree_add_51_79_groupi_n_4301, csa_tree_add_51_79_groupi_n_4302, csa_tree_add_51_79_groupi_n_4303;
  wire csa_tree_add_51_79_groupi_n_4304, csa_tree_add_51_79_groupi_n_4305, csa_tree_add_51_79_groupi_n_4306, csa_tree_add_51_79_groupi_n_4307, csa_tree_add_51_79_groupi_n_4308, csa_tree_add_51_79_groupi_n_4309, csa_tree_add_51_79_groupi_n_4310, csa_tree_add_51_79_groupi_n_4311;
  wire csa_tree_add_51_79_groupi_n_4312, csa_tree_add_51_79_groupi_n_4313, csa_tree_add_51_79_groupi_n_4314, csa_tree_add_51_79_groupi_n_4315, csa_tree_add_51_79_groupi_n_4316, csa_tree_add_51_79_groupi_n_4317, csa_tree_add_51_79_groupi_n_4318, csa_tree_add_51_79_groupi_n_4319;
  wire csa_tree_add_51_79_groupi_n_4320, csa_tree_add_51_79_groupi_n_4321, csa_tree_add_51_79_groupi_n_4322, csa_tree_add_51_79_groupi_n_4323, csa_tree_add_51_79_groupi_n_4324, csa_tree_add_51_79_groupi_n_4325, csa_tree_add_51_79_groupi_n_4326, csa_tree_add_51_79_groupi_n_4327;
  wire csa_tree_add_51_79_groupi_n_4328, csa_tree_add_51_79_groupi_n_4329, csa_tree_add_51_79_groupi_n_4330, csa_tree_add_51_79_groupi_n_4331, csa_tree_add_51_79_groupi_n_4332, csa_tree_add_51_79_groupi_n_4333, csa_tree_add_51_79_groupi_n_4334, csa_tree_add_51_79_groupi_n_4335;
  wire csa_tree_add_51_79_groupi_n_4336, csa_tree_add_51_79_groupi_n_4337, csa_tree_add_51_79_groupi_n_4338, csa_tree_add_51_79_groupi_n_4339, csa_tree_add_51_79_groupi_n_4340, csa_tree_add_51_79_groupi_n_4341, csa_tree_add_51_79_groupi_n_4342, csa_tree_add_51_79_groupi_n_4343;
  wire csa_tree_add_51_79_groupi_n_4344, csa_tree_add_51_79_groupi_n_4345, csa_tree_add_51_79_groupi_n_4346, csa_tree_add_51_79_groupi_n_4347, csa_tree_add_51_79_groupi_n_4348, csa_tree_add_51_79_groupi_n_4349, csa_tree_add_51_79_groupi_n_4350, csa_tree_add_51_79_groupi_n_4351;
  wire csa_tree_add_51_79_groupi_n_4352, csa_tree_add_51_79_groupi_n_4353, csa_tree_add_51_79_groupi_n_4354, csa_tree_add_51_79_groupi_n_4355, csa_tree_add_51_79_groupi_n_4356, csa_tree_add_51_79_groupi_n_4357, csa_tree_add_51_79_groupi_n_4358, csa_tree_add_51_79_groupi_n_4359;
  wire csa_tree_add_51_79_groupi_n_4360, csa_tree_add_51_79_groupi_n_4361, csa_tree_add_51_79_groupi_n_4362, csa_tree_add_51_79_groupi_n_4363, csa_tree_add_51_79_groupi_n_4364, csa_tree_add_51_79_groupi_n_4365, csa_tree_add_51_79_groupi_n_4366, csa_tree_add_51_79_groupi_n_4367;
  wire csa_tree_add_51_79_groupi_n_4368, csa_tree_add_51_79_groupi_n_4369, csa_tree_add_51_79_groupi_n_4370, csa_tree_add_51_79_groupi_n_4371, csa_tree_add_51_79_groupi_n_4372, csa_tree_add_51_79_groupi_n_4373, csa_tree_add_51_79_groupi_n_4374, csa_tree_add_51_79_groupi_n_4375;
  wire csa_tree_add_51_79_groupi_n_4376, csa_tree_add_51_79_groupi_n_4377, csa_tree_add_51_79_groupi_n_4378, csa_tree_add_51_79_groupi_n_4379, csa_tree_add_51_79_groupi_n_4380, csa_tree_add_51_79_groupi_n_4381, csa_tree_add_51_79_groupi_n_4382, csa_tree_add_51_79_groupi_n_4383;
  wire csa_tree_add_51_79_groupi_n_4384, csa_tree_add_51_79_groupi_n_4385, csa_tree_add_51_79_groupi_n_4386, csa_tree_add_51_79_groupi_n_4387, csa_tree_add_51_79_groupi_n_4388, csa_tree_add_51_79_groupi_n_4389, csa_tree_add_51_79_groupi_n_4390, csa_tree_add_51_79_groupi_n_4391;
  wire csa_tree_add_51_79_groupi_n_4392, csa_tree_add_51_79_groupi_n_4393, csa_tree_add_51_79_groupi_n_4394, csa_tree_add_51_79_groupi_n_4395, csa_tree_add_51_79_groupi_n_4396, csa_tree_add_51_79_groupi_n_4397, csa_tree_add_51_79_groupi_n_4398, csa_tree_add_51_79_groupi_n_4399;
  wire csa_tree_add_51_79_groupi_n_4400, csa_tree_add_51_79_groupi_n_4401, csa_tree_add_51_79_groupi_n_4402, csa_tree_add_51_79_groupi_n_4403, csa_tree_add_51_79_groupi_n_4404, csa_tree_add_51_79_groupi_n_4405, csa_tree_add_51_79_groupi_n_4406, csa_tree_add_51_79_groupi_n_4407;
  wire csa_tree_add_51_79_groupi_n_4408, csa_tree_add_51_79_groupi_n_4409, csa_tree_add_51_79_groupi_n_4410, csa_tree_add_51_79_groupi_n_4411, csa_tree_add_51_79_groupi_n_4412, csa_tree_add_51_79_groupi_n_4413, csa_tree_add_51_79_groupi_n_4414, csa_tree_add_51_79_groupi_n_4415;
  wire csa_tree_add_51_79_groupi_n_4416, csa_tree_add_51_79_groupi_n_4417, csa_tree_add_51_79_groupi_n_4418, csa_tree_add_51_79_groupi_n_4419, csa_tree_add_51_79_groupi_n_4420, csa_tree_add_51_79_groupi_n_4421, csa_tree_add_51_79_groupi_n_4422, csa_tree_add_51_79_groupi_n_4423;
  wire csa_tree_add_51_79_groupi_n_4424, csa_tree_add_51_79_groupi_n_4425, csa_tree_add_51_79_groupi_n_4426, csa_tree_add_51_79_groupi_n_4427, csa_tree_add_51_79_groupi_n_4428, csa_tree_add_51_79_groupi_n_4429, csa_tree_add_51_79_groupi_n_4430, csa_tree_add_51_79_groupi_n_4431;
  wire csa_tree_add_51_79_groupi_n_4432, csa_tree_add_51_79_groupi_n_4433, csa_tree_add_51_79_groupi_n_4434, csa_tree_add_51_79_groupi_n_4435, csa_tree_add_51_79_groupi_n_4436, csa_tree_add_51_79_groupi_n_4437, csa_tree_add_51_79_groupi_n_4438, csa_tree_add_51_79_groupi_n_4439;
  wire csa_tree_add_51_79_groupi_n_4440, csa_tree_add_51_79_groupi_n_4441, csa_tree_add_51_79_groupi_n_4442, csa_tree_add_51_79_groupi_n_4443, csa_tree_add_51_79_groupi_n_4444, csa_tree_add_51_79_groupi_n_4445, csa_tree_add_51_79_groupi_n_4446, csa_tree_add_51_79_groupi_n_4447;
  wire csa_tree_add_51_79_groupi_n_4448, csa_tree_add_51_79_groupi_n_4449, csa_tree_add_51_79_groupi_n_4450, csa_tree_add_51_79_groupi_n_4451, csa_tree_add_51_79_groupi_n_4452, csa_tree_add_51_79_groupi_n_4453, csa_tree_add_51_79_groupi_n_4454, csa_tree_add_51_79_groupi_n_4455;
  wire csa_tree_add_51_79_groupi_n_4456, csa_tree_add_51_79_groupi_n_4457, csa_tree_add_51_79_groupi_n_4458, csa_tree_add_51_79_groupi_n_4459, csa_tree_add_51_79_groupi_n_4460, csa_tree_add_51_79_groupi_n_4461, csa_tree_add_51_79_groupi_n_4462, csa_tree_add_51_79_groupi_n_4463;
  wire csa_tree_add_51_79_groupi_n_4464, csa_tree_add_51_79_groupi_n_4465, csa_tree_add_51_79_groupi_n_4466, csa_tree_add_51_79_groupi_n_4467, csa_tree_add_51_79_groupi_n_4468, csa_tree_add_51_79_groupi_n_4469, csa_tree_add_51_79_groupi_n_4470, csa_tree_add_51_79_groupi_n_4471;
  wire csa_tree_add_51_79_groupi_n_4472, csa_tree_add_51_79_groupi_n_4473, csa_tree_add_51_79_groupi_n_4474, csa_tree_add_51_79_groupi_n_4475, csa_tree_add_51_79_groupi_n_4476, csa_tree_add_51_79_groupi_n_4477, csa_tree_add_51_79_groupi_n_4478, csa_tree_add_51_79_groupi_n_4479;
  wire csa_tree_add_51_79_groupi_n_4480, csa_tree_add_51_79_groupi_n_4481, csa_tree_add_51_79_groupi_n_4482, csa_tree_add_51_79_groupi_n_4483, csa_tree_add_51_79_groupi_n_4484, csa_tree_add_51_79_groupi_n_4485, csa_tree_add_51_79_groupi_n_4486, csa_tree_add_51_79_groupi_n_4487;
  wire csa_tree_add_51_79_groupi_n_4488, csa_tree_add_51_79_groupi_n_4489, csa_tree_add_51_79_groupi_n_4490, csa_tree_add_51_79_groupi_n_4491, csa_tree_add_51_79_groupi_n_4492, csa_tree_add_51_79_groupi_n_4493, csa_tree_add_51_79_groupi_n_4494, csa_tree_add_51_79_groupi_n_4495;
  wire csa_tree_add_51_79_groupi_n_4496, csa_tree_add_51_79_groupi_n_4497, csa_tree_add_51_79_groupi_n_4498, csa_tree_add_51_79_groupi_n_4499, csa_tree_add_51_79_groupi_n_4500, csa_tree_add_51_79_groupi_n_4501, csa_tree_add_51_79_groupi_n_4502, csa_tree_add_51_79_groupi_n_4503;
  wire csa_tree_add_51_79_groupi_n_4504, csa_tree_add_51_79_groupi_n_4505, csa_tree_add_51_79_groupi_n_4506, csa_tree_add_51_79_groupi_n_4507, csa_tree_add_51_79_groupi_n_4508, csa_tree_add_51_79_groupi_n_4509, csa_tree_add_51_79_groupi_n_4510, csa_tree_add_51_79_groupi_n_4511;
  wire csa_tree_add_51_79_groupi_n_4512, csa_tree_add_51_79_groupi_n_4513, csa_tree_add_51_79_groupi_n_4514, csa_tree_add_51_79_groupi_n_4515, csa_tree_add_51_79_groupi_n_4516, csa_tree_add_51_79_groupi_n_4517, csa_tree_add_51_79_groupi_n_4518, csa_tree_add_51_79_groupi_n_4519;
  wire csa_tree_add_51_79_groupi_n_4520, csa_tree_add_51_79_groupi_n_4521, csa_tree_add_51_79_groupi_n_4522, csa_tree_add_51_79_groupi_n_4523, csa_tree_add_51_79_groupi_n_4524, csa_tree_add_51_79_groupi_n_4525, csa_tree_add_51_79_groupi_n_4526, csa_tree_add_51_79_groupi_n_4527;
  wire csa_tree_add_51_79_groupi_n_4528, csa_tree_add_51_79_groupi_n_4529, csa_tree_add_51_79_groupi_n_4530, csa_tree_add_51_79_groupi_n_4531, csa_tree_add_51_79_groupi_n_4532, csa_tree_add_51_79_groupi_n_4533, csa_tree_add_51_79_groupi_n_4534, csa_tree_add_51_79_groupi_n_4535;
  wire csa_tree_add_51_79_groupi_n_4536, csa_tree_add_51_79_groupi_n_4537, csa_tree_add_51_79_groupi_n_4538, csa_tree_add_51_79_groupi_n_4539, csa_tree_add_51_79_groupi_n_4540, csa_tree_add_51_79_groupi_n_4541, csa_tree_add_51_79_groupi_n_4542, csa_tree_add_51_79_groupi_n_4543;
  wire csa_tree_add_51_79_groupi_n_4544, csa_tree_add_51_79_groupi_n_4545, csa_tree_add_51_79_groupi_n_4546, csa_tree_add_51_79_groupi_n_4547, csa_tree_add_51_79_groupi_n_4548, csa_tree_add_51_79_groupi_n_4549, csa_tree_add_51_79_groupi_n_4550, csa_tree_add_51_79_groupi_n_4551;
  wire csa_tree_add_51_79_groupi_n_4552, csa_tree_add_51_79_groupi_n_4553, csa_tree_add_51_79_groupi_n_4554, csa_tree_add_51_79_groupi_n_4555, csa_tree_add_51_79_groupi_n_4556, csa_tree_add_51_79_groupi_n_4557, csa_tree_add_51_79_groupi_n_4558, csa_tree_add_51_79_groupi_n_4559;
  wire csa_tree_add_51_79_groupi_n_4560, csa_tree_add_51_79_groupi_n_4561, csa_tree_add_51_79_groupi_n_4562, csa_tree_add_51_79_groupi_n_4563, csa_tree_add_51_79_groupi_n_4564, csa_tree_add_51_79_groupi_n_4565, csa_tree_add_51_79_groupi_n_4566, csa_tree_add_51_79_groupi_n_4567;
  wire csa_tree_add_51_79_groupi_n_4568, csa_tree_add_51_79_groupi_n_4569, csa_tree_add_51_79_groupi_n_4570, csa_tree_add_51_79_groupi_n_4571, csa_tree_add_51_79_groupi_n_4572, csa_tree_add_51_79_groupi_n_4573, csa_tree_add_51_79_groupi_n_4574, csa_tree_add_51_79_groupi_n_4575;
  wire csa_tree_add_51_79_groupi_n_4576, csa_tree_add_51_79_groupi_n_4577, csa_tree_add_51_79_groupi_n_4578, csa_tree_add_51_79_groupi_n_4579, csa_tree_add_51_79_groupi_n_4580, csa_tree_add_51_79_groupi_n_4581, csa_tree_add_51_79_groupi_n_4582, csa_tree_add_51_79_groupi_n_4583;
  wire csa_tree_add_51_79_groupi_n_4584, csa_tree_add_51_79_groupi_n_4585, csa_tree_add_51_79_groupi_n_4586, csa_tree_add_51_79_groupi_n_4587, csa_tree_add_51_79_groupi_n_4588, csa_tree_add_51_79_groupi_n_4589, csa_tree_add_51_79_groupi_n_4590, csa_tree_add_51_79_groupi_n_4591;
  wire csa_tree_add_51_79_groupi_n_4592, csa_tree_add_51_79_groupi_n_4593, csa_tree_add_51_79_groupi_n_4594, csa_tree_add_51_79_groupi_n_4595, csa_tree_add_51_79_groupi_n_4596, csa_tree_add_51_79_groupi_n_4597, csa_tree_add_51_79_groupi_n_4598, csa_tree_add_51_79_groupi_n_4599;
  wire csa_tree_add_51_79_groupi_n_4600, csa_tree_add_51_79_groupi_n_4601, csa_tree_add_51_79_groupi_n_4602, csa_tree_add_51_79_groupi_n_4603, csa_tree_add_51_79_groupi_n_4604, csa_tree_add_51_79_groupi_n_4605, csa_tree_add_51_79_groupi_n_4606, csa_tree_add_51_79_groupi_n_4607;
  wire csa_tree_add_51_79_groupi_n_4608, csa_tree_add_51_79_groupi_n_4609, csa_tree_add_51_79_groupi_n_4610, csa_tree_add_51_79_groupi_n_4611, csa_tree_add_51_79_groupi_n_4612, csa_tree_add_51_79_groupi_n_4613, csa_tree_add_51_79_groupi_n_4614, csa_tree_add_51_79_groupi_n_4615;
  wire csa_tree_add_51_79_groupi_n_4616, csa_tree_add_51_79_groupi_n_4617, csa_tree_add_51_79_groupi_n_4618, csa_tree_add_51_79_groupi_n_4619, csa_tree_add_51_79_groupi_n_4620, csa_tree_add_51_79_groupi_n_4621, csa_tree_add_51_79_groupi_n_4622, csa_tree_add_51_79_groupi_n_4623;
  wire csa_tree_add_51_79_groupi_n_4624, csa_tree_add_51_79_groupi_n_4625, csa_tree_add_51_79_groupi_n_4626, csa_tree_add_51_79_groupi_n_4627, csa_tree_add_51_79_groupi_n_4628, csa_tree_add_51_79_groupi_n_4629, csa_tree_add_51_79_groupi_n_4630, csa_tree_add_51_79_groupi_n_4631;
  wire csa_tree_add_51_79_groupi_n_4632, csa_tree_add_51_79_groupi_n_4633, csa_tree_add_51_79_groupi_n_4634, csa_tree_add_51_79_groupi_n_4635, csa_tree_add_51_79_groupi_n_4636, csa_tree_add_51_79_groupi_n_4637, csa_tree_add_51_79_groupi_n_4638, csa_tree_add_51_79_groupi_n_4639;
  wire csa_tree_add_51_79_groupi_n_4640, csa_tree_add_51_79_groupi_n_4641, csa_tree_add_51_79_groupi_n_4642, csa_tree_add_51_79_groupi_n_4643, csa_tree_add_51_79_groupi_n_4644, csa_tree_add_51_79_groupi_n_4645, csa_tree_add_51_79_groupi_n_4646, csa_tree_add_51_79_groupi_n_4647;
  wire csa_tree_add_51_79_groupi_n_4648, csa_tree_add_51_79_groupi_n_4649, csa_tree_add_51_79_groupi_n_4650, csa_tree_add_51_79_groupi_n_4651, csa_tree_add_51_79_groupi_n_4652, csa_tree_add_51_79_groupi_n_4653, csa_tree_add_51_79_groupi_n_4654, csa_tree_add_51_79_groupi_n_4655;
  wire csa_tree_add_51_79_groupi_n_4656, csa_tree_add_51_79_groupi_n_4657, csa_tree_add_51_79_groupi_n_4658, csa_tree_add_51_79_groupi_n_4659, csa_tree_add_51_79_groupi_n_4660, csa_tree_add_51_79_groupi_n_4661, csa_tree_add_51_79_groupi_n_4662, csa_tree_add_51_79_groupi_n_4663;
  wire csa_tree_add_51_79_groupi_n_4664, csa_tree_add_51_79_groupi_n_4665, csa_tree_add_51_79_groupi_n_4666, csa_tree_add_51_79_groupi_n_4667, csa_tree_add_51_79_groupi_n_4668, csa_tree_add_51_79_groupi_n_4669, csa_tree_add_51_79_groupi_n_4670, csa_tree_add_51_79_groupi_n_4671;
  wire csa_tree_add_51_79_groupi_n_4672, csa_tree_add_51_79_groupi_n_4673, csa_tree_add_51_79_groupi_n_4674, csa_tree_add_51_79_groupi_n_4675, csa_tree_add_51_79_groupi_n_4676, csa_tree_add_51_79_groupi_n_4677, csa_tree_add_51_79_groupi_n_4678, csa_tree_add_51_79_groupi_n_4679;
  wire csa_tree_add_51_79_groupi_n_4680, csa_tree_add_51_79_groupi_n_4681, csa_tree_add_51_79_groupi_n_4682, csa_tree_add_51_79_groupi_n_4683, csa_tree_add_51_79_groupi_n_4684, csa_tree_add_51_79_groupi_n_4685, csa_tree_add_51_79_groupi_n_4686, csa_tree_add_51_79_groupi_n_4687;
  wire csa_tree_add_51_79_groupi_n_4688, csa_tree_add_51_79_groupi_n_4689, csa_tree_add_51_79_groupi_n_4690, csa_tree_add_51_79_groupi_n_4691, csa_tree_add_51_79_groupi_n_4692, csa_tree_add_51_79_groupi_n_4693, csa_tree_add_51_79_groupi_n_4694, csa_tree_add_51_79_groupi_n_4695;
  wire csa_tree_add_51_79_groupi_n_4696, csa_tree_add_51_79_groupi_n_4697, csa_tree_add_51_79_groupi_n_4698, csa_tree_add_51_79_groupi_n_4699, csa_tree_add_51_79_groupi_n_4700, csa_tree_add_51_79_groupi_n_4701, csa_tree_add_51_79_groupi_n_4702, csa_tree_add_51_79_groupi_n_4703;
  wire csa_tree_add_51_79_groupi_n_4704, csa_tree_add_51_79_groupi_n_4705, csa_tree_add_51_79_groupi_n_4706, csa_tree_add_51_79_groupi_n_4707, csa_tree_add_51_79_groupi_n_4708, csa_tree_add_51_79_groupi_n_4709, csa_tree_add_51_79_groupi_n_4710, csa_tree_add_51_79_groupi_n_4711;
  wire csa_tree_add_51_79_groupi_n_4712, csa_tree_add_51_79_groupi_n_4713, csa_tree_add_51_79_groupi_n_4714, csa_tree_add_51_79_groupi_n_4715, csa_tree_add_51_79_groupi_n_4716, csa_tree_add_51_79_groupi_n_4717, csa_tree_add_51_79_groupi_n_4718, csa_tree_add_51_79_groupi_n_4719;
  wire csa_tree_add_51_79_groupi_n_4720, csa_tree_add_51_79_groupi_n_4721, csa_tree_add_51_79_groupi_n_4722, csa_tree_add_51_79_groupi_n_4723, csa_tree_add_51_79_groupi_n_4724, csa_tree_add_51_79_groupi_n_4725, csa_tree_add_51_79_groupi_n_4726, csa_tree_add_51_79_groupi_n_4727;
  wire csa_tree_add_51_79_groupi_n_4728, csa_tree_add_51_79_groupi_n_4729, csa_tree_add_51_79_groupi_n_4730, csa_tree_add_51_79_groupi_n_4731, csa_tree_add_51_79_groupi_n_4732, csa_tree_add_51_79_groupi_n_4733, csa_tree_add_51_79_groupi_n_4734, csa_tree_add_51_79_groupi_n_4735;
  wire csa_tree_add_51_79_groupi_n_4736, csa_tree_add_51_79_groupi_n_4737, csa_tree_add_51_79_groupi_n_4738, csa_tree_add_51_79_groupi_n_4739, csa_tree_add_51_79_groupi_n_4740, csa_tree_add_51_79_groupi_n_4741, csa_tree_add_51_79_groupi_n_4742, csa_tree_add_51_79_groupi_n_4743;
  wire csa_tree_add_51_79_groupi_n_4744, csa_tree_add_51_79_groupi_n_4745, csa_tree_add_51_79_groupi_n_4746, csa_tree_add_51_79_groupi_n_4747, csa_tree_add_51_79_groupi_n_4748, csa_tree_add_51_79_groupi_n_4749, csa_tree_add_51_79_groupi_n_4750, csa_tree_add_51_79_groupi_n_4751;
  wire csa_tree_add_51_79_groupi_n_4752, csa_tree_add_51_79_groupi_n_4753, csa_tree_add_51_79_groupi_n_4754, csa_tree_add_51_79_groupi_n_4755, csa_tree_add_51_79_groupi_n_4756, csa_tree_add_51_79_groupi_n_4757, csa_tree_add_51_79_groupi_n_4758, csa_tree_add_51_79_groupi_n_4759;
  wire csa_tree_add_51_79_groupi_n_4760, csa_tree_add_51_79_groupi_n_4761, csa_tree_add_51_79_groupi_n_4762, csa_tree_add_51_79_groupi_n_4763, csa_tree_add_51_79_groupi_n_4764, csa_tree_add_51_79_groupi_n_4765, csa_tree_add_51_79_groupi_n_4766, csa_tree_add_51_79_groupi_n_4767;
  wire csa_tree_add_51_79_groupi_n_4768, csa_tree_add_51_79_groupi_n_4769, csa_tree_add_51_79_groupi_n_4770, csa_tree_add_51_79_groupi_n_4771, csa_tree_add_51_79_groupi_n_4772, csa_tree_add_51_79_groupi_n_4773, csa_tree_add_51_79_groupi_n_4774, csa_tree_add_51_79_groupi_n_4775;
  wire csa_tree_add_51_79_groupi_n_4776, csa_tree_add_51_79_groupi_n_4777, csa_tree_add_51_79_groupi_n_4778, csa_tree_add_51_79_groupi_n_4779, csa_tree_add_51_79_groupi_n_4780, csa_tree_add_51_79_groupi_n_4781, csa_tree_add_51_79_groupi_n_4782, csa_tree_add_51_79_groupi_n_4783;
  wire csa_tree_add_51_79_groupi_n_4784, csa_tree_add_51_79_groupi_n_4785, csa_tree_add_51_79_groupi_n_4786, csa_tree_add_51_79_groupi_n_4787, csa_tree_add_51_79_groupi_n_4788, csa_tree_add_51_79_groupi_n_4789, csa_tree_add_51_79_groupi_n_4790, csa_tree_add_51_79_groupi_n_4791;
  wire csa_tree_add_51_79_groupi_n_4792, csa_tree_add_51_79_groupi_n_4793, csa_tree_add_51_79_groupi_n_4794, csa_tree_add_51_79_groupi_n_4795, csa_tree_add_51_79_groupi_n_4796, csa_tree_add_51_79_groupi_n_4797, csa_tree_add_51_79_groupi_n_4798, csa_tree_add_51_79_groupi_n_4799;
  wire csa_tree_add_51_79_groupi_n_4800, csa_tree_add_51_79_groupi_n_4801, csa_tree_add_51_79_groupi_n_4802, csa_tree_add_51_79_groupi_n_4803, csa_tree_add_51_79_groupi_n_4804, csa_tree_add_51_79_groupi_n_4805, csa_tree_add_51_79_groupi_n_4806, csa_tree_add_51_79_groupi_n_4807;
  wire csa_tree_add_51_79_groupi_n_4808, csa_tree_add_51_79_groupi_n_4809, csa_tree_add_51_79_groupi_n_4810, csa_tree_add_51_79_groupi_n_4811, csa_tree_add_51_79_groupi_n_4812, csa_tree_add_51_79_groupi_n_4813, csa_tree_add_51_79_groupi_n_4814, csa_tree_add_51_79_groupi_n_4815;
  wire csa_tree_add_51_79_groupi_n_4816, csa_tree_add_51_79_groupi_n_4817, csa_tree_add_51_79_groupi_n_4818, csa_tree_add_51_79_groupi_n_4819, csa_tree_add_51_79_groupi_n_4820, csa_tree_add_51_79_groupi_n_4821, csa_tree_add_51_79_groupi_n_4822, csa_tree_add_51_79_groupi_n_4823;
  wire csa_tree_add_51_79_groupi_n_4824, csa_tree_add_51_79_groupi_n_4825, csa_tree_add_51_79_groupi_n_4826, csa_tree_add_51_79_groupi_n_4827, csa_tree_add_51_79_groupi_n_4828, csa_tree_add_51_79_groupi_n_4829, csa_tree_add_51_79_groupi_n_4830, csa_tree_add_51_79_groupi_n_4831;
  wire csa_tree_add_51_79_groupi_n_4832, csa_tree_add_51_79_groupi_n_4833, csa_tree_add_51_79_groupi_n_4834, csa_tree_add_51_79_groupi_n_4835, csa_tree_add_51_79_groupi_n_4836, csa_tree_add_51_79_groupi_n_4837, csa_tree_add_51_79_groupi_n_4838, csa_tree_add_51_79_groupi_n_4839;
  wire csa_tree_add_51_79_groupi_n_4840, csa_tree_add_51_79_groupi_n_4841, csa_tree_add_51_79_groupi_n_4842, csa_tree_add_51_79_groupi_n_4843, csa_tree_add_51_79_groupi_n_4844, csa_tree_add_51_79_groupi_n_4845, csa_tree_add_51_79_groupi_n_4846, csa_tree_add_51_79_groupi_n_4847;
  wire csa_tree_add_51_79_groupi_n_4848, csa_tree_add_51_79_groupi_n_4849, csa_tree_add_51_79_groupi_n_4850, csa_tree_add_51_79_groupi_n_4851, csa_tree_add_51_79_groupi_n_4852, csa_tree_add_51_79_groupi_n_4853, csa_tree_add_51_79_groupi_n_4854, csa_tree_add_51_79_groupi_n_4855;
  wire csa_tree_add_51_79_groupi_n_4856, csa_tree_add_51_79_groupi_n_4857, csa_tree_add_51_79_groupi_n_4858, csa_tree_add_51_79_groupi_n_4859, csa_tree_add_51_79_groupi_n_4860, csa_tree_add_51_79_groupi_n_4861, csa_tree_add_51_79_groupi_n_4862, csa_tree_add_51_79_groupi_n_4863;
  wire csa_tree_add_51_79_groupi_n_4864, csa_tree_add_51_79_groupi_n_4865, csa_tree_add_51_79_groupi_n_4866, csa_tree_add_51_79_groupi_n_4867, csa_tree_add_51_79_groupi_n_4868, csa_tree_add_51_79_groupi_n_4869, csa_tree_add_51_79_groupi_n_4870, csa_tree_add_51_79_groupi_n_4871;
  wire csa_tree_add_51_79_groupi_n_4872, csa_tree_add_51_79_groupi_n_4873, csa_tree_add_51_79_groupi_n_4874, csa_tree_add_51_79_groupi_n_4875, csa_tree_add_51_79_groupi_n_4876, csa_tree_add_51_79_groupi_n_4877, csa_tree_add_51_79_groupi_n_4878, csa_tree_add_51_79_groupi_n_4879;
  wire csa_tree_add_51_79_groupi_n_4880, csa_tree_add_51_79_groupi_n_4881, csa_tree_add_51_79_groupi_n_4882, csa_tree_add_51_79_groupi_n_4883, csa_tree_add_51_79_groupi_n_4884, csa_tree_add_51_79_groupi_n_4885, csa_tree_add_51_79_groupi_n_4886, csa_tree_add_51_79_groupi_n_4887;
  wire csa_tree_add_51_79_groupi_n_4888, csa_tree_add_51_79_groupi_n_4889, csa_tree_add_51_79_groupi_n_4890, csa_tree_add_51_79_groupi_n_4891, csa_tree_add_51_79_groupi_n_4892, csa_tree_add_51_79_groupi_n_4893, csa_tree_add_51_79_groupi_n_4894, csa_tree_add_51_79_groupi_n_4895;
  wire csa_tree_add_51_79_groupi_n_4896, csa_tree_add_51_79_groupi_n_4897, csa_tree_add_51_79_groupi_n_4898, csa_tree_add_51_79_groupi_n_4899, csa_tree_add_51_79_groupi_n_4900, csa_tree_add_51_79_groupi_n_4901, csa_tree_add_51_79_groupi_n_4902, csa_tree_add_51_79_groupi_n_4903;
  wire csa_tree_add_51_79_groupi_n_4904, csa_tree_add_51_79_groupi_n_4905, csa_tree_add_51_79_groupi_n_4906, csa_tree_add_51_79_groupi_n_4907, csa_tree_add_51_79_groupi_n_4908, csa_tree_add_51_79_groupi_n_4909, csa_tree_add_51_79_groupi_n_4910, csa_tree_add_51_79_groupi_n_4911;
  wire csa_tree_add_51_79_groupi_n_4912, csa_tree_add_51_79_groupi_n_4913, csa_tree_add_51_79_groupi_n_4914, csa_tree_add_51_79_groupi_n_4915, csa_tree_add_51_79_groupi_n_4916, csa_tree_add_51_79_groupi_n_4917, csa_tree_add_51_79_groupi_n_4918, csa_tree_add_51_79_groupi_n_4919;
  wire csa_tree_add_51_79_groupi_n_4920, csa_tree_add_51_79_groupi_n_4921, csa_tree_add_51_79_groupi_n_4922, csa_tree_add_51_79_groupi_n_4923, csa_tree_add_51_79_groupi_n_4924, csa_tree_add_51_79_groupi_n_4925, csa_tree_add_51_79_groupi_n_4926, csa_tree_add_51_79_groupi_n_4927;
  wire csa_tree_add_51_79_groupi_n_4928, csa_tree_add_51_79_groupi_n_4929, csa_tree_add_51_79_groupi_n_4930, csa_tree_add_51_79_groupi_n_4931, csa_tree_add_51_79_groupi_n_4932, csa_tree_add_51_79_groupi_n_4933, csa_tree_add_51_79_groupi_n_4934, csa_tree_add_51_79_groupi_n_4935;
  wire csa_tree_add_51_79_groupi_n_4936, csa_tree_add_51_79_groupi_n_4937, csa_tree_add_51_79_groupi_n_4938, csa_tree_add_51_79_groupi_n_4939, csa_tree_add_51_79_groupi_n_4940, csa_tree_add_51_79_groupi_n_4941, csa_tree_add_51_79_groupi_n_4942, csa_tree_add_51_79_groupi_n_4943;
  wire csa_tree_add_51_79_groupi_n_4944, csa_tree_add_51_79_groupi_n_4945, csa_tree_add_51_79_groupi_n_4946, csa_tree_add_51_79_groupi_n_4947, csa_tree_add_51_79_groupi_n_4948, csa_tree_add_51_79_groupi_n_4949, csa_tree_add_51_79_groupi_n_4950, csa_tree_add_51_79_groupi_n_4951;
  wire csa_tree_add_51_79_groupi_n_4952, csa_tree_add_51_79_groupi_n_4953, csa_tree_add_51_79_groupi_n_4954, csa_tree_add_51_79_groupi_n_4955, csa_tree_add_51_79_groupi_n_4956, csa_tree_add_51_79_groupi_n_4957, csa_tree_add_51_79_groupi_n_4958, csa_tree_add_51_79_groupi_n_4959;
  wire csa_tree_add_51_79_groupi_n_4960, csa_tree_add_51_79_groupi_n_4961, csa_tree_add_51_79_groupi_n_4962, csa_tree_add_51_79_groupi_n_4963, csa_tree_add_51_79_groupi_n_4964, csa_tree_add_51_79_groupi_n_4965, csa_tree_add_51_79_groupi_n_4966, csa_tree_add_51_79_groupi_n_4967;
  wire csa_tree_add_51_79_groupi_n_4968, csa_tree_add_51_79_groupi_n_4969, csa_tree_add_51_79_groupi_n_4970, csa_tree_add_51_79_groupi_n_4971, csa_tree_add_51_79_groupi_n_4972, csa_tree_add_51_79_groupi_n_4973, csa_tree_add_51_79_groupi_n_4974, csa_tree_add_51_79_groupi_n_4975;
  wire csa_tree_add_51_79_groupi_n_4976, csa_tree_add_51_79_groupi_n_4977, csa_tree_add_51_79_groupi_n_4978, csa_tree_add_51_79_groupi_n_4979, csa_tree_add_51_79_groupi_n_4980, csa_tree_add_51_79_groupi_n_4981, csa_tree_add_51_79_groupi_n_4982, csa_tree_add_51_79_groupi_n_4983;
  wire csa_tree_add_51_79_groupi_n_4984, csa_tree_add_51_79_groupi_n_4985, csa_tree_add_51_79_groupi_n_4986, csa_tree_add_51_79_groupi_n_4987, csa_tree_add_51_79_groupi_n_4988, csa_tree_add_51_79_groupi_n_4989, csa_tree_add_51_79_groupi_n_4990, csa_tree_add_51_79_groupi_n_4991;
  wire csa_tree_add_51_79_groupi_n_4992, csa_tree_add_51_79_groupi_n_4993, csa_tree_add_51_79_groupi_n_4994, csa_tree_add_51_79_groupi_n_4995, csa_tree_add_51_79_groupi_n_4996, csa_tree_add_51_79_groupi_n_4997, csa_tree_add_51_79_groupi_n_4998, csa_tree_add_51_79_groupi_n_4999;
  wire csa_tree_add_51_79_groupi_n_5000, csa_tree_add_51_79_groupi_n_5001, csa_tree_add_51_79_groupi_n_5002, csa_tree_add_51_79_groupi_n_5003, csa_tree_add_51_79_groupi_n_5004, csa_tree_add_51_79_groupi_n_5005, csa_tree_add_51_79_groupi_n_5006, csa_tree_add_51_79_groupi_n_5007;
  wire csa_tree_add_51_79_groupi_n_5008, csa_tree_add_51_79_groupi_n_5009, csa_tree_add_51_79_groupi_n_5010, csa_tree_add_51_79_groupi_n_5011, csa_tree_add_51_79_groupi_n_5012, csa_tree_add_51_79_groupi_n_5013, csa_tree_add_51_79_groupi_n_5014, csa_tree_add_51_79_groupi_n_5015;
  wire csa_tree_add_51_79_groupi_n_5016, csa_tree_add_51_79_groupi_n_5017, csa_tree_add_51_79_groupi_n_5018, csa_tree_add_51_79_groupi_n_5019, csa_tree_add_51_79_groupi_n_5020, csa_tree_add_51_79_groupi_n_5021, csa_tree_add_51_79_groupi_n_5022, csa_tree_add_51_79_groupi_n_5023;
  wire csa_tree_add_51_79_groupi_n_5024, csa_tree_add_51_79_groupi_n_5025, csa_tree_add_51_79_groupi_n_5026, csa_tree_add_51_79_groupi_n_5027, csa_tree_add_51_79_groupi_n_5028, csa_tree_add_51_79_groupi_n_5029, csa_tree_add_51_79_groupi_n_5030, csa_tree_add_51_79_groupi_n_5031;
  wire csa_tree_add_51_79_groupi_n_5032, csa_tree_add_51_79_groupi_n_5033, csa_tree_add_51_79_groupi_n_5034, csa_tree_add_51_79_groupi_n_5035, csa_tree_add_51_79_groupi_n_5036, csa_tree_add_51_79_groupi_n_5037, csa_tree_add_51_79_groupi_n_5038, csa_tree_add_51_79_groupi_n_5039;
  wire csa_tree_add_51_79_groupi_n_5040, csa_tree_add_51_79_groupi_n_5041, csa_tree_add_51_79_groupi_n_5042, csa_tree_add_51_79_groupi_n_5043, csa_tree_add_51_79_groupi_n_5044, csa_tree_add_51_79_groupi_n_5045, csa_tree_add_51_79_groupi_n_5046, csa_tree_add_51_79_groupi_n_5047;
  wire csa_tree_add_51_79_groupi_n_5048, csa_tree_add_51_79_groupi_n_5049, csa_tree_add_51_79_groupi_n_5050, csa_tree_add_51_79_groupi_n_5051, csa_tree_add_51_79_groupi_n_5052, csa_tree_add_51_79_groupi_n_5053, csa_tree_add_51_79_groupi_n_5054, csa_tree_add_51_79_groupi_n_5055;
  wire csa_tree_add_51_79_groupi_n_5056, csa_tree_add_51_79_groupi_n_5057, csa_tree_add_51_79_groupi_n_5058, csa_tree_add_51_79_groupi_n_5059, csa_tree_add_51_79_groupi_n_5060, csa_tree_add_51_79_groupi_n_5061, csa_tree_add_51_79_groupi_n_5062, csa_tree_add_51_79_groupi_n_5063;
  wire csa_tree_add_51_79_groupi_n_5064, csa_tree_add_51_79_groupi_n_5065, csa_tree_add_51_79_groupi_n_5066, csa_tree_add_51_79_groupi_n_5067, csa_tree_add_51_79_groupi_n_5068, csa_tree_add_51_79_groupi_n_5069, csa_tree_add_51_79_groupi_n_5070, csa_tree_add_51_79_groupi_n_5071;
  wire csa_tree_add_51_79_groupi_n_5072, csa_tree_add_51_79_groupi_n_5073, csa_tree_add_51_79_groupi_n_5074, csa_tree_add_51_79_groupi_n_5075, csa_tree_add_51_79_groupi_n_5076, csa_tree_add_51_79_groupi_n_5077, csa_tree_add_51_79_groupi_n_5078, csa_tree_add_51_79_groupi_n_5079;
  wire csa_tree_add_51_79_groupi_n_5080, csa_tree_add_51_79_groupi_n_5081, csa_tree_add_51_79_groupi_n_5082, csa_tree_add_51_79_groupi_n_5083, csa_tree_add_51_79_groupi_n_5084, csa_tree_add_51_79_groupi_n_5085, csa_tree_add_51_79_groupi_n_5086, csa_tree_add_51_79_groupi_n_5087;
  wire csa_tree_add_51_79_groupi_n_5088, csa_tree_add_51_79_groupi_n_5089, csa_tree_add_51_79_groupi_n_5090, csa_tree_add_51_79_groupi_n_5091, csa_tree_add_51_79_groupi_n_5092, csa_tree_add_51_79_groupi_n_5093, csa_tree_add_51_79_groupi_n_5094, csa_tree_add_51_79_groupi_n_5095;
  wire csa_tree_add_51_79_groupi_n_5096, csa_tree_add_51_79_groupi_n_5097, csa_tree_add_51_79_groupi_n_5098, csa_tree_add_51_79_groupi_n_5099, csa_tree_add_51_79_groupi_n_5100, csa_tree_add_51_79_groupi_n_5101, csa_tree_add_51_79_groupi_n_5102, csa_tree_add_51_79_groupi_n_5103;
  wire csa_tree_add_51_79_groupi_n_5104, csa_tree_add_51_79_groupi_n_5105, csa_tree_add_51_79_groupi_n_5106, csa_tree_add_51_79_groupi_n_5107, csa_tree_add_51_79_groupi_n_5108, csa_tree_add_51_79_groupi_n_5109, csa_tree_add_51_79_groupi_n_5110, csa_tree_add_51_79_groupi_n_5111;
  wire csa_tree_add_51_79_groupi_n_5112, csa_tree_add_51_79_groupi_n_5113, csa_tree_add_51_79_groupi_n_5114, csa_tree_add_51_79_groupi_n_5115, csa_tree_add_51_79_groupi_n_5116, csa_tree_add_51_79_groupi_n_5117, csa_tree_add_51_79_groupi_n_5118, csa_tree_add_51_79_groupi_n_5119;
  wire csa_tree_add_51_79_groupi_n_5120, csa_tree_add_51_79_groupi_n_5121, csa_tree_add_51_79_groupi_n_5122, csa_tree_add_51_79_groupi_n_5123, csa_tree_add_51_79_groupi_n_5124, csa_tree_add_51_79_groupi_n_5125, csa_tree_add_51_79_groupi_n_5126, csa_tree_add_51_79_groupi_n_5127;
  wire csa_tree_add_51_79_groupi_n_5128, csa_tree_add_51_79_groupi_n_5129, csa_tree_add_51_79_groupi_n_5130, csa_tree_add_51_79_groupi_n_5131, csa_tree_add_51_79_groupi_n_5132, csa_tree_add_51_79_groupi_n_5133, csa_tree_add_51_79_groupi_n_5134, csa_tree_add_51_79_groupi_n_5135;
  wire csa_tree_add_51_79_groupi_n_5136, csa_tree_add_51_79_groupi_n_5137, csa_tree_add_51_79_groupi_n_5138, csa_tree_add_51_79_groupi_n_5139, csa_tree_add_51_79_groupi_n_5140, csa_tree_add_51_79_groupi_n_5141, csa_tree_add_51_79_groupi_n_5142, csa_tree_add_51_79_groupi_n_5143;
  wire csa_tree_add_51_79_groupi_n_5144, csa_tree_add_51_79_groupi_n_5145, csa_tree_add_51_79_groupi_n_5146, csa_tree_add_51_79_groupi_n_5147, csa_tree_add_51_79_groupi_n_5148, csa_tree_add_51_79_groupi_n_5149, csa_tree_add_51_79_groupi_n_5150, csa_tree_add_51_79_groupi_n_5151;
  wire csa_tree_add_51_79_groupi_n_5152, csa_tree_add_51_79_groupi_n_5153, csa_tree_add_51_79_groupi_n_5154, csa_tree_add_51_79_groupi_n_5155, csa_tree_add_51_79_groupi_n_5156, csa_tree_add_51_79_groupi_n_5157, csa_tree_add_51_79_groupi_n_5158, csa_tree_add_51_79_groupi_n_5159;
  wire csa_tree_add_51_79_groupi_n_5160, csa_tree_add_51_79_groupi_n_5161, csa_tree_add_51_79_groupi_n_5162, csa_tree_add_51_79_groupi_n_5163, csa_tree_add_51_79_groupi_n_5164, csa_tree_add_51_79_groupi_n_5165, csa_tree_add_51_79_groupi_n_5166, csa_tree_add_51_79_groupi_n_5167;
  wire csa_tree_add_51_79_groupi_n_5168, csa_tree_add_51_79_groupi_n_5169, csa_tree_add_51_79_groupi_n_5170, csa_tree_add_51_79_groupi_n_5171, csa_tree_add_51_79_groupi_n_5172, csa_tree_add_51_79_groupi_n_5173, csa_tree_add_51_79_groupi_n_5174, csa_tree_add_51_79_groupi_n_5175;
  wire csa_tree_add_51_79_groupi_n_5176, csa_tree_add_51_79_groupi_n_5177, csa_tree_add_51_79_groupi_n_5178, csa_tree_add_51_79_groupi_n_5179, csa_tree_add_51_79_groupi_n_5180, csa_tree_add_51_79_groupi_n_5181, csa_tree_add_51_79_groupi_n_5182, csa_tree_add_51_79_groupi_n_5183;
  wire csa_tree_add_51_79_groupi_n_5184, csa_tree_add_51_79_groupi_n_5185, csa_tree_add_51_79_groupi_n_5186, csa_tree_add_51_79_groupi_n_5187, csa_tree_add_51_79_groupi_n_5188, csa_tree_add_51_79_groupi_n_5189, csa_tree_add_51_79_groupi_n_5190, csa_tree_add_51_79_groupi_n_5191;
  wire csa_tree_add_51_79_groupi_n_5192, csa_tree_add_51_79_groupi_n_5193, csa_tree_add_51_79_groupi_n_5194, csa_tree_add_51_79_groupi_n_5195, csa_tree_add_51_79_groupi_n_5196, csa_tree_add_51_79_groupi_n_5197, csa_tree_add_51_79_groupi_n_5198, csa_tree_add_51_79_groupi_n_5199;
  wire csa_tree_add_51_79_groupi_n_5200, csa_tree_add_51_79_groupi_n_5201, csa_tree_add_51_79_groupi_n_5202, csa_tree_add_51_79_groupi_n_5203, csa_tree_add_51_79_groupi_n_5204, csa_tree_add_51_79_groupi_n_5205, csa_tree_add_51_79_groupi_n_5206, csa_tree_add_51_79_groupi_n_5207;
  wire csa_tree_add_51_79_groupi_n_5208, csa_tree_add_51_79_groupi_n_5209, csa_tree_add_51_79_groupi_n_5210, csa_tree_add_51_79_groupi_n_5211, csa_tree_add_51_79_groupi_n_5212, csa_tree_add_51_79_groupi_n_5213, csa_tree_add_51_79_groupi_n_5214, csa_tree_add_51_79_groupi_n_5215;
  wire csa_tree_add_51_79_groupi_n_5216, csa_tree_add_51_79_groupi_n_5217, csa_tree_add_51_79_groupi_n_5218, csa_tree_add_51_79_groupi_n_5219, csa_tree_add_51_79_groupi_n_5220, csa_tree_add_51_79_groupi_n_5221, csa_tree_add_51_79_groupi_n_5222, csa_tree_add_51_79_groupi_n_5223;
  wire csa_tree_add_51_79_groupi_n_5224, csa_tree_add_51_79_groupi_n_5225, csa_tree_add_51_79_groupi_n_5226, csa_tree_add_51_79_groupi_n_5227, csa_tree_add_51_79_groupi_n_5228, csa_tree_add_51_79_groupi_n_5229, csa_tree_add_51_79_groupi_n_5230, csa_tree_add_51_79_groupi_n_5231;
  wire csa_tree_add_51_79_groupi_n_5232, csa_tree_add_51_79_groupi_n_5233, csa_tree_add_51_79_groupi_n_5234, csa_tree_add_51_79_groupi_n_5235, csa_tree_add_51_79_groupi_n_5236, csa_tree_add_51_79_groupi_n_5237, csa_tree_add_51_79_groupi_n_5238, csa_tree_add_51_79_groupi_n_5239;
  wire csa_tree_add_51_79_groupi_n_5240, csa_tree_add_51_79_groupi_n_5241, csa_tree_add_51_79_groupi_n_5242, csa_tree_add_51_79_groupi_n_5243, csa_tree_add_51_79_groupi_n_5244, csa_tree_add_51_79_groupi_n_5245, csa_tree_add_51_79_groupi_n_5246, csa_tree_add_51_79_groupi_n_5247;
  wire csa_tree_add_51_79_groupi_n_5248, csa_tree_add_51_79_groupi_n_5249, csa_tree_add_51_79_groupi_n_5250, csa_tree_add_51_79_groupi_n_5251, csa_tree_add_51_79_groupi_n_5252, csa_tree_add_51_79_groupi_n_5253, csa_tree_add_51_79_groupi_n_5254, csa_tree_add_51_79_groupi_n_5255;
  wire csa_tree_add_51_79_groupi_n_5256, csa_tree_add_51_79_groupi_n_5257, csa_tree_add_51_79_groupi_n_5258, csa_tree_add_51_79_groupi_n_5259, csa_tree_add_51_79_groupi_n_5260, csa_tree_add_51_79_groupi_n_5261, csa_tree_add_51_79_groupi_n_5262, csa_tree_add_51_79_groupi_n_5263;
  wire csa_tree_add_51_79_groupi_n_5264, csa_tree_add_51_79_groupi_n_5265, csa_tree_add_51_79_groupi_n_5266, csa_tree_add_51_79_groupi_n_5267, csa_tree_add_51_79_groupi_n_5268, csa_tree_add_51_79_groupi_n_5269, csa_tree_add_51_79_groupi_n_5270, csa_tree_add_51_79_groupi_n_5271;
  wire csa_tree_add_51_79_groupi_n_5272, csa_tree_add_51_79_groupi_n_5273, csa_tree_add_51_79_groupi_n_5274, csa_tree_add_51_79_groupi_n_5275, csa_tree_add_51_79_groupi_n_5276, csa_tree_add_51_79_groupi_n_5277, csa_tree_add_51_79_groupi_n_5278, csa_tree_add_51_79_groupi_n_5279;
  wire csa_tree_add_51_79_groupi_n_5280, csa_tree_add_51_79_groupi_n_5281, csa_tree_add_51_79_groupi_n_5282, csa_tree_add_51_79_groupi_n_5283, csa_tree_add_51_79_groupi_n_5284, csa_tree_add_51_79_groupi_n_5285, csa_tree_add_51_79_groupi_n_5286, csa_tree_add_51_79_groupi_n_5287;
  wire csa_tree_add_51_79_groupi_n_5288, csa_tree_add_51_79_groupi_n_5289, csa_tree_add_51_79_groupi_n_5290, csa_tree_add_51_79_groupi_n_5291, csa_tree_add_51_79_groupi_n_5292, csa_tree_add_51_79_groupi_n_5293, csa_tree_add_51_79_groupi_n_5294, csa_tree_add_51_79_groupi_n_5295;
  wire csa_tree_add_51_79_groupi_n_5296, csa_tree_add_51_79_groupi_n_5297, csa_tree_add_51_79_groupi_n_5298, csa_tree_add_51_79_groupi_n_5299, csa_tree_add_51_79_groupi_n_5300, csa_tree_add_51_79_groupi_n_5301, csa_tree_add_51_79_groupi_n_5302, csa_tree_add_51_79_groupi_n_5303;
  wire csa_tree_add_51_79_groupi_n_5304, csa_tree_add_51_79_groupi_n_5305, csa_tree_add_51_79_groupi_n_5306, csa_tree_add_51_79_groupi_n_5307, csa_tree_add_51_79_groupi_n_5308, csa_tree_add_51_79_groupi_n_5309, csa_tree_add_51_79_groupi_n_5310, csa_tree_add_51_79_groupi_n_5311;
  wire csa_tree_add_51_79_groupi_n_5312, csa_tree_add_51_79_groupi_n_5313, csa_tree_add_51_79_groupi_n_5314, csa_tree_add_51_79_groupi_n_5315, csa_tree_add_51_79_groupi_n_5316, csa_tree_add_51_79_groupi_n_5317, csa_tree_add_51_79_groupi_n_5318, csa_tree_add_51_79_groupi_n_5319;
  wire csa_tree_add_51_79_groupi_n_5320, csa_tree_add_51_79_groupi_n_5321, csa_tree_add_51_79_groupi_n_5322, csa_tree_add_51_79_groupi_n_5323, csa_tree_add_51_79_groupi_n_5324, csa_tree_add_51_79_groupi_n_5325, csa_tree_add_51_79_groupi_n_5326, csa_tree_add_51_79_groupi_n_5327;
  wire csa_tree_add_51_79_groupi_n_5328, csa_tree_add_51_79_groupi_n_5329, csa_tree_add_51_79_groupi_n_5330, csa_tree_add_51_79_groupi_n_5331, csa_tree_add_51_79_groupi_n_5332, csa_tree_add_51_79_groupi_n_5333, csa_tree_add_51_79_groupi_n_5334, csa_tree_add_51_79_groupi_n_5335;
  wire csa_tree_add_51_79_groupi_n_5336, csa_tree_add_51_79_groupi_n_5337, csa_tree_add_51_79_groupi_n_5338, csa_tree_add_51_79_groupi_n_5339, csa_tree_add_51_79_groupi_n_5340, csa_tree_add_51_79_groupi_n_5341, csa_tree_add_51_79_groupi_n_5342, csa_tree_add_51_79_groupi_n_5343;
  wire csa_tree_add_51_79_groupi_n_5344, csa_tree_add_51_79_groupi_n_5345, csa_tree_add_51_79_groupi_n_5346, csa_tree_add_51_79_groupi_n_5347, csa_tree_add_51_79_groupi_n_5348, csa_tree_add_51_79_groupi_n_5349, csa_tree_add_51_79_groupi_n_5350, csa_tree_add_51_79_groupi_n_5351;
  wire csa_tree_add_51_79_groupi_n_5352, csa_tree_add_51_79_groupi_n_5353, csa_tree_add_51_79_groupi_n_5354, csa_tree_add_51_79_groupi_n_5355, csa_tree_add_51_79_groupi_n_5356, csa_tree_add_51_79_groupi_n_5357, csa_tree_add_51_79_groupi_n_5358, csa_tree_add_51_79_groupi_n_5359;
  wire csa_tree_add_51_79_groupi_n_5360, csa_tree_add_51_79_groupi_n_5361, csa_tree_add_51_79_groupi_n_5362, csa_tree_add_51_79_groupi_n_5363, csa_tree_add_51_79_groupi_n_5364, csa_tree_add_51_79_groupi_n_5365, csa_tree_add_51_79_groupi_n_5366, csa_tree_add_51_79_groupi_n_5367;
  wire csa_tree_add_51_79_groupi_n_5368, csa_tree_add_51_79_groupi_n_5369, csa_tree_add_51_79_groupi_n_5370, csa_tree_add_51_79_groupi_n_5371, csa_tree_add_51_79_groupi_n_5372, csa_tree_add_51_79_groupi_n_5373, csa_tree_add_51_79_groupi_n_5374, csa_tree_add_51_79_groupi_n_5375;
  wire csa_tree_add_51_79_groupi_n_5376, csa_tree_add_51_79_groupi_n_5377, csa_tree_add_51_79_groupi_n_5378, csa_tree_add_51_79_groupi_n_5379, csa_tree_add_51_79_groupi_n_5380, csa_tree_add_51_79_groupi_n_5381, csa_tree_add_51_79_groupi_n_5382, csa_tree_add_51_79_groupi_n_5383;
  wire csa_tree_add_51_79_groupi_n_5384, csa_tree_add_51_79_groupi_n_5385, csa_tree_add_51_79_groupi_n_5386, csa_tree_add_51_79_groupi_n_5387, csa_tree_add_51_79_groupi_n_5388, csa_tree_add_51_79_groupi_n_5389, csa_tree_add_51_79_groupi_n_5390, csa_tree_add_51_79_groupi_n_5391;
  wire csa_tree_add_51_79_groupi_n_5392, csa_tree_add_51_79_groupi_n_5393, csa_tree_add_51_79_groupi_n_5394, csa_tree_add_51_79_groupi_n_5395, csa_tree_add_51_79_groupi_n_5396, csa_tree_add_51_79_groupi_n_5397, csa_tree_add_51_79_groupi_n_5398, csa_tree_add_51_79_groupi_n_5399;
  wire csa_tree_add_51_79_groupi_n_5400, csa_tree_add_51_79_groupi_n_5401, csa_tree_add_51_79_groupi_n_5402, csa_tree_add_51_79_groupi_n_5403, csa_tree_add_51_79_groupi_n_5404, csa_tree_add_51_79_groupi_n_5405, csa_tree_add_51_79_groupi_n_5406, csa_tree_add_51_79_groupi_n_5407;
  wire csa_tree_add_51_79_groupi_n_5408, csa_tree_add_51_79_groupi_n_5409, csa_tree_add_51_79_groupi_n_5410, csa_tree_add_51_79_groupi_n_5411, csa_tree_add_51_79_groupi_n_5412, csa_tree_add_51_79_groupi_n_5413, csa_tree_add_51_79_groupi_n_5414, csa_tree_add_51_79_groupi_n_5415;
  wire csa_tree_add_51_79_groupi_n_5416, csa_tree_add_51_79_groupi_n_5417, csa_tree_add_51_79_groupi_n_5418, csa_tree_add_51_79_groupi_n_5419, csa_tree_add_51_79_groupi_n_5420, csa_tree_add_51_79_groupi_n_5421, csa_tree_add_51_79_groupi_n_5422, csa_tree_add_51_79_groupi_n_5423;
  wire csa_tree_add_51_79_groupi_n_5424, csa_tree_add_51_79_groupi_n_5425, csa_tree_add_51_79_groupi_n_5426, csa_tree_add_51_79_groupi_n_5427, csa_tree_add_51_79_groupi_n_5428, csa_tree_add_51_79_groupi_n_5429, csa_tree_add_51_79_groupi_n_5430, csa_tree_add_51_79_groupi_n_5431;
  wire csa_tree_add_51_79_groupi_n_5432, csa_tree_add_51_79_groupi_n_5433, csa_tree_add_51_79_groupi_n_5434, csa_tree_add_51_79_groupi_n_5435, csa_tree_add_51_79_groupi_n_5436, csa_tree_add_51_79_groupi_n_5437, csa_tree_add_51_79_groupi_n_5438, csa_tree_add_51_79_groupi_n_5439;
  wire csa_tree_add_51_79_groupi_n_5440, csa_tree_add_51_79_groupi_n_5441, csa_tree_add_51_79_groupi_n_5442, csa_tree_add_51_79_groupi_n_5443, csa_tree_add_51_79_groupi_n_5444, csa_tree_add_51_79_groupi_n_5445, csa_tree_add_51_79_groupi_n_5446, csa_tree_add_51_79_groupi_n_5447;
  wire csa_tree_add_51_79_groupi_n_5448, csa_tree_add_51_79_groupi_n_5449, csa_tree_add_51_79_groupi_n_5450, csa_tree_add_51_79_groupi_n_5451, csa_tree_add_51_79_groupi_n_5452, csa_tree_add_51_79_groupi_n_5453, csa_tree_add_51_79_groupi_n_5454, csa_tree_add_51_79_groupi_n_5455;
  wire csa_tree_add_51_79_groupi_n_5456, csa_tree_add_51_79_groupi_n_5457, csa_tree_add_51_79_groupi_n_5458, csa_tree_add_51_79_groupi_n_5459, csa_tree_add_51_79_groupi_n_5460, csa_tree_add_51_79_groupi_n_5461, csa_tree_add_51_79_groupi_n_5462, csa_tree_add_51_79_groupi_n_5463;
  wire csa_tree_add_51_79_groupi_n_5464, csa_tree_add_51_79_groupi_n_5465, csa_tree_add_51_79_groupi_n_5466, csa_tree_add_51_79_groupi_n_5467, csa_tree_add_51_79_groupi_n_5468, csa_tree_add_51_79_groupi_n_5469, csa_tree_add_51_79_groupi_n_5470, csa_tree_add_51_79_groupi_n_5471;
  wire csa_tree_add_51_79_groupi_n_5472, csa_tree_add_51_79_groupi_n_5473, csa_tree_add_51_79_groupi_n_5474, csa_tree_add_51_79_groupi_n_5475, csa_tree_add_51_79_groupi_n_5476, csa_tree_add_51_79_groupi_n_5477, csa_tree_add_51_79_groupi_n_5478, csa_tree_add_51_79_groupi_n_5479;
  wire csa_tree_add_51_79_groupi_n_5480, csa_tree_add_51_79_groupi_n_5481, csa_tree_add_51_79_groupi_n_5482, csa_tree_add_51_79_groupi_n_5483, csa_tree_add_51_79_groupi_n_5484, csa_tree_add_51_79_groupi_n_5485, csa_tree_add_51_79_groupi_n_5486, csa_tree_add_51_79_groupi_n_5487;
  wire csa_tree_add_51_79_groupi_n_5488, csa_tree_add_51_79_groupi_n_5489, csa_tree_add_51_79_groupi_n_5490, csa_tree_add_51_79_groupi_n_5491, csa_tree_add_51_79_groupi_n_5492, csa_tree_add_51_79_groupi_n_5493, csa_tree_add_51_79_groupi_n_5494, csa_tree_add_51_79_groupi_n_5495;
  wire csa_tree_add_51_79_groupi_n_5496, csa_tree_add_51_79_groupi_n_5497, csa_tree_add_51_79_groupi_n_5498, csa_tree_add_51_79_groupi_n_5499, csa_tree_add_51_79_groupi_n_5500, csa_tree_add_51_79_groupi_n_5501, csa_tree_add_51_79_groupi_n_5502, csa_tree_add_51_79_groupi_n_5503;
  wire csa_tree_add_51_79_groupi_n_5504, csa_tree_add_51_79_groupi_n_5505, csa_tree_add_51_79_groupi_n_5506, csa_tree_add_51_79_groupi_n_5507, csa_tree_add_51_79_groupi_n_5508, csa_tree_add_51_79_groupi_n_5509, csa_tree_add_51_79_groupi_n_5510, csa_tree_add_51_79_groupi_n_5511;
  wire csa_tree_add_51_79_groupi_n_5512, csa_tree_add_51_79_groupi_n_5513, csa_tree_add_51_79_groupi_n_5514, csa_tree_add_51_79_groupi_n_5515, csa_tree_add_51_79_groupi_n_5516, csa_tree_add_51_79_groupi_n_5517, csa_tree_add_51_79_groupi_n_5518, csa_tree_add_51_79_groupi_n_5519;
  wire csa_tree_add_51_79_groupi_n_5520, csa_tree_add_51_79_groupi_n_5521, csa_tree_add_51_79_groupi_n_5522, csa_tree_add_51_79_groupi_n_5523, csa_tree_add_51_79_groupi_n_5524, csa_tree_add_51_79_groupi_n_5525, csa_tree_add_51_79_groupi_n_5526, csa_tree_add_51_79_groupi_n_5527;
  wire csa_tree_add_51_79_groupi_n_5528, csa_tree_add_51_79_groupi_n_5529, csa_tree_add_51_79_groupi_n_5530, csa_tree_add_51_79_groupi_n_5531, csa_tree_add_51_79_groupi_n_5532, csa_tree_add_51_79_groupi_n_5533, csa_tree_add_51_79_groupi_n_5534, csa_tree_add_51_79_groupi_n_5535;
  wire csa_tree_add_51_79_groupi_n_5536, csa_tree_add_51_79_groupi_n_5537, csa_tree_add_51_79_groupi_n_5538, csa_tree_add_51_79_groupi_n_5539, csa_tree_add_51_79_groupi_n_5540, csa_tree_add_51_79_groupi_n_5541, csa_tree_add_51_79_groupi_n_5542, csa_tree_add_51_79_groupi_n_5543;
  wire csa_tree_add_51_79_groupi_n_5544, csa_tree_add_51_79_groupi_n_5545, csa_tree_add_51_79_groupi_n_5546, csa_tree_add_51_79_groupi_n_5547, csa_tree_add_51_79_groupi_n_5548, csa_tree_add_51_79_groupi_n_5549, csa_tree_add_51_79_groupi_n_5550, csa_tree_add_51_79_groupi_n_5551;
  wire csa_tree_add_51_79_groupi_n_5552, csa_tree_add_51_79_groupi_n_5553, csa_tree_add_51_79_groupi_n_5554, csa_tree_add_51_79_groupi_n_5555, csa_tree_add_51_79_groupi_n_5556, csa_tree_add_51_79_groupi_n_5557, csa_tree_add_51_79_groupi_n_5558, csa_tree_add_51_79_groupi_n_5559;
  wire csa_tree_add_51_79_groupi_n_5560, csa_tree_add_51_79_groupi_n_5561, csa_tree_add_51_79_groupi_n_5562, csa_tree_add_51_79_groupi_n_5563, csa_tree_add_51_79_groupi_n_5564, csa_tree_add_51_79_groupi_n_5565, csa_tree_add_51_79_groupi_n_5566, csa_tree_add_51_79_groupi_n_5567;
  wire csa_tree_add_51_79_groupi_n_5568, csa_tree_add_51_79_groupi_n_5569, csa_tree_add_51_79_groupi_n_5570, csa_tree_add_51_79_groupi_n_5571, csa_tree_add_51_79_groupi_n_5572, csa_tree_add_51_79_groupi_n_5573, csa_tree_add_51_79_groupi_n_5574, csa_tree_add_51_79_groupi_n_5575;
  wire csa_tree_add_51_79_groupi_n_5576, csa_tree_add_51_79_groupi_n_5577, csa_tree_add_51_79_groupi_n_5578, csa_tree_add_51_79_groupi_n_5579, csa_tree_add_51_79_groupi_n_5580, csa_tree_add_51_79_groupi_n_5581, csa_tree_add_51_79_groupi_n_5582, csa_tree_add_51_79_groupi_n_5583;
  wire csa_tree_add_51_79_groupi_n_5584, csa_tree_add_51_79_groupi_n_5585, csa_tree_add_51_79_groupi_n_5586, csa_tree_add_51_79_groupi_n_5587, csa_tree_add_51_79_groupi_n_5588, csa_tree_add_51_79_groupi_n_5589, csa_tree_add_51_79_groupi_n_5590, csa_tree_add_51_79_groupi_n_5591;
  wire csa_tree_add_51_79_groupi_n_5592, csa_tree_add_51_79_groupi_n_5593, csa_tree_add_51_79_groupi_n_5594, csa_tree_add_51_79_groupi_n_5595, csa_tree_add_51_79_groupi_n_5596, csa_tree_add_51_79_groupi_n_5597, csa_tree_add_51_79_groupi_n_5598, csa_tree_add_51_79_groupi_n_5599;
  wire csa_tree_add_51_79_groupi_n_5600, csa_tree_add_51_79_groupi_n_5601, csa_tree_add_51_79_groupi_n_5602, csa_tree_add_51_79_groupi_n_5603, csa_tree_add_51_79_groupi_n_5604, csa_tree_add_51_79_groupi_n_5605, csa_tree_add_51_79_groupi_n_5606, csa_tree_add_51_79_groupi_n_5607;
  wire csa_tree_add_51_79_groupi_n_5608, csa_tree_add_51_79_groupi_n_5609, csa_tree_add_51_79_groupi_n_5610, csa_tree_add_51_79_groupi_n_5611, csa_tree_add_51_79_groupi_n_5612, csa_tree_add_51_79_groupi_n_5613, csa_tree_add_51_79_groupi_n_5614, csa_tree_add_51_79_groupi_n_5615;
  wire csa_tree_add_51_79_groupi_n_5616, csa_tree_add_51_79_groupi_n_5617, csa_tree_add_51_79_groupi_n_5618, csa_tree_add_51_79_groupi_n_5619, csa_tree_add_51_79_groupi_n_5620, csa_tree_add_51_79_groupi_n_5621, csa_tree_add_51_79_groupi_n_5622, csa_tree_add_51_79_groupi_n_5623;
  wire csa_tree_add_51_79_groupi_n_5624, csa_tree_add_51_79_groupi_n_5625, csa_tree_add_51_79_groupi_n_5626, csa_tree_add_51_79_groupi_n_5627, csa_tree_add_51_79_groupi_n_5628, csa_tree_add_51_79_groupi_n_5629, csa_tree_add_51_79_groupi_n_5630, csa_tree_add_51_79_groupi_n_5631;
  wire csa_tree_add_51_79_groupi_n_5632, csa_tree_add_51_79_groupi_n_5633, csa_tree_add_51_79_groupi_n_5634, csa_tree_add_51_79_groupi_n_5635, csa_tree_add_51_79_groupi_n_5636, csa_tree_add_51_79_groupi_n_5637, csa_tree_add_51_79_groupi_n_5638, csa_tree_add_51_79_groupi_n_5639;
  wire csa_tree_add_51_79_groupi_n_5640, csa_tree_add_51_79_groupi_n_5641, csa_tree_add_51_79_groupi_n_5642, csa_tree_add_51_79_groupi_n_5643, csa_tree_add_51_79_groupi_n_5644, csa_tree_add_51_79_groupi_n_5645, csa_tree_add_51_79_groupi_n_5646, csa_tree_add_51_79_groupi_n_5647;
  wire csa_tree_add_51_79_groupi_n_5648, csa_tree_add_51_79_groupi_n_5649, csa_tree_add_51_79_groupi_n_5650, csa_tree_add_51_79_groupi_n_5651, csa_tree_add_51_79_groupi_n_5652, csa_tree_add_51_79_groupi_n_5653, csa_tree_add_51_79_groupi_n_5654, csa_tree_add_51_79_groupi_n_5655;
  wire csa_tree_add_51_79_groupi_n_5656, csa_tree_add_51_79_groupi_n_5657, csa_tree_add_51_79_groupi_n_5658, csa_tree_add_51_79_groupi_n_5659, csa_tree_add_51_79_groupi_n_5660, csa_tree_add_51_79_groupi_n_5661, csa_tree_add_51_79_groupi_n_5662, csa_tree_add_51_79_groupi_n_5663;
  wire csa_tree_add_51_79_groupi_n_5664, csa_tree_add_51_79_groupi_n_5665, csa_tree_add_51_79_groupi_n_5666, csa_tree_add_51_79_groupi_n_5667, csa_tree_add_51_79_groupi_n_5668, csa_tree_add_51_79_groupi_n_5669, csa_tree_add_51_79_groupi_n_5670, csa_tree_add_51_79_groupi_n_5671;
  wire csa_tree_add_51_79_groupi_n_5672, csa_tree_add_51_79_groupi_n_5673, csa_tree_add_51_79_groupi_n_5674, csa_tree_add_51_79_groupi_n_5675, csa_tree_add_51_79_groupi_n_5676, csa_tree_add_51_79_groupi_n_5677, csa_tree_add_51_79_groupi_n_5678, csa_tree_add_51_79_groupi_n_5679;
  wire csa_tree_add_51_79_groupi_n_5680, csa_tree_add_51_79_groupi_n_5681, csa_tree_add_51_79_groupi_n_5682, csa_tree_add_51_79_groupi_n_5683, csa_tree_add_51_79_groupi_n_5684, csa_tree_add_51_79_groupi_n_5685, csa_tree_add_51_79_groupi_n_5686, csa_tree_add_51_79_groupi_n_5687;
  wire csa_tree_add_51_79_groupi_n_5688, csa_tree_add_51_79_groupi_n_5689, csa_tree_add_51_79_groupi_n_5690, csa_tree_add_51_79_groupi_n_5691, csa_tree_add_51_79_groupi_n_5692, csa_tree_add_51_79_groupi_n_5693, csa_tree_add_51_79_groupi_n_5694, csa_tree_add_51_79_groupi_n_5695;
  wire csa_tree_add_51_79_groupi_n_5696, csa_tree_add_51_79_groupi_n_5697, csa_tree_add_51_79_groupi_n_5698, csa_tree_add_51_79_groupi_n_5699, csa_tree_add_51_79_groupi_n_5700, csa_tree_add_51_79_groupi_n_5701, csa_tree_add_51_79_groupi_n_5702, csa_tree_add_51_79_groupi_n_5703;
  wire csa_tree_add_51_79_groupi_n_5704, csa_tree_add_51_79_groupi_n_5705, csa_tree_add_51_79_groupi_n_5706, csa_tree_add_51_79_groupi_n_5707, csa_tree_add_51_79_groupi_n_5708, csa_tree_add_51_79_groupi_n_5709, csa_tree_add_51_79_groupi_n_5710, csa_tree_add_51_79_groupi_n_5711;
  wire csa_tree_add_51_79_groupi_n_5712, csa_tree_add_51_79_groupi_n_5713, csa_tree_add_51_79_groupi_n_5714, csa_tree_add_51_79_groupi_n_5715, csa_tree_add_51_79_groupi_n_5716, csa_tree_add_51_79_groupi_n_5717, csa_tree_add_51_79_groupi_n_5718, csa_tree_add_51_79_groupi_n_5719;
  wire csa_tree_add_51_79_groupi_n_5720, csa_tree_add_51_79_groupi_n_5721, csa_tree_add_51_79_groupi_n_5722, csa_tree_add_51_79_groupi_n_5723, csa_tree_add_51_79_groupi_n_5724, csa_tree_add_51_79_groupi_n_5725, csa_tree_add_51_79_groupi_n_5726, csa_tree_add_51_79_groupi_n_5727;
  wire csa_tree_add_51_79_groupi_n_5728, csa_tree_add_51_79_groupi_n_5729, csa_tree_add_51_79_groupi_n_5730, csa_tree_add_51_79_groupi_n_5731, csa_tree_add_51_79_groupi_n_5732, csa_tree_add_51_79_groupi_n_5733, csa_tree_add_51_79_groupi_n_5734, csa_tree_add_51_79_groupi_n_5735;
  wire csa_tree_add_51_79_groupi_n_5736, csa_tree_add_51_79_groupi_n_5737, csa_tree_add_51_79_groupi_n_5738, csa_tree_add_51_79_groupi_n_5739, csa_tree_add_51_79_groupi_n_5740, csa_tree_add_51_79_groupi_n_5741, csa_tree_add_51_79_groupi_n_5742, csa_tree_add_51_79_groupi_n_5743;
  wire csa_tree_add_51_79_groupi_n_5744, csa_tree_add_51_79_groupi_n_5745, csa_tree_add_51_79_groupi_n_5746, csa_tree_add_51_79_groupi_n_5747, csa_tree_add_51_79_groupi_n_5748, csa_tree_add_51_79_groupi_n_5749, csa_tree_add_51_79_groupi_n_5750, csa_tree_add_51_79_groupi_n_5751;
  wire csa_tree_add_51_79_groupi_n_5752, csa_tree_add_51_79_groupi_n_5753, csa_tree_add_51_79_groupi_n_5754, csa_tree_add_51_79_groupi_n_5755, csa_tree_add_51_79_groupi_n_5756, csa_tree_add_51_79_groupi_n_5757, csa_tree_add_51_79_groupi_n_5758, csa_tree_add_51_79_groupi_n_5759;
  wire csa_tree_add_51_79_groupi_n_5760, csa_tree_add_51_79_groupi_n_5761, csa_tree_add_51_79_groupi_n_5762, csa_tree_add_51_79_groupi_n_5763, csa_tree_add_51_79_groupi_n_5764, csa_tree_add_51_79_groupi_n_5765, csa_tree_add_51_79_groupi_n_5766, csa_tree_add_51_79_groupi_n_5767;
  wire csa_tree_add_51_79_groupi_n_5768, csa_tree_add_51_79_groupi_n_5769, csa_tree_add_51_79_groupi_n_5770, csa_tree_add_51_79_groupi_n_5771, csa_tree_add_51_79_groupi_n_5772, csa_tree_add_51_79_groupi_n_5773, csa_tree_add_51_79_groupi_n_5774, csa_tree_add_51_79_groupi_n_5775;
  wire csa_tree_add_51_79_groupi_n_5776, csa_tree_add_51_79_groupi_n_5777, csa_tree_add_51_79_groupi_n_5778, csa_tree_add_51_79_groupi_n_5779, csa_tree_add_51_79_groupi_n_5780, csa_tree_add_51_79_groupi_n_5781, csa_tree_add_51_79_groupi_n_5782, csa_tree_add_51_79_groupi_n_5783;
  wire csa_tree_add_51_79_groupi_n_5784, csa_tree_add_51_79_groupi_n_5785, csa_tree_add_51_79_groupi_n_5786, csa_tree_add_51_79_groupi_n_5787, csa_tree_add_51_79_groupi_n_5788, csa_tree_add_51_79_groupi_n_5789, csa_tree_add_51_79_groupi_n_5790, csa_tree_add_51_79_groupi_n_5791;
  wire csa_tree_add_51_79_groupi_n_5792, csa_tree_add_51_79_groupi_n_5793, csa_tree_add_51_79_groupi_n_5794, csa_tree_add_51_79_groupi_n_5795, csa_tree_add_51_79_groupi_n_5796, csa_tree_add_51_79_groupi_n_5797, csa_tree_add_51_79_groupi_n_5798, csa_tree_add_51_79_groupi_n_5799;
  wire csa_tree_add_51_79_groupi_n_5800, csa_tree_add_51_79_groupi_n_5801, csa_tree_add_51_79_groupi_n_5802, csa_tree_add_51_79_groupi_n_5803, csa_tree_add_51_79_groupi_n_5804, csa_tree_add_51_79_groupi_n_5805, csa_tree_add_51_79_groupi_n_5806, csa_tree_add_51_79_groupi_n_5807;
  wire csa_tree_add_51_79_groupi_n_5808, csa_tree_add_51_79_groupi_n_5809, csa_tree_add_51_79_groupi_n_5810, csa_tree_add_51_79_groupi_n_5811, csa_tree_add_51_79_groupi_n_5812, csa_tree_add_51_79_groupi_n_5813, csa_tree_add_51_79_groupi_n_5814, csa_tree_add_51_79_groupi_n_5815;
  wire csa_tree_add_51_79_groupi_n_5816, csa_tree_add_51_79_groupi_n_5817, csa_tree_add_51_79_groupi_n_5818, csa_tree_add_51_79_groupi_n_5819, csa_tree_add_51_79_groupi_n_5820, csa_tree_add_51_79_groupi_n_5821, csa_tree_add_51_79_groupi_n_5822, csa_tree_add_51_79_groupi_n_5823;
  wire csa_tree_add_51_79_groupi_n_5824, csa_tree_add_51_79_groupi_n_5825, csa_tree_add_51_79_groupi_n_5826, csa_tree_add_51_79_groupi_n_5827, csa_tree_add_51_79_groupi_n_5828, csa_tree_add_51_79_groupi_n_5829, csa_tree_add_51_79_groupi_n_5830, csa_tree_add_51_79_groupi_n_5831;
  wire csa_tree_add_51_79_groupi_n_5832, csa_tree_add_51_79_groupi_n_5833, csa_tree_add_51_79_groupi_n_5834, csa_tree_add_51_79_groupi_n_5835, csa_tree_add_51_79_groupi_n_5836, csa_tree_add_51_79_groupi_n_5837, csa_tree_add_51_79_groupi_n_5838, csa_tree_add_51_79_groupi_n_5839;
  wire csa_tree_add_51_79_groupi_n_5840, csa_tree_add_51_79_groupi_n_5841, csa_tree_add_51_79_groupi_n_5842, csa_tree_add_51_79_groupi_n_5843, csa_tree_add_51_79_groupi_n_5844, csa_tree_add_51_79_groupi_n_5845, csa_tree_add_51_79_groupi_n_5846, csa_tree_add_51_79_groupi_n_5847;
  wire csa_tree_add_51_79_groupi_n_5848, csa_tree_add_51_79_groupi_n_5849, csa_tree_add_51_79_groupi_n_5850, csa_tree_add_51_79_groupi_n_5851, csa_tree_add_51_79_groupi_n_5852, csa_tree_add_51_79_groupi_n_5853, csa_tree_add_51_79_groupi_n_5854, csa_tree_add_51_79_groupi_n_5855;
  wire csa_tree_add_51_79_groupi_n_5856, csa_tree_add_51_79_groupi_n_5857, csa_tree_add_51_79_groupi_n_5858, csa_tree_add_51_79_groupi_n_5859, csa_tree_add_51_79_groupi_n_5860, csa_tree_add_51_79_groupi_n_5861, csa_tree_add_51_79_groupi_n_5862, csa_tree_add_51_79_groupi_n_5863;
  wire csa_tree_add_51_79_groupi_n_5864, csa_tree_add_51_79_groupi_n_5865, csa_tree_add_51_79_groupi_n_5866, csa_tree_add_51_79_groupi_n_5867, csa_tree_add_51_79_groupi_n_5868, csa_tree_add_51_79_groupi_n_5869, csa_tree_add_51_79_groupi_n_5870, csa_tree_add_51_79_groupi_n_5871;
  wire csa_tree_add_51_79_groupi_n_5872, csa_tree_add_51_79_groupi_n_5873, csa_tree_add_51_79_groupi_n_5874, csa_tree_add_51_79_groupi_n_5875, csa_tree_add_51_79_groupi_n_5876, csa_tree_add_51_79_groupi_n_5877, csa_tree_add_51_79_groupi_n_5878, csa_tree_add_51_79_groupi_n_5879;
  wire csa_tree_add_51_79_groupi_n_5880, csa_tree_add_51_79_groupi_n_5881, csa_tree_add_51_79_groupi_n_5882, csa_tree_add_51_79_groupi_n_5883, csa_tree_add_51_79_groupi_n_5884, csa_tree_add_51_79_groupi_n_5885, csa_tree_add_51_79_groupi_n_5886, csa_tree_add_51_79_groupi_n_5887;
  wire csa_tree_add_51_79_groupi_n_5888, csa_tree_add_51_79_groupi_n_5889, csa_tree_add_51_79_groupi_n_5890, csa_tree_add_51_79_groupi_n_5891, csa_tree_add_51_79_groupi_n_5892, csa_tree_add_51_79_groupi_n_5893, csa_tree_add_51_79_groupi_n_5894, csa_tree_add_51_79_groupi_n_5895;
  wire csa_tree_add_51_79_groupi_n_5896, csa_tree_add_51_79_groupi_n_5897, csa_tree_add_51_79_groupi_n_5898, csa_tree_add_51_79_groupi_n_5899, csa_tree_add_51_79_groupi_n_5900, csa_tree_add_51_79_groupi_n_5901, csa_tree_add_51_79_groupi_n_5902, csa_tree_add_51_79_groupi_n_5903;
  wire csa_tree_add_51_79_groupi_n_5904, csa_tree_add_51_79_groupi_n_5905, csa_tree_add_51_79_groupi_n_5906, csa_tree_add_51_79_groupi_n_5907, csa_tree_add_51_79_groupi_n_5908, csa_tree_add_51_79_groupi_n_5909, csa_tree_add_51_79_groupi_n_5910, csa_tree_add_51_79_groupi_n_5911;
  wire csa_tree_add_51_79_groupi_n_5912, csa_tree_add_51_79_groupi_n_5913, csa_tree_add_51_79_groupi_n_5914, csa_tree_add_51_79_groupi_n_5915, csa_tree_add_51_79_groupi_n_5916, csa_tree_add_51_79_groupi_n_5917, csa_tree_add_51_79_groupi_n_5918, csa_tree_add_51_79_groupi_n_5919;
  wire csa_tree_add_51_79_groupi_n_5920, csa_tree_add_51_79_groupi_n_5921, csa_tree_add_51_79_groupi_n_5922, csa_tree_add_51_79_groupi_n_5923, csa_tree_add_51_79_groupi_n_5924, csa_tree_add_51_79_groupi_n_5925, csa_tree_add_51_79_groupi_n_5926, csa_tree_add_51_79_groupi_n_5927;
  wire csa_tree_add_51_79_groupi_n_5928, csa_tree_add_51_79_groupi_n_5929, csa_tree_add_51_79_groupi_n_5930, csa_tree_add_51_79_groupi_n_5931, csa_tree_add_51_79_groupi_n_5932, csa_tree_add_51_79_groupi_n_5933, csa_tree_add_51_79_groupi_n_5934, csa_tree_add_51_79_groupi_n_5935;
  wire csa_tree_add_51_79_groupi_n_5936, csa_tree_add_51_79_groupi_n_5937, csa_tree_add_51_79_groupi_n_5938, csa_tree_add_51_79_groupi_n_5939, csa_tree_add_51_79_groupi_n_5940, csa_tree_add_51_79_groupi_n_5941, csa_tree_add_51_79_groupi_n_5942, csa_tree_add_51_79_groupi_n_5943;
  wire csa_tree_add_51_79_groupi_n_5944, csa_tree_add_51_79_groupi_n_5945, csa_tree_add_51_79_groupi_n_5946, csa_tree_add_51_79_groupi_n_5947, csa_tree_add_51_79_groupi_n_5948, csa_tree_add_51_79_groupi_n_5949, csa_tree_add_51_79_groupi_n_5950, csa_tree_add_51_79_groupi_n_5951;
  wire csa_tree_add_51_79_groupi_n_5952, csa_tree_add_51_79_groupi_n_5953, csa_tree_add_51_79_groupi_n_5954, csa_tree_add_51_79_groupi_n_5955, csa_tree_add_51_79_groupi_n_5956, csa_tree_add_51_79_groupi_n_5957, csa_tree_add_51_79_groupi_n_5958, csa_tree_add_51_79_groupi_n_5959;
  wire csa_tree_add_51_79_groupi_n_5960, csa_tree_add_51_79_groupi_n_5961, csa_tree_add_51_79_groupi_n_5962, csa_tree_add_51_79_groupi_n_5963, csa_tree_add_51_79_groupi_n_5964, csa_tree_add_51_79_groupi_n_5965, csa_tree_add_51_79_groupi_n_5966, csa_tree_add_51_79_groupi_n_5967;
  wire csa_tree_add_51_79_groupi_n_5968, csa_tree_add_51_79_groupi_n_5969, csa_tree_add_51_79_groupi_n_5970, csa_tree_add_51_79_groupi_n_5971, csa_tree_add_51_79_groupi_n_5972, csa_tree_add_51_79_groupi_n_5973, csa_tree_add_51_79_groupi_n_5974, csa_tree_add_51_79_groupi_n_5975;
  wire csa_tree_add_51_79_groupi_n_5976, csa_tree_add_51_79_groupi_n_5977, csa_tree_add_51_79_groupi_n_5978, csa_tree_add_51_79_groupi_n_5979, csa_tree_add_51_79_groupi_n_5980, csa_tree_add_51_79_groupi_n_5981, csa_tree_add_51_79_groupi_n_5982, csa_tree_add_51_79_groupi_n_5983;
  wire csa_tree_add_51_79_groupi_n_5984, csa_tree_add_51_79_groupi_n_5985, csa_tree_add_51_79_groupi_n_5986, csa_tree_add_51_79_groupi_n_5987, csa_tree_add_51_79_groupi_n_5988, csa_tree_add_51_79_groupi_n_5989, csa_tree_add_51_79_groupi_n_5990, csa_tree_add_51_79_groupi_n_5991;
  wire csa_tree_add_51_79_groupi_n_5992, csa_tree_add_51_79_groupi_n_5993, csa_tree_add_51_79_groupi_n_5994, csa_tree_add_51_79_groupi_n_5995, csa_tree_add_51_79_groupi_n_5996, csa_tree_add_51_79_groupi_n_5997, csa_tree_add_51_79_groupi_n_5998, csa_tree_add_51_79_groupi_n_5999;
  wire csa_tree_add_51_79_groupi_n_6000, csa_tree_add_51_79_groupi_n_6001, csa_tree_add_51_79_groupi_n_6002, csa_tree_add_51_79_groupi_n_6003, csa_tree_add_51_79_groupi_n_6004, csa_tree_add_51_79_groupi_n_6005, csa_tree_add_51_79_groupi_n_6006, csa_tree_add_51_79_groupi_n_6007;
  wire csa_tree_add_51_79_groupi_n_6008, csa_tree_add_51_79_groupi_n_6009, csa_tree_add_51_79_groupi_n_6010, csa_tree_add_51_79_groupi_n_6011, csa_tree_add_51_79_groupi_n_6012, csa_tree_add_51_79_groupi_n_6013, csa_tree_add_51_79_groupi_n_6014, csa_tree_add_51_79_groupi_n_6015;
  wire csa_tree_add_51_79_groupi_n_6016, csa_tree_add_51_79_groupi_n_6017, csa_tree_add_51_79_groupi_n_6018, csa_tree_add_51_79_groupi_n_6019, csa_tree_add_51_79_groupi_n_6020, csa_tree_add_51_79_groupi_n_6021, csa_tree_add_51_79_groupi_n_6022, csa_tree_add_51_79_groupi_n_6023;
  wire csa_tree_add_51_79_groupi_n_6024, csa_tree_add_51_79_groupi_n_6025, csa_tree_add_51_79_groupi_n_6026, csa_tree_add_51_79_groupi_n_6027, csa_tree_add_51_79_groupi_n_6028, csa_tree_add_51_79_groupi_n_6029, csa_tree_add_51_79_groupi_n_6030, csa_tree_add_51_79_groupi_n_6031;
  wire csa_tree_add_51_79_groupi_n_6032, csa_tree_add_51_79_groupi_n_6033, csa_tree_add_51_79_groupi_n_6034, csa_tree_add_51_79_groupi_n_6035, csa_tree_add_51_79_groupi_n_6036, csa_tree_add_51_79_groupi_n_6037, csa_tree_add_51_79_groupi_n_6038, csa_tree_add_51_79_groupi_n_6039;
  wire csa_tree_add_51_79_groupi_n_6040, csa_tree_add_51_79_groupi_n_6041, csa_tree_add_51_79_groupi_n_6042, csa_tree_add_51_79_groupi_n_6043, csa_tree_add_51_79_groupi_n_6044, csa_tree_add_51_79_groupi_n_6045, csa_tree_add_51_79_groupi_n_6046, csa_tree_add_51_79_groupi_n_6047;
  wire csa_tree_add_51_79_groupi_n_6048, csa_tree_add_51_79_groupi_n_6049, csa_tree_add_51_79_groupi_n_6050, csa_tree_add_51_79_groupi_n_6051, csa_tree_add_51_79_groupi_n_6052, csa_tree_add_51_79_groupi_n_6053, csa_tree_add_51_79_groupi_n_6054, csa_tree_add_51_79_groupi_n_6055;
  wire csa_tree_add_51_79_groupi_n_6056, csa_tree_add_51_79_groupi_n_6057, csa_tree_add_51_79_groupi_n_6058, csa_tree_add_51_79_groupi_n_6059, csa_tree_add_51_79_groupi_n_6060, csa_tree_add_51_79_groupi_n_6061, csa_tree_add_51_79_groupi_n_6062, csa_tree_add_51_79_groupi_n_6063;
  wire csa_tree_add_51_79_groupi_n_6064, csa_tree_add_51_79_groupi_n_6065, csa_tree_add_51_79_groupi_n_6066, csa_tree_add_51_79_groupi_n_6067, csa_tree_add_51_79_groupi_n_6068, csa_tree_add_51_79_groupi_n_6069, csa_tree_add_51_79_groupi_n_6070, csa_tree_add_51_79_groupi_n_6071;
  wire csa_tree_add_51_79_groupi_n_6072, csa_tree_add_51_79_groupi_n_6073, csa_tree_add_51_79_groupi_n_6074, csa_tree_add_51_79_groupi_n_6075, csa_tree_add_51_79_groupi_n_6076, csa_tree_add_51_79_groupi_n_6077, csa_tree_add_51_79_groupi_n_6078, csa_tree_add_51_79_groupi_n_6079;
  wire csa_tree_add_51_79_groupi_n_6080, csa_tree_add_51_79_groupi_n_6081, csa_tree_add_51_79_groupi_n_6082, csa_tree_add_51_79_groupi_n_6083, csa_tree_add_51_79_groupi_n_6084, csa_tree_add_51_79_groupi_n_6085, csa_tree_add_51_79_groupi_n_6086, csa_tree_add_51_79_groupi_n_6087;
  wire csa_tree_add_51_79_groupi_n_6088, csa_tree_add_51_79_groupi_n_6089, csa_tree_add_51_79_groupi_n_6090, csa_tree_add_51_79_groupi_n_6091, csa_tree_add_51_79_groupi_n_6092, csa_tree_add_51_79_groupi_n_6093, csa_tree_add_51_79_groupi_n_6094, csa_tree_add_51_79_groupi_n_6095;
  wire csa_tree_add_51_79_groupi_n_6096, csa_tree_add_51_79_groupi_n_6097, csa_tree_add_51_79_groupi_n_6098, csa_tree_add_51_79_groupi_n_6099, csa_tree_add_51_79_groupi_n_6100, csa_tree_add_51_79_groupi_n_6101, csa_tree_add_51_79_groupi_n_6102, csa_tree_add_51_79_groupi_n_6103;
  wire csa_tree_add_51_79_groupi_n_6104, csa_tree_add_51_79_groupi_n_6105, csa_tree_add_51_79_groupi_n_6106, csa_tree_add_51_79_groupi_n_6107, csa_tree_add_51_79_groupi_n_6108, csa_tree_add_51_79_groupi_n_6109, csa_tree_add_51_79_groupi_n_6110, csa_tree_add_51_79_groupi_n_6111;
  wire csa_tree_add_51_79_groupi_n_6112, csa_tree_add_51_79_groupi_n_6113, csa_tree_add_51_79_groupi_n_6114, csa_tree_add_51_79_groupi_n_6115, csa_tree_add_51_79_groupi_n_6116, csa_tree_add_51_79_groupi_n_6117, csa_tree_add_51_79_groupi_n_6118, csa_tree_add_51_79_groupi_n_6119;
  wire csa_tree_add_51_79_groupi_n_6120, csa_tree_add_51_79_groupi_n_6121, csa_tree_add_51_79_groupi_n_6122, csa_tree_add_51_79_groupi_n_6123, csa_tree_add_51_79_groupi_n_6124, csa_tree_add_51_79_groupi_n_6125, csa_tree_add_51_79_groupi_n_6126, csa_tree_add_51_79_groupi_n_6127;
  wire csa_tree_add_51_79_groupi_n_6128, csa_tree_add_51_79_groupi_n_6129, csa_tree_add_51_79_groupi_n_6130, csa_tree_add_51_79_groupi_n_6131, csa_tree_add_51_79_groupi_n_6132, csa_tree_add_51_79_groupi_n_6133, csa_tree_add_51_79_groupi_n_6134, csa_tree_add_51_79_groupi_n_6135;
  wire csa_tree_add_51_79_groupi_n_6136, csa_tree_add_51_79_groupi_n_6137, csa_tree_add_51_79_groupi_n_6138, csa_tree_add_51_79_groupi_n_6139, csa_tree_add_51_79_groupi_n_6140, csa_tree_add_51_79_groupi_n_6141, csa_tree_add_51_79_groupi_n_6142, csa_tree_add_51_79_groupi_n_6143;
  wire csa_tree_add_51_79_groupi_n_6144, csa_tree_add_51_79_groupi_n_6145, csa_tree_add_51_79_groupi_n_6146, csa_tree_add_51_79_groupi_n_6147, csa_tree_add_51_79_groupi_n_6148, csa_tree_add_51_79_groupi_n_6149, csa_tree_add_51_79_groupi_n_6150, csa_tree_add_51_79_groupi_n_6151;
  wire csa_tree_add_51_79_groupi_n_6152, csa_tree_add_51_79_groupi_n_6153, csa_tree_add_51_79_groupi_n_6154, csa_tree_add_51_79_groupi_n_6155, csa_tree_add_51_79_groupi_n_6156, csa_tree_add_51_79_groupi_n_6157, csa_tree_add_51_79_groupi_n_6158, csa_tree_add_51_79_groupi_n_6159;
  wire csa_tree_add_51_79_groupi_n_6160, csa_tree_add_51_79_groupi_n_6161, csa_tree_add_51_79_groupi_n_6162, csa_tree_add_51_79_groupi_n_6163, csa_tree_add_51_79_groupi_n_6164, csa_tree_add_51_79_groupi_n_6165, csa_tree_add_51_79_groupi_n_6166, csa_tree_add_51_79_groupi_n_6167;
  wire csa_tree_add_51_79_groupi_n_6168, csa_tree_add_51_79_groupi_n_6169, csa_tree_add_51_79_groupi_n_6170, csa_tree_add_51_79_groupi_n_6171, csa_tree_add_51_79_groupi_n_6172, csa_tree_add_51_79_groupi_n_6173, csa_tree_add_51_79_groupi_n_6174, csa_tree_add_51_79_groupi_n_6175;
  wire csa_tree_add_51_79_groupi_n_6176, csa_tree_add_51_79_groupi_n_6177, csa_tree_add_51_79_groupi_n_6178, csa_tree_add_51_79_groupi_n_6179, csa_tree_add_51_79_groupi_n_6180, csa_tree_add_51_79_groupi_n_6181, csa_tree_add_51_79_groupi_n_6182, csa_tree_add_51_79_groupi_n_6183;
  wire csa_tree_add_51_79_groupi_n_6184, csa_tree_add_51_79_groupi_n_6185, csa_tree_add_51_79_groupi_n_6186, csa_tree_add_51_79_groupi_n_6187, csa_tree_add_51_79_groupi_n_6188, csa_tree_add_51_79_groupi_n_6189, csa_tree_add_51_79_groupi_n_6190, csa_tree_add_51_79_groupi_n_6191;
  wire csa_tree_add_51_79_groupi_n_6192, csa_tree_add_51_79_groupi_n_6193, csa_tree_add_51_79_groupi_n_6194, csa_tree_add_51_79_groupi_n_6195, csa_tree_add_51_79_groupi_n_6196, csa_tree_add_51_79_groupi_n_6197, csa_tree_add_51_79_groupi_n_6198, csa_tree_add_51_79_groupi_n_6199;
  wire csa_tree_add_51_79_groupi_n_6200, csa_tree_add_51_79_groupi_n_6201, csa_tree_add_51_79_groupi_n_6202, csa_tree_add_51_79_groupi_n_6203, csa_tree_add_51_79_groupi_n_6204, csa_tree_add_51_79_groupi_n_6205, csa_tree_add_51_79_groupi_n_6206, csa_tree_add_51_79_groupi_n_6207;
  wire csa_tree_add_51_79_groupi_n_6208, csa_tree_add_51_79_groupi_n_6209, csa_tree_add_51_79_groupi_n_6210, csa_tree_add_51_79_groupi_n_6211, csa_tree_add_51_79_groupi_n_6212, csa_tree_add_51_79_groupi_n_6213, csa_tree_add_51_79_groupi_n_6214, csa_tree_add_51_79_groupi_n_6215;
  wire csa_tree_add_51_79_groupi_n_6216, csa_tree_add_51_79_groupi_n_6217, csa_tree_add_51_79_groupi_n_6218, csa_tree_add_51_79_groupi_n_6219, csa_tree_add_51_79_groupi_n_6220, csa_tree_add_51_79_groupi_n_6221, csa_tree_add_51_79_groupi_n_6222, csa_tree_add_51_79_groupi_n_6223;
  wire csa_tree_add_51_79_groupi_n_6224, csa_tree_add_51_79_groupi_n_6225, csa_tree_add_51_79_groupi_n_6226, csa_tree_add_51_79_groupi_n_6227, csa_tree_add_51_79_groupi_n_6228, csa_tree_add_51_79_groupi_n_6229, csa_tree_add_51_79_groupi_n_6230, csa_tree_add_51_79_groupi_n_6231;
  wire csa_tree_add_51_79_groupi_n_6232, csa_tree_add_51_79_groupi_n_6233, csa_tree_add_51_79_groupi_n_6234, csa_tree_add_51_79_groupi_n_6235, csa_tree_add_51_79_groupi_n_6236, csa_tree_add_51_79_groupi_n_6237, csa_tree_add_51_79_groupi_n_6238, csa_tree_add_51_79_groupi_n_6239;
  wire csa_tree_add_51_79_groupi_n_6240, csa_tree_add_51_79_groupi_n_6241, csa_tree_add_51_79_groupi_n_6242, csa_tree_add_51_79_groupi_n_6243, csa_tree_add_51_79_groupi_n_6244, csa_tree_add_51_79_groupi_n_6245, csa_tree_add_51_79_groupi_n_6246, csa_tree_add_51_79_groupi_n_6247;
  wire csa_tree_add_51_79_groupi_n_6248, csa_tree_add_51_79_groupi_n_6249, csa_tree_add_51_79_groupi_n_6250, csa_tree_add_51_79_groupi_n_6251, csa_tree_add_51_79_groupi_n_6252, csa_tree_add_51_79_groupi_n_6253, csa_tree_add_51_79_groupi_n_6254, csa_tree_add_51_79_groupi_n_6255;
  wire csa_tree_add_51_79_groupi_n_6256, csa_tree_add_51_79_groupi_n_6257, csa_tree_add_51_79_groupi_n_6258, csa_tree_add_51_79_groupi_n_6259, csa_tree_add_51_79_groupi_n_6260, csa_tree_add_51_79_groupi_n_6261, csa_tree_add_51_79_groupi_n_6262, csa_tree_add_51_79_groupi_n_6263;
  wire csa_tree_add_51_79_groupi_n_6264, csa_tree_add_51_79_groupi_n_6265, csa_tree_add_51_79_groupi_n_6266, csa_tree_add_51_79_groupi_n_6267, csa_tree_add_51_79_groupi_n_6268, csa_tree_add_51_79_groupi_n_6269, csa_tree_add_51_79_groupi_n_6270, csa_tree_add_51_79_groupi_n_6271;
  wire csa_tree_add_51_79_groupi_n_6272, csa_tree_add_51_79_groupi_n_6273, csa_tree_add_51_79_groupi_n_6274, csa_tree_add_51_79_groupi_n_6275, csa_tree_add_51_79_groupi_n_6276, csa_tree_add_51_79_groupi_n_6277, csa_tree_add_51_79_groupi_n_6278, csa_tree_add_51_79_groupi_n_6279;
  wire csa_tree_add_51_79_groupi_n_6280, csa_tree_add_51_79_groupi_n_6281, csa_tree_add_51_79_groupi_n_6282, csa_tree_add_51_79_groupi_n_6283, csa_tree_add_51_79_groupi_n_6284, csa_tree_add_51_79_groupi_n_6285, csa_tree_add_51_79_groupi_n_6286, csa_tree_add_51_79_groupi_n_6287;
  wire csa_tree_add_51_79_groupi_n_6288, csa_tree_add_51_79_groupi_n_6289, csa_tree_add_51_79_groupi_n_6290, csa_tree_add_51_79_groupi_n_6291, csa_tree_add_51_79_groupi_n_6292, csa_tree_add_51_79_groupi_n_6293, csa_tree_add_51_79_groupi_n_6294, csa_tree_add_51_79_groupi_n_6295;
  wire csa_tree_add_51_79_groupi_n_6296, csa_tree_add_51_79_groupi_n_6297, csa_tree_add_51_79_groupi_n_6298, csa_tree_add_51_79_groupi_n_6299, csa_tree_add_51_79_groupi_n_6300, csa_tree_add_51_79_groupi_n_6301, csa_tree_add_51_79_groupi_n_6302, csa_tree_add_51_79_groupi_n_6303;
  wire csa_tree_add_51_79_groupi_n_6304, csa_tree_add_51_79_groupi_n_6305, csa_tree_add_51_79_groupi_n_6306, csa_tree_add_51_79_groupi_n_6307, csa_tree_add_51_79_groupi_n_6308, csa_tree_add_51_79_groupi_n_6309, csa_tree_add_51_79_groupi_n_6310, csa_tree_add_51_79_groupi_n_6311;
  wire csa_tree_add_51_79_groupi_n_6312, csa_tree_add_51_79_groupi_n_6313, csa_tree_add_51_79_groupi_n_6314, csa_tree_add_51_79_groupi_n_6315, csa_tree_add_51_79_groupi_n_6316, csa_tree_add_51_79_groupi_n_6317, csa_tree_add_51_79_groupi_n_6318, csa_tree_add_51_79_groupi_n_6319;
  wire csa_tree_add_51_79_groupi_n_6320, csa_tree_add_51_79_groupi_n_6321, csa_tree_add_51_79_groupi_n_6322, csa_tree_add_51_79_groupi_n_6323, csa_tree_add_51_79_groupi_n_6324, csa_tree_add_51_79_groupi_n_6325, csa_tree_add_51_79_groupi_n_6326, csa_tree_add_51_79_groupi_n_6327;
  wire csa_tree_add_51_79_groupi_n_6328, csa_tree_add_51_79_groupi_n_6329, csa_tree_add_51_79_groupi_n_6330, csa_tree_add_51_79_groupi_n_6331, csa_tree_add_51_79_groupi_n_6332, csa_tree_add_51_79_groupi_n_6333, csa_tree_add_51_79_groupi_n_6334, csa_tree_add_51_79_groupi_n_6335;
  wire csa_tree_add_51_79_groupi_n_6336, csa_tree_add_51_79_groupi_n_6337, csa_tree_add_51_79_groupi_n_6338, csa_tree_add_51_79_groupi_n_6339, csa_tree_add_51_79_groupi_n_6340, csa_tree_add_51_79_groupi_n_6341, csa_tree_add_51_79_groupi_n_6342, csa_tree_add_51_79_groupi_n_6343;
  wire csa_tree_add_51_79_groupi_n_6344, csa_tree_add_51_79_groupi_n_6345, csa_tree_add_51_79_groupi_n_6346, csa_tree_add_51_79_groupi_n_6347, csa_tree_add_51_79_groupi_n_6348, csa_tree_add_51_79_groupi_n_6349, csa_tree_add_51_79_groupi_n_6350, csa_tree_add_51_79_groupi_n_6351;
  wire csa_tree_add_51_79_groupi_n_6352, csa_tree_add_51_79_groupi_n_6353, csa_tree_add_51_79_groupi_n_6354, csa_tree_add_51_79_groupi_n_6355, csa_tree_add_51_79_groupi_n_6356, csa_tree_add_51_79_groupi_n_6357, csa_tree_add_51_79_groupi_n_6358, csa_tree_add_51_79_groupi_n_6359;
  wire csa_tree_add_51_79_groupi_n_6360, csa_tree_add_51_79_groupi_n_6361, csa_tree_add_51_79_groupi_n_6362, csa_tree_add_51_79_groupi_n_6363, csa_tree_add_51_79_groupi_n_6364, csa_tree_add_51_79_groupi_n_6365, csa_tree_add_51_79_groupi_n_6366, csa_tree_add_51_79_groupi_n_6367;
  wire csa_tree_add_51_79_groupi_n_6368, csa_tree_add_51_79_groupi_n_6369, csa_tree_add_51_79_groupi_n_6370, csa_tree_add_51_79_groupi_n_6371, csa_tree_add_51_79_groupi_n_6372, csa_tree_add_51_79_groupi_n_6373, csa_tree_add_51_79_groupi_n_6374, csa_tree_add_51_79_groupi_n_6375;
  wire csa_tree_add_51_79_groupi_n_6376, csa_tree_add_51_79_groupi_n_6377, csa_tree_add_51_79_groupi_n_6378, csa_tree_add_51_79_groupi_n_6379, csa_tree_add_51_79_groupi_n_6380, csa_tree_add_51_79_groupi_n_6381, csa_tree_add_51_79_groupi_n_6382, csa_tree_add_51_79_groupi_n_6383;
  wire csa_tree_add_51_79_groupi_n_6384, csa_tree_add_51_79_groupi_n_6385, csa_tree_add_51_79_groupi_n_6386, csa_tree_add_51_79_groupi_n_6387, csa_tree_add_51_79_groupi_n_6388, csa_tree_add_51_79_groupi_n_6389, csa_tree_add_51_79_groupi_n_6390, csa_tree_add_51_79_groupi_n_6391;
  wire csa_tree_add_51_79_groupi_n_6392, csa_tree_add_51_79_groupi_n_6393, csa_tree_add_51_79_groupi_n_6394, csa_tree_add_51_79_groupi_n_6395, csa_tree_add_51_79_groupi_n_6396, csa_tree_add_51_79_groupi_n_6397, csa_tree_add_51_79_groupi_n_6398, csa_tree_add_51_79_groupi_n_6399;
  wire csa_tree_add_51_79_groupi_n_6400, csa_tree_add_51_79_groupi_n_6401, csa_tree_add_51_79_groupi_n_6402, csa_tree_add_51_79_groupi_n_6403, csa_tree_add_51_79_groupi_n_6404, csa_tree_add_51_79_groupi_n_6405, csa_tree_add_51_79_groupi_n_6406, csa_tree_add_51_79_groupi_n_6407;
  wire csa_tree_add_51_79_groupi_n_6408, csa_tree_add_51_79_groupi_n_6409, csa_tree_add_51_79_groupi_n_6410, csa_tree_add_51_79_groupi_n_6411, csa_tree_add_51_79_groupi_n_6412, csa_tree_add_51_79_groupi_n_6413, csa_tree_add_51_79_groupi_n_6414, csa_tree_add_51_79_groupi_n_6415;
  wire csa_tree_add_51_79_groupi_n_6416, csa_tree_add_51_79_groupi_n_6417, csa_tree_add_51_79_groupi_n_6418, csa_tree_add_51_79_groupi_n_6419, csa_tree_add_51_79_groupi_n_6420, csa_tree_add_51_79_groupi_n_6421, csa_tree_add_51_79_groupi_n_6422, csa_tree_add_51_79_groupi_n_6423;
  wire csa_tree_add_51_79_groupi_n_6424, csa_tree_add_51_79_groupi_n_6425, csa_tree_add_51_79_groupi_n_6426, csa_tree_add_51_79_groupi_n_6427, csa_tree_add_51_79_groupi_n_6428, csa_tree_add_51_79_groupi_n_6429, csa_tree_add_51_79_groupi_n_6430, csa_tree_add_51_79_groupi_n_6431;
  wire csa_tree_add_51_79_groupi_n_6432, csa_tree_add_51_79_groupi_n_6433, csa_tree_add_51_79_groupi_n_6434, csa_tree_add_51_79_groupi_n_6435, csa_tree_add_51_79_groupi_n_6436, csa_tree_add_51_79_groupi_n_6437, csa_tree_add_51_79_groupi_n_6438, csa_tree_add_51_79_groupi_n_6439;
  wire csa_tree_add_51_79_groupi_n_6440, csa_tree_add_51_79_groupi_n_6441, csa_tree_add_51_79_groupi_n_6442, csa_tree_add_51_79_groupi_n_6443, csa_tree_add_51_79_groupi_n_6444, csa_tree_add_51_79_groupi_n_6445, csa_tree_add_51_79_groupi_n_6446, csa_tree_add_51_79_groupi_n_6447;
  wire csa_tree_add_51_79_groupi_n_6448, csa_tree_add_51_79_groupi_n_6449, csa_tree_add_51_79_groupi_n_6450, csa_tree_add_51_79_groupi_n_6451, csa_tree_add_51_79_groupi_n_6452, csa_tree_add_51_79_groupi_n_6453, csa_tree_add_51_79_groupi_n_6454, csa_tree_add_51_79_groupi_n_6455;
  wire csa_tree_add_51_79_groupi_n_6456, csa_tree_add_51_79_groupi_n_6457, csa_tree_add_51_79_groupi_n_6458, csa_tree_add_51_79_groupi_n_6459, csa_tree_add_51_79_groupi_n_6460, csa_tree_add_51_79_groupi_n_6461, csa_tree_add_51_79_groupi_n_6462, csa_tree_add_51_79_groupi_n_6463;
  wire csa_tree_add_51_79_groupi_n_6464, csa_tree_add_51_79_groupi_n_6465, csa_tree_add_51_79_groupi_n_6466, csa_tree_add_51_79_groupi_n_6467, csa_tree_add_51_79_groupi_n_6468, csa_tree_add_51_79_groupi_n_6469, csa_tree_add_51_79_groupi_n_6470, csa_tree_add_51_79_groupi_n_6471;
  wire csa_tree_add_51_79_groupi_n_6472, csa_tree_add_51_79_groupi_n_6473, csa_tree_add_51_79_groupi_n_6474, csa_tree_add_51_79_groupi_n_6475, csa_tree_add_51_79_groupi_n_6476, csa_tree_add_51_79_groupi_n_6477, csa_tree_add_51_79_groupi_n_6478, csa_tree_add_51_79_groupi_n_6479;
  wire csa_tree_add_51_79_groupi_n_6480, csa_tree_add_51_79_groupi_n_6481, csa_tree_add_51_79_groupi_n_6482, csa_tree_add_51_79_groupi_n_6483, csa_tree_add_51_79_groupi_n_6484, csa_tree_add_51_79_groupi_n_6485, csa_tree_add_51_79_groupi_n_6486, csa_tree_add_51_79_groupi_n_6487;
  wire csa_tree_add_51_79_groupi_n_6488, csa_tree_add_51_79_groupi_n_6489, csa_tree_add_51_79_groupi_n_6490, csa_tree_add_51_79_groupi_n_6491, csa_tree_add_51_79_groupi_n_6492, csa_tree_add_51_79_groupi_n_6493, csa_tree_add_51_79_groupi_n_6494, csa_tree_add_51_79_groupi_n_6495;
  wire csa_tree_add_51_79_groupi_n_6496, csa_tree_add_51_79_groupi_n_6497, csa_tree_add_51_79_groupi_n_6498, csa_tree_add_51_79_groupi_n_6499, csa_tree_add_51_79_groupi_n_6500, csa_tree_add_51_79_groupi_n_6501, csa_tree_add_51_79_groupi_n_6502, csa_tree_add_51_79_groupi_n_6503;
  wire csa_tree_add_51_79_groupi_n_6504, csa_tree_add_51_79_groupi_n_6505, csa_tree_add_51_79_groupi_n_6506, csa_tree_add_51_79_groupi_n_6507, csa_tree_add_51_79_groupi_n_6508, csa_tree_add_51_79_groupi_n_6509, csa_tree_add_51_79_groupi_n_6510, csa_tree_add_51_79_groupi_n_6511;
  wire csa_tree_add_51_79_groupi_n_6512, csa_tree_add_51_79_groupi_n_6513, csa_tree_add_51_79_groupi_n_6514, csa_tree_add_51_79_groupi_n_6515, csa_tree_add_51_79_groupi_n_6516, csa_tree_add_51_79_groupi_n_6517, csa_tree_add_51_79_groupi_n_6518, csa_tree_add_51_79_groupi_n_6519;
  wire csa_tree_add_51_79_groupi_n_6520, csa_tree_add_51_79_groupi_n_6521, csa_tree_add_51_79_groupi_n_6522, csa_tree_add_51_79_groupi_n_6523, csa_tree_add_51_79_groupi_n_6524, csa_tree_add_51_79_groupi_n_6525, csa_tree_add_51_79_groupi_n_6526, csa_tree_add_51_79_groupi_n_6527;
  wire csa_tree_add_51_79_groupi_n_6528, csa_tree_add_51_79_groupi_n_6529, csa_tree_add_51_79_groupi_n_6530, csa_tree_add_51_79_groupi_n_6531, csa_tree_add_51_79_groupi_n_6532, csa_tree_add_51_79_groupi_n_6533, csa_tree_add_51_79_groupi_n_6534, csa_tree_add_51_79_groupi_n_6535;
  wire csa_tree_add_51_79_groupi_n_6536, csa_tree_add_51_79_groupi_n_6537, csa_tree_add_51_79_groupi_n_6538, csa_tree_add_51_79_groupi_n_6539, csa_tree_add_51_79_groupi_n_6540, csa_tree_add_51_79_groupi_n_6541, csa_tree_add_51_79_groupi_n_6542, csa_tree_add_51_79_groupi_n_6543;
  wire csa_tree_add_51_79_groupi_n_6544, csa_tree_add_51_79_groupi_n_6545, csa_tree_add_51_79_groupi_n_6546, csa_tree_add_51_79_groupi_n_6547, csa_tree_add_51_79_groupi_n_6548, csa_tree_add_51_79_groupi_n_6549, csa_tree_add_51_79_groupi_n_6550, csa_tree_add_51_79_groupi_n_6551;
  wire csa_tree_add_51_79_groupi_n_6552, csa_tree_add_51_79_groupi_n_6553, csa_tree_add_51_79_groupi_n_6554, csa_tree_add_51_79_groupi_n_6555, csa_tree_add_51_79_groupi_n_6556, csa_tree_add_51_79_groupi_n_6557, csa_tree_add_51_79_groupi_n_6558, csa_tree_add_51_79_groupi_n_6559;
  wire csa_tree_add_51_79_groupi_n_6560, csa_tree_add_51_79_groupi_n_6561, csa_tree_add_51_79_groupi_n_6562, csa_tree_add_51_79_groupi_n_6563, csa_tree_add_51_79_groupi_n_6564, csa_tree_add_51_79_groupi_n_6565, csa_tree_add_51_79_groupi_n_6566, csa_tree_add_51_79_groupi_n_6567;
  wire csa_tree_add_51_79_groupi_n_6568, csa_tree_add_51_79_groupi_n_6569, csa_tree_add_51_79_groupi_n_6570, csa_tree_add_51_79_groupi_n_6571, csa_tree_add_51_79_groupi_n_6572, csa_tree_add_51_79_groupi_n_6573, csa_tree_add_51_79_groupi_n_6574, csa_tree_add_51_79_groupi_n_6575;
  wire csa_tree_add_51_79_groupi_n_6576, csa_tree_add_51_79_groupi_n_6577, csa_tree_add_51_79_groupi_n_6578, csa_tree_add_51_79_groupi_n_6579, csa_tree_add_51_79_groupi_n_6580, csa_tree_add_51_79_groupi_n_6581, csa_tree_add_51_79_groupi_n_6582, csa_tree_add_51_79_groupi_n_6583;
  wire csa_tree_add_51_79_groupi_n_6584, csa_tree_add_51_79_groupi_n_6585, csa_tree_add_51_79_groupi_n_6586, csa_tree_add_51_79_groupi_n_6587, csa_tree_add_51_79_groupi_n_6588, csa_tree_add_51_79_groupi_n_6589, csa_tree_add_51_79_groupi_n_6590, csa_tree_add_51_79_groupi_n_6591;
  wire csa_tree_add_51_79_groupi_n_6592, csa_tree_add_51_79_groupi_n_6593, csa_tree_add_51_79_groupi_n_6594, csa_tree_add_51_79_groupi_n_6595, csa_tree_add_51_79_groupi_n_6596, csa_tree_add_51_79_groupi_n_6597, csa_tree_add_51_79_groupi_n_6598, csa_tree_add_51_79_groupi_n_6599;
  wire csa_tree_add_51_79_groupi_n_6600, csa_tree_add_51_79_groupi_n_6601, csa_tree_add_51_79_groupi_n_6602, csa_tree_add_51_79_groupi_n_6603, csa_tree_add_51_79_groupi_n_6604, csa_tree_add_51_79_groupi_n_6605, csa_tree_add_51_79_groupi_n_6606, csa_tree_add_51_79_groupi_n_6607;
  wire csa_tree_add_51_79_groupi_n_6608, csa_tree_add_51_79_groupi_n_6609, csa_tree_add_51_79_groupi_n_6610, csa_tree_add_51_79_groupi_n_6611, csa_tree_add_51_79_groupi_n_6612, csa_tree_add_51_79_groupi_n_6613, csa_tree_add_51_79_groupi_n_6614, csa_tree_add_51_79_groupi_n_6615;
  wire csa_tree_add_51_79_groupi_n_6616, csa_tree_add_51_79_groupi_n_6617, csa_tree_add_51_79_groupi_n_6618, csa_tree_add_51_79_groupi_n_6619, csa_tree_add_51_79_groupi_n_6620, csa_tree_add_51_79_groupi_n_6621, csa_tree_add_51_79_groupi_n_6622, csa_tree_add_51_79_groupi_n_6623;
  wire csa_tree_add_51_79_groupi_n_6624, csa_tree_add_51_79_groupi_n_6625, csa_tree_add_51_79_groupi_n_6626, csa_tree_add_51_79_groupi_n_6627, csa_tree_add_51_79_groupi_n_6628, csa_tree_add_51_79_groupi_n_6629, csa_tree_add_51_79_groupi_n_6630, csa_tree_add_51_79_groupi_n_6631;
  wire csa_tree_add_51_79_groupi_n_6632, csa_tree_add_51_79_groupi_n_6633, csa_tree_add_51_79_groupi_n_6634, csa_tree_add_51_79_groupi_n_6635, csa_tree_add_51_79_groupi_n_6636, csa_tree_add_51_79_groupi_n_6637, csa_tree_add_51_79_groupi_n_6638, csa_tree_add_51_79_groupi_n_6639;
  wire csa_tree_add_51_79_groupi_n_6640, csa_tree_add_51_79_groupi_n_6641, csa_tree_add_51_79_groupi_n_6642, csa_tree_add_51_79_groupi_n_6643, csa_tree_add_51_79_groupi_n_6644, csa_tree_add_51_79_groupi_n_6645, csa_tree_add_51_79_groupi_n_6646, csa_tree_add_51_79_groupi_n_6647;
  wire csa_tree_add_51_79_groupi_n_6648, csa_tree_add_51_79_groupi_n_6649, csa_tree_add_51_79_groupi_n_6650, csa_tree_add_51_79_groupi_n_6651, csa_tree_add_51_79_groupi_n_6652, csa_tree_add_51_79_groupi_n_6653, csa_tree_add_51_79_groupi_n_6654, csa_tree_add_51_79_groupi_n_6655;
  wire csa_tree_add_51_79_groupi_n_6656, csa_tree_add_51_79_groupi_n_6657, csa_tree_add_51_79_groupi_n_6658, csa_tree_add_51_79_groupi_n_6659, csa_tree_add_51_79_groupi_n_6660, csa_tree_add_51_79_groupi_n_6661, csa_tree_add_51_79_groupi_n_6662, csa_tree_add_51_79_groupi_n_6663;
  wire csa_tree_add_51_79_groupi_n_6664, csa_tree_add_51_79_groupi_n_6665, csa_tree_add_51_79_groupi_n_6666, csa_tree_add_51_79_groupi_n_6667, csa_tree_add_51_79_groupi_n_6668, csa_tree_add_51_79_groupi_n_6669, csa_tree_add_51_79_groupi_n_6670, csa_tree_add_51_79_groupi_n_6671;
  wire csa_tree_add_51_79_groupi_n_6672, csa_tree_add_51_79_groupi_n_6673, csa_tree_add_51_79_groupi_n_6674, csa_tree_add_51_79_groupi_n_6675, csa_tree_add_51_79_groupi_n_6676, csa_tree_add_51_79_groupi_n_6677, csa_tree_add_51_79_groupi_n_6678, csa_tree_add_51_79_groupi_n_6679;
  wire csa_tree_add_51_79_groupi_n_6680, csa_tree_add_51_79_groupi_n_6681, csa_tree_add_51_79_groupi_n_6682, csa_tree_add_51_79_groupi_n_6683, csa_tree_add_51_79_groupi_n_6684, csa_tree_add_51_79_groupi_n_6685, csa_tree_add_51_79_groupi_n_6686, csa_tree_add_51_79_groupi_n_6687;
  wire csa_tree_add_51_79_groupi_n_6688, csa_tree_add_51_79_groupi_n_6689, csa_tree_add_51_79_groupi_n_6690, csa_tree_add_51_79_groupi_n_6691, csa_tree_add_51_79_groupi_n_6692, csa_tree_add_51_79_groupi_n_6693, csa_tree_add_51_79_groupi_n_6694, csa_tree_add_51_79_groupi_n_6695;
  wire csa_tree_add_51_79_groupi_n_6696, csa_tree_add_51_79_groupi_n_6697, csa_tree_add_51_79_groupi_n_6698, csa_tree_add_51_79_groupi_n_6699, csa_tree_add_51_79_groupi_n_6700, csa_tree_add_51_79_groupi_n_6701, csa_tree_add_51_79_groupi_n_6702, csa_tree_add_51_79_groupi_n_6703;
  wire csa_tree_add_51_79_groupi_n_6704, csa_tree_add_51_79_groupi_n_6705, csa_tree_add_51_79_groupi_n_6706, csa_tree_add_51_79_groupi_n_6707, csa_tree_add_51_79_groupi_n_6708, csa_tree_add_51_79_groupi_n_6709, csa_tree_add_51_79_groupi_n_6710, csa_tree_add_51_79_groupi_n_6711;
  wire csa_tree_add_51_79_groupi_n_6712, csa_tree_add_51_79_groupi_n_6713, csa_tree_add_51_79_groupi_n_6714, csa_tree_add_51_79_groupi_n_6715, csa_tree_add_51_79_groupi_n_6716, csa_tree_add_51_79_groupi_n_6717, csa_tree_add_51_79_groupi_n_6718, csa_tree_add_51_79_groupi_n_6719;
  wire csa_tree_add_51_79_groupi_n_6720, csa_tree_add_51_79_groupi_n_6721, csa_tree_add_51_79_groupi_n_6722, csa_tree_add_51_79_groupi_n_6723, csa_tree_add_51_79_groupi_n_6724, csa_tree_add_51_79_groupi_n_6725, csa_tree_add_51_79_groupi_n_6726, csa_tree_add_51_79_groupi_n_6727;
  wire csa_tree_add_51_79_groupi_n_6728, csa_tree_add_51_79_groupi_n_6729, csa_tree_add_51_79_groupi_n_6730, csa_tree_add_51_79_groupi_n_6731, csa_tree_add_51_79_groupi_n_6732, csa_tree_add_51_79_groupi_n_6733, csa_tree_add_51_79_groupi_n_6734, csa_tree_add_51_79_groupi_n_6735;
  wire csa_tree_add_51_79_groupi_n_6736, csa_tree_add_51_79_groupi_n_6737, csa_tree_add_51_79_groupi_n_6738, csa_tree_add_51_79_groupi_n_6739, csa_tree_add_51_79_groupi_n_6740, csa_tree_add_51_79_groupi_n_6741, csa_tree_add_51_79_groupi_n_6742, csa_tree_add_51_79_groupi_n_6743;
  wire csa_tree_add_51_79_groupi_n_6744, csa_tree_add_51_79_groupi_n_6745, csa_tree_add_51_79_groupi_n_6746, csa_tree_add_51_79_groupi_n_6747, csa_tree_add_51_79_groupi_n_6748, csa_tree_add_51_79_groupi_n_6749, csa_tree_add_51_79_groupi_n_6750, csa_tree_add_51_79_groupi_n_6751;
  wire csa_tree_add_51_79_groupi_n_6752, csa_tree_add_51_79_groupi_n_6753, csa_tree_add_51_79_groupi_n_6754, csa_tree_add_51_79_groupi_n_6755, csa_tree_add_51_79_groupi_n_6756, csa_tree_add_51_79_groupi_n_6757, csa_tree_add_51_79_groupi_n_6758, csa_tree_add_51_79_groupi_n_6759;
  wire csa_tree_add_51_79_groupi_n_6760, csa_tree_add_51_79_groupi_n_6761, csa_tree_add_51_79_groupi_n_6762, csa_tree_add_51_79_groupi_n_6763, csa_tree_add_51_79_groupi_n_6764, csa_tree_add_51_79_groupi_n_6765, csa_tree_add_51_79_groupi_n_6766, csa_tree_add_51_79_groupi_n_6767;
  wire csa_tree_add_51_79_groupi_n_6768, csa_tree_add_51_79_groupi_n_6769, csa_tree_add_51_79_groupi_n_6770, csa_tree_add_51_79_groupi_n_6771, csa_tree_add_51_79_groupi_n_6772, csa_tree_add_51_79_groupi_n_6773, csa_tree_add_51_79_groupi_n_6774, csa_tree_add_51_79_groupi_n_6775;
  wire csa_tree_add_51_79_groupi_n_6776, csa_tree_add_51_79_groupi_n_6777, csa_tree_add_51_79_groupi_n_6778, csa_tree_add_51_79_groupi_n_6779, csa_tree_add_51_79_groupi_n_6780, csa_tree_add_51_79_groupi_n_6781, csa_tree_add_51_79_groupi_n_6782, csa_tree_add_51_79_groupi_n_6783;
  wire csa_tree_add_51_79_groupi_n_6784, csa_tree_add_51_79_groupi_n_6785, csa_tree_add_51_79_groupi_n_6786, csa_tree_add_51_79_groupi_n_6787, csa_tree_add_51_79_groupi_n_6788, csa_tree_add_51_79_groupi_n_6789, csa_tree_add_51_79_groupi_n_6790, csa_tree_add_51_79_groupi_n_6791;
  wire csa_tree_add_51_79_groupi_n_6792, csa_tree_add_51_79_groupi_n_6793, csa_tree_add_51_79_groupi_n_6794, csa_tree_add_51_79_groupi_n_6795, csa_tree_add_51_79_groupi_n_6796, csa_tree_add_51_79_groupi_n_6797, csa_tree_add_51_79_groupi_n_6798, csa_tree_add_51_79_groupi_n_6799;
  wire csa_tree_add_51_79_groupi_n_6800, csa_tree_add_51_79_groupi_n_6801, csa_tree_add_51_79_groupi_n_6802, csa_tree_add_51_79_groupi_n_6803, csa_tree_add_51_79_groupi_n_6804, csa_tree_add_51_79_groupi_n_6805, csa_tree_add_51_79_groupi_n_6806, csa_tree_add_51_79_groupi_n_6807;
  wire csa_tree_add_51_79_groupi_n_6808, csa_tree_add_51_79_groupi_n_6809, csa_tree_add_51_79_groupi_n_6810, csa_tree_add_51_79_groupi_n_6811, csa_tree_add_51_79_groupi_n_6812, csa_tree_add_51_79_groupi_n_6813, csa_tree_add_51_79_groupi_n_6814, csa_tree_add_51_79_groupi_n_6815;
  wire csa_tree_add_51_79_groupi_n_6816, csa_tree_add_51_79_groupi_n_6817, csa_tree_add_51_79_groupi_n_6818, csa_tree_add_51_79_groupi_n_6819, csa_tree_add_51_79_groupi_n_6820, csa_tree_add_51_79_groupi_n_6821, csa_tree_add_51_79_groupi_n_6822, csa_tree_add_51_79_groupi_n_6823;
  wire csa_tree_add_51_79_groupi_n_6824, csa_tree_add_51_79_groupi_n_6825, csa_tree_add_51_79_groupi_n_6826, csa_tree_add_51_79_groupi_n_6827, csa_tree_add_51_79_groupi_n_6828, csa_tree_add_51_79_groupi_n_6829, csa_tree_add_51_79_groupi_n_6830, csa_tree_add_51_79_groupi_n_6831;
  wire csa_tree_add_51_79_groupi_n_6832, csa_tree_add_51_79_groupi_n_6833, csa_tree_add_51_79_groupi_n_6834, csa_tree_add_51_79_groupi_n_6835, csa_tree_add_51_79_groupi_n_6836, csa_tree_add_51_79_groupi_n_6837, csa_tree_add_51_79_groupi_n_6838, csa_tree_add_51_79_groupi_n_6839;
  wire csa_tree_add_51_79_groupi_n_6840, csa_tree_add_51_79_groupi_n_6841, csa_tree_add_51_79_groupi_n_6842, csa_tree_add_51_79_groupi_n_6843, csa_tree_add_51_79_groupi_n_6844, csa_tree_add_51_79_groupi_n_6845, csa_tree_add_51_79_groupi_n_6846, csa_tree_add_51_79_groupi_n_6847;
  wire csa_tree_add_51_79_groupi_n_6848, csa_tree_add_51_79_groupi_n_6849, csa_tree_add_51_79_groupi_n_6850, csa_tree_add_51_79_groupi_n_6851, csa_tree_add_51_79_groupi_n_6852, csa_tree_add_51_79_groupi_n_6853, csa_tree_add_51_79_groupi_n_6854, csa_tree_add_51_79_groupi_n_6855;
  wire csa_tree_add_51_79_groupi_n_6856, csa_tree_add_51_79_groupi_n_6857, csa_tree_add_51_79_groupi_n_6858, csa_tree_add_51_79_groupi_n_6859, csa_tree_add_51_79_groupi_n_6860, csa_tree_add_51_79_groupi_n_6861, csa_tree_add_51_79_groupi_n_6862, csa_tree_add_51_79_groupi_n_6863;
  wire csa_tree_add_51_79_groupi_n_6864, csa_tree_add_51_79_groupi_n_6865, csa_tree_add_51_79_groupi_n_6866, csa_tree_add_51_79_groupi_n_6867, csa_tree_add_51_79_groupi_n_6868, csa_tree_add_51_79_groupi_n_6869, csa_tree_add_51_79_groupi_n_6870, csa_tree_add_51_79_groupi_n_6871;
  wire csa_tree_add_51_79_groupi_n_6872, csa_tree_add_51_79_groupi_n_6873, csa_tree_add_51_79_groupi_n_6874, csa_tree_add_51_79_groupi_n_6875, csa_tree_add_51_79_groupi_n_6876, csa_tree_add_51_79_groupi_n_6877, csa_tree_add_51_79_groupi_n_6878, csa_tree_add_51_79_groupi_n_6879;
  wire csa_tree_add_51_79_groupi_n_6880, csa_tree_add_51_79_groupi_n_6881, csa_tree_add_51_79_groupi_n_6882, csa_tree_add_51_79_groupi_n_6883, csa_tree_add_51_79_groupi_n_6884, csa_tree_add_51_79_groupi_n_6885, csa_tree_add_51_79_groupi_n_6886, csa_tree_add_51_79_groupi_n_6887;
  wire csa_tree_add_51_79_groupi_n_6888, csa_tree_add_51_79_groupi_n_6889, csa_tree_add_51_79_groupi_n_6890, csa_tree_add_51_79_groupi_n_6891, csa_tree_add_51_79_groupi_n_6892, csa_tree_add_51_79_groupi_n_6893, csa_tree_add_51_79_groupi_n_6894, csa_tree_add_51_79_groupi_n_6895;
  wire csa_tree_add_51_79_groupi_n_6896, csa_tree_add_51_79_groupi_n_6897, csa_tree_add_51_79_groupi_n_6898, csa_tree_add_51_79_groupi_n_6899, csa_tree_add_51_79_groupi_n_6900, csa_tree_add_51_79_groupi_n_6901, csa_tree_add_51_79_groupi_n_6902, csa_tree_add_51_79_groupi_n_6903;
  wire csa_tree_add_51_79_groupi_n_6904, csa_tree_add_51_79_groupi_n_6905, csa_tree_add_51_79_groupi_n_6906, csa_tree_add_51_79_groupi_n_6907, csa_tree_add_51_79_groupi_n_6908, csa_tree_add_51_79_groupi_n_6909, csa_tree_add_51_79_groupi_n_6910, csa_tree_add_51_79_groupi_n_6911;
  wire csa_tree_add_51_79_groupi_n_6912, csa_tree_add_51_79_groupi_n_6913, csa_tree_add_51_79_groupi_n_6914, csa_tree_add_51_79_groupi_n_6915, csa_tree_add_51_79_groupi_n_6916, csa_tree_add_51_79_groupi_n_6917, csa_tree_add_51_79_groupi_n_6918, csa_tree_add_51_79_groupi_n_6919;
  wire csa_tree_add_51_79_groupi_n_6920, csa_tree_add_51_79_groupi_n_6921, csa_tree_add_51_79_groupi_n_6922, csa_tree_add_51_79_groupi_n_6923, csa_tree_add_51_79_groupi_n_6924, csa_tree_add_51_79_groupi_n_6925, csa_tree_add_51_79_groupi_n_6926, csa_tree_add_51_79_groupi_n_6927;
  wire csa_tree_add_51_79_groupi_n_6928, csa_tree_add_51_79_groupi_n_6929, csa_tree_add_51_79_groupi_n_6930, csa_tree_add_51_79_groupi_n_6931, csa_tree_add_51_79_groupi_n_6932, csa_tree_add_51_79_groupi_n_6933, csa_tree_add_51_79_groupi_n_6934, csa_tree_add_51_79_groupi_n_6935;
  wire csa_tree_add_51_79_groupi_n_6936, csa_tree_add_51_79_groupi_n_6937, csa_tree_add_51_79_groupi_n_6938, csa_tree_add_51_79_groupi_n_6939, csa_tree_add_51_79_groupi_n_6940, csa_tree_add_51_79_groupi_n_6941, csa_tree_add_51_79_groupi_n_6942, csa_tree_add_51_79_groupi_n_6943;
  wire csa_tree_add_51_79_groupi_n_6944, csa_tree_add_51_79_groupi_n_6945, csa_tree_add_51_79_groupi_n_6946, csa_tree_add_51_79_groupi_n_6947, csa_tree_add_51_79_groupi_n_6948, csa_tree_add_51_79_groupi_n_6949, csa_tree_add_51_79_groupi_n_6950, csa_tree_add_51_79_groupi_n_6951;
  wire csa_tree_add_51_79_groupi_n_6952, csa_tree_add_51_79_groupi_n_6953, csa_tree_add_51_79_groupi_n_6954, csa_tree_add_51_79_groupi_n_6955, csa_tree_add_51_79_groupi_n_6956, csa_tree_add_51_79_groupi_n_6957, csa_tree_add_51_79_groupi_n_6958, csa_tree_add_51_79_groupi_n_6959;
  wire csa_tree_add_51_79_groupi_n_6960, csa_tree_add_51_79_groupi_n_6961, csa_tree_add_51_79_groupi_n_6962, csa_tree_add_51_79_groupi_n_6963, csa_tree_add_51_79_groupi_n_6964, csa_tree_add_51_79_groupi_n_6965, csa_tree_add_51_79_groupi_n_6966, csa_tree_add_51_79_groupi_n_6967;
  wire csa_tree_add_51_79_groupi_n_6968, csa_tree_add_51_79_groupi_n_6969, csa_tree_add_51_79_groupi_n_6970, csa_tree_add_51_79_groupi_n_6971, csa_tree_add_51_79_groupi_n_6972, csa_tree_add_51_79_groupi_n_6973, csa_tree_add_51_79_groupi_n_6974, csa_tree_add_51_79_groupi_n_6975;
  wire csa_tree_add_51_79_groupi_n_6976, csa_tree_add_51_79_groupi_n_6977, csa_tree_add_51_79_groupi_n_6978, csa_tree_add_51_79_groupi_n_6979, csa_tree_add_51_79_groupi_n_6980, csa_tree_add_51_79_groupi_n_6981, csa_tree_add_51_79_groupi_n_6982, csa_tree_add_51_79_groupi_n_6983;
  wire csa_tree_add_51_79_groupi_n_6984, csa_tree_add_51_79_groupi_n_6985, csa_tree_add_51_79_groupi_n_6986, csa_tree_add_51_79_groupi_n_6987, csa_tree_add_51_79_groupi_n_6988, csa_tree_add_51_79_groupi_n_6989, csa_tree_add_51_79_groupi_n_6990, csa_tree_add_51_79_groupi_n_6991;
  wire csa_tree_add_51_79_groupi_n_6992, csa_tree_add_51_79_groupi_n_6993, csa_tree_add_51_79_groupi_n_6994, csa_tree_add_51_79_groupi_n_6995, csa_tree_add_51_79_groupi_n_6996, csa_tree_add_51_79_groupi_n_6997, csa_tree_add_51_79_groupi_n_6998, csa_tree_add_51_79_groupi_n_6999;
  wire csa_tree_add_51_79_groupi_n_7000, csa_tree_add_51_79_groupi_n_7001, csa_tree_add_51_79_groupi_n_7002, csa_tree_add_51_79_groupi_n_7003, csa_tree_add_51_79_groupi_n_7004, csa_tree_add_51_79_groupi_n_7005, csa_tree_add_51_79_groupi_n_7006, csa_tree_add_51_79_groupi_n_7007;
  wire csa_tree_add_51_79_groupi_n_7008, csa_tree_add_51_79_groupi_n_7009, csa_tree_add_51_79_groupi_n_7010, csa_tree_add_51_79_groupi_n_7011, csa_tree_add_51_79_groupi_n_7012, csa_tree_add_51_79_groupi_n_7013, csa_tree_add_51_79_groupi_n_7014, csa_tree_add_51_79_groupi_n_7015;
  wire csa_tree_add_51_79_groupi_n_7016, csa_tree_add_51_79_groupi_n_7017, csa_tree_add_51_79_groupi_n_7018, csa_tree_add_51_79_groupi_n_7019, csa_tree_add_51_79_groupi_n_7020, csa_tree_add_51_79_groupi_n_7021, csa_tree_add_51_79_groupi_n_7022, csa_tree_add_51_79_groupi_n_7023;
  wire csa_tree_add_51_79_groupi_n_7024, csa_tree_add_51_79_groupi_n_7025, csa_tree_add_51_79_groupi_n_7026, csa_tree_add_51_79_groupi_n_7027, csa_tree_add_51_79_groupi_n_7028, csa_tree_add_51_79_groupi_n_7029, csa_tree_add_51_79_groupi_n_7030, csa_tree_add_51_79_groupi_n_7031;
  wire csa_tree_add_51_79_groupi_n_7032, csa_tree_add_51_79_groupi_n_7033, csa_tree_add_51_79_groupi_n_7034, csa_tree_add_51_79_groupi_n_7035, csa_tree_add_51_79_groupi_n_7036, csa_tree_add_51_79_groupi_n_7037, csa_tree_add_51_79_groupi_n_7038, csa_tree_add_51_79_groupi_n_7039;
  wire csa_tree_add_51_79_groupi_n_7040, csa_tree_add_51_79_groupi_n_7041, csa_tree_add_51_79_groupi_n_7042, csa_tree_add_51_79_groupi_n_7043, csa_tree_add_51_79_groupi_n_7044, csa_tree_add_51_79_groupi_n_7045, csa_tree_add_51_79_groupi_n_7046, csa_tree_add_51_79_groupi_n_7047;
  wire csa_tree_add_51_79_groupi_n_7048, csa_tree_add_51_79_groupi_n_7049, csa_tree_add_51_79_groupi_n_7050, csa_tree_add_51_79_groupi_n_7051, csa_tree_add_51_79_groupi_n_7052, csa_tree_add_51_79_groupi_n_7053, csa_tree_add_51_79_groupi_n_7054, csa_tree_add_51_79_groupi_n_7055;
  wire csa_tree_add_51_79_groupi_n_7056, csa_tree_add_51_79_groupi_n_7057, csa_tree_add_51_79_groupi_n_7058, csa_tree_add_51_79_groupi_n_7059, csa_tree_add_51_79_groupi_n_7060, csa_tree_add_51_79_groupi_n_7061, csa_tree_add_51_79_groupi_n_7062, csa_tree_add_51_79_groupi_n_7063;
  wire csa_tree_add_51_79_groupi_n_7064, csa_tree_add_51_79_groupi_n_7065, csa_tree_add_51_79_groupi_n_7066, csa_tree_add_51_79_groupi_n_7067, csa_tree_add_51_79_groupi_n_7068, csa_tree_add_51_79_groupi_n_7069, csa_tree_add_51_79_groupi_n_7070, csa_tree_add_51_79_groupi_n_7071;
  wire csa_tree_add_51_79_groupi_n_7072, csa_tree_add_51_79_groupi_n_7073, csa_tree_add_51_79_groupi_n_7074, csa_tree_add_51_79_groupi_n_7075, csa_tree_add_51_79_groupi_n_7076, csa_tree_add_51_79_groupi_n_7077, csa_tree_add_51_79_groupi_n_7078, csa_tree_add_51_79_groupi_n_7079;
  wire csa_tree_add_51_79_groupi_n_7080, csa_tree_add_51_79_groupi_n_7081, csa_tree_add_51_79_groupi_n_7082, csa_tree_add_51_79_groupi_n_7083, csa_tree_add_51_79_groupi_n_7084, csa_tree_add_51_79_groupi_n_7085, csa_tree_add_51_79_groupi_n_7086, csa_tree_add_51_79_groupi_n_7087;
  wire csa_tree_add_51_79_groupi_n_7088, csa_tree_add_51_79_groupi_n_7089, csa_tree_add_51_79_groupi_n_7090, csa_tree_add_51_79_groupi_n_7091, csa_tree_add_51_79_groupi_n_7092, csa_tree_add_51_79_groupi_n_7093, csa_tree_add_51_79_groupi_n_7094, csa_tree_add_51_79_groupi_n_7095;
  wire csa_tree_add_51_79_groupi_n_7096, csa_tree_add_51_79_groupi_n_7097, csa_tree_add_51_79_groupi_n_7098, csa_tree_add_51_79_groupi_n_7099, csa_tree_add_51_79_groupi_n_7100, csa_tree_add_51_79_groupi_n_7101, csa_tree_add_51_79_groupi_n_7102, csa_tree_add_51_79_groupi_n_7103;
  wire csa_tree_add_51_79_groupi_n_7104, csa_tree_add_51_79_groupi_n_7105, csa_tree_add_51_79_groupi_n_7106, csa_tree_add_51_79_groupi_n_7107, csa_tree_add_51_79_groupi_n_7108, csa_tree_add_51_79_groupi_n_7109, csa_tree_add_51_79_groupi_n_7110, csa_tree_add_51_79_groupi_n_7111;
  wire csa_tree_add_51_79_groupi_n_7112, csa_tree_add_51_79_groupi_n_7113, csa_tree_add_51_79_groupi_n_7114, csa_tree_add_51_79_groupi_n_7115, csa_tree_add_51_79_groupi_n_7116, csa_tree_add_51_79_groupi_n_7117, csa_tree_add_51_79_groupi_n_7118, csa_tree_add_51_79_groupi_n_7119;
  wire csa_tree_add_51_79_groupi_n_7120, csa_tree_add_51_79_groupi_n_7121, csa_tree_add_51_79_groupi_n_7122, csa_tree_add_51_79_groupi_n_7123, csa_tree_add_51_79_groupi_n_7124, csa_tree_add_51_79_groupi_n_7125, csa_tree_add_51_79_groupi_n_7126, csa_tree_add_51_79_groupi_n_7127;
  wire csa_tree_add_51_79_groupi_n_7128, csa_tree_add_51_79_groupi_n_7129, csa_tree_add_51_79_groupi_n_7130, csa_tree_add_51_79_groupi_n_7131, csa_tree_add_51_79_groupi_n_7132, csa_tree_add_51_79_groupi_n_7133, csa_tree_add_51_79_groupi_n_7134, csa_tree_add_51_79_groupi_n_7135;
  wire csa_tree_add_51_79_groupi_n_7136, csa_tree_add_51_79_groupi_n_7137, csa_tree_add_51_79_groupi_n_7138, csa_tree_add_51_79_groupi_n_7139, csa_tree_add_51_79_groupi_n_7140, csa_tree_add_51_79_groupi_n_7141, csa_tree_add_51_79_groupi_n_7142, csa_tree_add_51_79_groupi_n_7143;
  wire csa_tree_add_51_79_groupi_n_7144, csa_tree_add_51_79_groupi_n_7145, csa_tree_add_51_79_groupi_n_7146, csa_tree_add_51_79_groupi_n_7147, csa_tree_add_51_79_groupi_n_7148, csa_tree_add_51_79_groupi_n_7149, csa_tree_add_51_79_groupi_n_7150, csa_tree_add_51_79_groupi_n_7151;
  wire csa_tree_add_51_79_groupi_n_7152, csa_tree_add_51_79_groupi_n_7153, csa_tree_add_51_79_groupi_n_7154, csa_tree_add_51_79_groupi_n_7155, csa_tree_add_51_79_groupi_n_7156, csa_tree_add_51_79_groupi_n_7157, csa_tree_add_51_79_groupi_n_7158, csa_tree_add_51_79_groupi_n_7159;
  wire csa_tree_add_51_79_groupi_n_7160, csa_tree_add_51_79_groupi_n_7161, csa_tree_add_51_79_groupi_n_7162, csa_tree_add_51_79_groupi_n_7163, csa_tree_add_51_79_groupi_n_7164, csa_tree_add_51_79_groupi_n_7165, csa_tree_add_51_79_groupi_n_7166, csa_tree_add_51_79_groupi_n_7167;
  wire csa_tree_add_51_79_groupi_n_7168, csa_tree_add_51_79_groupi_n_7169, csa_tree_add_51_79_groupi_n_7170, csa_tree_add_51_79_groupi_n_7171, csa_tree_add_51_79_groupi_n_7172, csa_tree_add_51_79_groupi_n_7173, csa_tree_add_51_79_groupi_n_7174, csa_tree_add_51_79_groupi_n_7175;
  wire csa_tree_add_51_79_groupi_n_7176, csa_tree_add_51_79_groupi_n_7177, csa_tree_add_51_79_groupi_n_7178, csa_tree_add_51_79_groupi_n_7179, csa_tree_add_51_79_groupi_n_7180, csa_tree_add_51_79_groupi_n_7181, csa_tree_add_51_79_groupi_n_7182, csa_tree_add_51_79_groupi_n_7183;
  wire csa_tree_add_51_79_groupi_n_7184, csa_tree_add_51_79_groupi_n_7185, csa_tree_add_51_79_groupi_n_7186, csa_tree_add_51_79_groupi_n_7187, csa_tree_add_51_79_groupi_n_7188, csa_tree_add_51_79_groupi_n_7189, csa_tree_add_51_79_groupi_n_7190, csa_tree_add_51_79_groupi_n_7191;
  wire csa_tree_add_51_79_groupi_n_7192, csa_tree_add_51_79_groupi_n_7193, csa_tree_add_51_79_groupi_n_7194, csa_tree_add_51_79_groupi_n_7195, csa_tree_add_51_79_groupi_n_7196, csa_tree_add_51_79_groupi_n_7197, csa_tree_add_51_79_groupi_n_7198, csa_tree_add_51_79_groupi_n_7199;
  wire csa_tree_add_51_79_groupi_n_7200, csa_tree_add_51_79_groupi_n_7201, csa_tree_add_51_79_groupi_n_7202, csa_tree_add_51_79_groupi_n_7203, csa_tree_add_51_79_groupi_n_7204, csa_tree_add_51_79_groupi_n_7205, csa_tree_add_51_79_groupi_n_7206, csa_tree_add_51_79_groupi_n_7207;
  wire csa_tree_add_51_79_groupi_n_7208, csa_tree_add_51_79_groupi_n_7209, csa_tree_add_51_79_groupi_n_7210, csa_tree_add_51_79_groupi_n_7211, csa_tree_add_51_79_groupi_n_7212, csa_tree_add_51_79_groupi_n_7213, csa_tree_add_51_79_groupi_n_7214, csa_tree_add_51_79_groupi_n_7215;
  wire csa_tree_add_51_79_groupi_n_7216, csa_tree_add_51_79_groupi_n_7217, csa_tree_add_51_79_groupi_n_7218, csa_tree_add_51_79_groupi_n_7219, csa_tree_add_51_79_groupi_n_7220, csa_tree_add_51_79_groupi_n_7221, csa_tree_add_51_79_groupi_n_7222, csa_tree_add_51_79_groupi_n_7223;
  wire csa_tree_add_51_79_groupi_n_7224, csa_tree_add_51_79_groupi_n_7225, csa_tree_add_51_79_groupi_n_7226, csa_tree_add_51_79_groupi_n_7227, csa_tree_add_51_79_groupi_n_7228, csa_tree_add_51_79_groupi_n_7229, csa_tree_add_51_79_groupi_n_7230, csa_tree_add_51_79_groupi_n_7231;
  wire csa_tree_add_51_79_groupi_n_7232, csa_tree_add_51_79_groupi_n_7233, csa_tree_add_51_79_groupi_n_7234, csa_tree_add_51_79_groupi_n_7235, csa_tree_add_51_79_groupi_n_7236, csa_tree_add_51_79_groupi_n_7237, csa_tree_add_51_79_groupi_n_7238, csa_tree_add_51_79_groupi_n_7239;
  wire csa_tree_add_51_79_groupi_n_7240, csa_tree_add_51_79_groupi_n_7241, csa_tree_add_51_79_groupi_n_7242, csa_tree_add_51_79_groupi_n_7243, csa_tree_add_51_79_groupi_n_7244, csa_tree_add_51_79_groupi_n_7245, csa_tree_add_51_79_groupi_n_7246, csa_tree_add_51_79_groupi_n_7247;
  wire csa_tree_add_51_79_groupi_n_7248, csa_tree_add_51_79_groupi_n_7249, csa_tree_add_51_79_groupi_n_7250, csa_tree_add_51_79_groupi_n_7251, csa_tree_add_51_79_groupi_n_7252, csa_tree_add_51_79_groupi_n_7253, csa_tree_add_51_79_groupi_n_7254, csa_tree_add_51_79_groupi_n_7255;
  wire csa_tree_add_51_79_groupi_n_7256, csa_tree_add_51_79_groupi_n_7257, csa_tree_add_51_79_groupi_n_7258, csa_tree_add_51_79_groupi_n_7259, csa_tree_add_51_79_groupi_n_7260, csa_tree_add_51_79_groupi_n_7261, csa_tree_add_51_79_groupi_n_7262, csa_tree_add_51_79_groupi_n_7263;
  wire csa_tree_add_51_79_groupi_n_7264, csa_tree_add_51_79_groupi_n_7265, csa_tree_add_51_79_groupi_n_7266, csa_tree_add_51_79_groupi_n_7267, csa_tree_add_51_79_groupi_n_7268, csa_tree_add_51_79_groupi_n_7269, csa_tree_add_51_79_groupi_n_7270, csa_tree_add_51_79_groupi_n_7271;
  wire csa_tree_add_51_79_groupi_n_7272, csa_tree_add_51_79_groupi_n_7273, csa_tree_add_51_79_groupi_n_7274, csa_tree_add_51_79_groupi_n_7275, csa_tree_add_51_79_groupi_n_7276, csa_tree_add_51_79_groupi_n_7277, csa_tree_add_51_79_groupi_n_7278, csa_tree_add_51_79_groupi_n_7279;
  wire csa_tree_add_51_79_groupi_n_7280, csa_tree_add_51_79_groupi_n_7281, csa_tree_add_51_79_groupi_n_7282, csa_tree_add_51_79_groupi_n_7283, csa_tree_add_51_79_groupi_n_7284, csa_tree_add_51_79_groupi_n_7285, csa_tree_add_51_79_groupi_n_7286, csa_tree_add_51_79_groupi_n_7287;
  wire csa_tree_add_51_79_groupi_n_7288, csa_tree_add_51_79_groupi_n_7289, csa_tree_add_51_79_groupi_n_7290, csa_tree_add_51_79_groupi_n_7291, csa_tree_add_51_79_groupi_n_7292, csa_tree_add_51_79_groupi_n_7293, csa_tree_add_51_79_groupi_n_7294, csa_tree_add_51_79_groupi_n_7295;
  wire csa_tree_add_51_79_groupi_n_7296, csa_tree_add_51_79_groupi_n_7297, csa_tree_add_51_79_groupi_n_7298, csa_tree_add_51_79_groupi_n_7299, csa_tree_add_51_79_groupi_n_7300, csa_tree_add_51_79_groupi_n_7301, csa_tree_add_51_79_groupi_n_7302, csa_tree_add_51_79_groupi_n_7303;
  wire csa_tree_add_51_79_groupi_n_7304, csa_tree_add_51_79_groupi_n_7305, csa_tree_add_51_79_groupi_n_7306, csa_tree_add_51_79_groupi_n_7307, csa_tree_add_51_79_groupi_n_7308, csa_tree_add_51_79_groupi_n_7309, csa_tree_add_51_79_groupi_n_7310, csa_tree_add_51_79_groupi_n_7311;
  wire csa_tree_add_51_79_groupi_n_7312, csa_tree_add_51_79_groupi_n_7313, csa_tree_add_51_79_groupi_n_7314, csa_tree_add_51_79_groupi_n_7315, csa_tree_add_51_79_groupi_n_7316, csa_tree_add_51_79_groupi_n_7317, csa_tree_add_51_79_groupi_n_7318, csa_tree_add_51_79_groupi_n_7319;
  wire csa_tree_add_51_79_groupi_n_7320, csa_tree_add_51_79_groupi_n_7321, csa_tree_add_51_79_groupi_n_7322, csa_tree_add_51_79_groupi_n_7323, csa_tree_add_51_79_groupi_n_7324, csa_tree_add_51_79_groupi_n_7325, csa_tree_add_51_79_groupi_n_7326, csa_tree_add_51_79_groupi_n_7327;
  wire csa_tree_add_51_79_groupi_n_7328, csa_tree_add_51_79_groupi_n_7329, csa_tree_add_51_79_groupi_n_7330, csa_tree_add_51_79_groupi_n_7331, csa_tree_add_51_79_groupi_n_7332, csa_tree_add_51_79_groupi_n_7333, csa_tree_add_51_79_groupi_n_7334, csa_tree_add_51_79_groupi_n_7335;
  wire csa_tree_add_51_79_groupi_n_7336, csa_tree_add_51_79_groupi_n_7337, csa_tree_add_51_79_groupi_n_7338, csa_tree_add_51_79_groupi_n_7339, csa_tree_add_51_79_groupi_n_7340, csa_tree_add_51_79_groupi_n_7341, csa_tree_add_51_79_groupi_n_7342, csa_tree_add_51_79_groupi_n_7343;
  wire csa_tree_add_51_79_groupi_n_7344, csa_tree_add_51_79_groupi_n_7345, csa_tree_add_51_79_groupi_n_7346, csa_tree_add_51_79_groupi_n_7347, csa_tree_add_51_79_groupi_n_7348, csa_tree_add_51_79_groupi_n_7349, csa_tree_add_51_79_groupi_n_7350, csa_tree_add_51_79_groupi_n_7351;
  wire csa_tree_add_51_79_groupi_n_7352, csa_tree_add_51_79_groupi_n_7353, csa_tree_add_51_79_groupi_n_7354, csa_tree_add_51_79_groupi_n_7355, csa_tree_add_51_79_groupi_n_7356, csa_tree_add_51_79_groupi_n_7357, csa_tree_add_51_79_groupi_n_7358, csa_tree_add_51_79_groupi_n_7359;
  wire csa_tree_add_51_79_groupi_n_7360, csa_tree_add_51_79_groupi_n_7361, csa_tree_add_51_79_groupi_n_7362, csa_tree_add_51_79_groupi_n_7363, csa_tree_add_51_79_groupi_n_7364, csa_tree_add_51_79_groupi_n_7365, csa_tree_add_51_79_groupi_n_7366, csa_tree_add_51_79_groupi_n_7367;
  wire csa_tree_add_51_79_groupi_n_7368, csa_tree_add_51_79_groupi_n_7369, csa_tree_add_51_79_groupi_n_7370, csa_tree_add_51_79_groupi_n_7371, csa_tree_add_51_79_groupi_n_7372, csa_tree_add_51_79_groupi_n_7373, csa_tree_add_51_79_groupi_n_7374, csa_tree_add_51_79_groupi_n_7375;
  wire csa_tree_add_51_79_groupi_n_7376, csa_tree_add_51_79_groupi_n_7377, csa_tree_add_51_79_groupi_n_7378, csa_tree_add_51_79_groupi_n_7379, csa_tree_add_51_79_groupi_n_7380, csa_tree_add_51_79_groupi_n_7381, csa_tree_add_51_79_groupi_n_7382, csa_tree_add_51_79_groupi_n_7383;
  wire csa_tree_add_51_79_groupi_n_7384, csa_tree_add_51_79_groupi_n_7385, csa_tree_add_51_79_groupi_n_7386, csa_tree_add_51_79_groupi_n_7387, csa_tree_add_51_79_groupi_n_7388, csa_tree_add_51_79_groupi_n_7389, csa_tree_add_51_79_groupi_n_7390, csa_tree_add_51_79_groupi_n_7391;
  wire csa_tree_add_51_79_groupi_n_7392, csa_tree_add_51_79_groupi_n_7393, csa_tree_add_51_79_groupi_n_7394, csa_tree_add_51_79_groupi_n_7395, csa_tree_add_51_79_groupi_n_7396, csa_tree_add_51_79_groupi_n_7397, csa_tree_add_51_79_groupi_n_7398, csa_tree_add_51_79_groupi_n_7399;
  wire csa_tree_add_51_79_groupi_n_7400, csa_tree_add_51_79_groupi_n_7401, csa_tree_add_51_79_groupi_n_7402, csa_tree_add_51_79_groupi_n_7403, csa_tree_add_51_79_groupi_n_7404, csa_tree_add_51_79_groupi_n_7405, csa_tree_add_51_79_groupi_n_7406, csa_tree_add_51_79_groupi_n_7407;
  wire csa_tree_add_51_79_groupi_n_7408, csa_tree_add_51_79_groupi_n_7409, csa_tree_add_51_79_groupi_n_7410, csa_tree_add_51_79_groupi_n_7411, csa_tree_add_51_79_groupi_n_7412, csa_tree_add_51_79_groupi_n_7413, csa_tree_add_51_79_groupi_n_7414, csa_tree_add_51_79_groupi_n_7415;
  wire csa_tree_add_51_79_groupi_n_7416, csa_tree_add_51_79_groupi_n_7417, csa_tree_add_51_79_groupi_n_7418, csa_tree_add_51_79_groupi_n_7419, csa_tree_add_51_79_groupi_n_7420, csa_tree_add_51_79_groupi_n_7421, csa_tree_add_51_79_groupi_n_7422, csa_tree_add_51_79_groupi_n_7423;
  wire csa_tree_add_51_79_groupi_n_7424, csa_tree_add_51_79_groupi_n_7425, csa_tree_add_51_79_groupi_n_7426, csa_tree_add_51_79_groupi_n_7427, csa_tree_add_51_79_groupi_n_7428, csa_tree_add_51_79_groupi_n_7429, csa_tree_add_51_79_groupi_n_7430, csa_tree_add_51_79_groupi_n_7431;
  wire csa_tree_add_51_79_groupi_n_7432, csa_tree_add_51_79_groupi_n_7433, csa_tree_add_51_79_groupi_n_7434, csa_tree_add_51_79_groupi_n_7435, csa_tree_add_51_79_groupi_n_7436, csa_tree_add_51_79_groupi_n_7437, csa_tree_add_51_79_groupi_n_7438, csa_tree_add_51_79_groupi_n_7439;
  wire csa_tree_add_51_79_groupi_n_7440, csa_tree_add_51_79_groupi_n_7441, csa_tree_add_51_79_groupi_n_7442, csa_tree_add_51_79_groupi_n_7443, csa_tree_add_51_79_groupi_n_7444, csa_tree_add_51_79_groupi_n_7445, csa_tree_add_51_79_groupi_n_7446, csa_tree_add_51_79_groupi_n_7447;
  wire csa_tree_add_51_79_groupi_n_7448, csa_tree_add_51_79_groupi_n_7449, csa_tree_add_51_79_groupi_n_7450, csa_tree_add_51_79_groupi_n_7451, csa_tree_add_51_79_groupi_n_7452, csa_tree_add_51_79_groupi_n_7453, csa_tree_add_51_79_groupi_n_7454, csa_tree_add_51_79_groupi_n_7455;
  wire csa_tree_add_51_79_groupi_n_7456, csa_tree_add_51_79_groupi_n_7457, csa_tree_add_51_79_groupi_n_7458, csa_tree_add_51_79_groupi_n_7459, csa_tree_add_51_79_groupi_n_7460, csa_tree_add_51_79_groupi_n_7461, csa_tree_add_51_79_groupi_n_7462, csa_tree_add_51_79_groupi_n_7463;
  wire csa_tree_add_51_79_groupi_n_7464, csa_tree_add_51_79_groupi_n_7465, csa_tree_add_51_79_groupi_n_7466, csa_tree_add_51_79_groupi_n_7467, csa_tree_add_51_79_groupi_n_7468, csa_tree_add_51_79_groupi_n_7469, csa_tree_add_51_79_groupi_n_7470, csa_tree_add_51_79_groupi_n_7471;
  wire csa_tree_add_51_79_groupi_n_7472, csa_tree_add_51_79_groupi_n_7473, csa_tree_add_51_79_groupi_n_7474, csa_tree_add_51_79_groupi_n_7475, csa_tree_add_51_79_groupi_n_7476, csa_tree_add_51_79_groupi_n_7477, csa_tree_add_51_79_groupi_n_7478, csa_tree_add_51_79_groupi_n_7479;
  wire csa_tree_add_51_79_groupi_n_7480, csa_tree_add_51_79_groupi_n_7481, csa_tree_add_51_79_groupi_n_7482, csa_tree_add_51_79_groupi_n_7483, csa_tree_add_51_79_groupi_n_7484, csa_tree_add_51_79_groupi_n_7485, csa_tree_add_51_79_groupi_n_7486, csa_tree_add_51_79_groupi_n_7487;
  wire csa_tree_add_51_79_groupi_n_7488, csa_tree_add_51_79_groupi_n_7489, csa_tree_add_51_79_groupi_n_7490, csa_tree_add_51_79_groupi_n_7491, csa_tree_add_51_79_groupi_n_7492, csa_tree_add_51_79_groupi_n_7493, csa_tree_add_51_79_groupi_n_7494, csa_tree_add_51_79_groupi_n_7495;
  wire csa_tree_add_51_79_groupi_n_7496, csa_tree_add_51_79_groupi_n_7497, csa_tree_add_51_79_groupi_n_7498, csa_tree_add_51_79_groupi_n_7499, csa_tree_add_51_79_groupi_n_7500, csa_tree_add_51_79_groupi_n_7501, csa_tree_add_51_79_groupi_n_7502, csa_tree_add_51_79_groupi_n_7503;
  wire csa_tree_add_51_79_groupi_n_7504, csa_tree_add_51_79_groupi_n_7505, csa_tree_add_51_79_groupi_n_7506, csa_tree_add_51_79_groupi_n_7507, csa_tree_add_51_79_groupi_n_7508, csa_tree_add_51_79_groupi_n_7509, csa_tree_add_51_79_groupi_n_7510, csa_tree_add_51_79_groupi_n_7511;
  wire csa_tree_add_51_79_groupi_n_7512, csa_tree_add_51_79_groupi_n_7513, csa_tree_add_51_79_groupi_n_7514, csa_tree_add_51_79_groupi_n_7515, csa_tree_add_51_79_groupi_n_7516, csa_tree_add_51_79_groupi_n_7517, csa_tree_add_51_79_groupi_n_7518, csa_tree_add_51_79_groupi_n_7519;
  wire csa_tree_add_51_79_groupi_n_7520, csa_tree_add_51_79_groupi_n_7521, csa_tree_add_51_79_groupi_n_7522, csa_tree_add_51_79_groupi_n_7523, csa_tree_add_51_79_groupi_n_7524, csa_tree_add_51_79_groupi_n_7525, csa_tree_add_51_79_groupi_n_7526, csa_tree_add_51_79_groupi_n_7527;
  wire csa_tree_add_51_79_groupi_n_7528, csa_tree_add_51_79_groupi_n_7529, csa_tree_add_51_79_groupi_n_7530, csa_tree_add_51_79_groupi_n_7531, csa_tree_add_51_79_groupi_n_7532, csa_tree_add_51_79_groupi_n_7533, csa_tree_add_51_79_groupi_n_7534, csa_tree_add_51_79_groupi_n_7535;
  wire csa_tree_add_51_79_groupi_n_7536, csa_tree_add_51_79_groupi_n_7537, csa_tree_add_51_79_groupi_n_7538, csa_tree_add_51_79_groupi_n_7539, csa_tree_add_51_79_groupi_n_7540, csa_tree_add_51_79_groupi_n_7541, csa_tree_add_51_79_groupi_n_7542, csa_tree_add_51_79_groupi_n_7543;
  wire csa_tree_add_51_79_groupi_n_7544, csa_tree_add_51_79_groupi_n_7545, csa_tree_add_51_79_groupi_n_7546, csa_tree_add_51_79_groupi_n_7547, csa_tree_add_51_79_groupi_n_7548, csa_tree_add_51_79_groupi_n_7549, csa_tree_add_51_79_groupi_n_7550, csa_tree_add_51_79_groupi_n_7551;
  wire csa_tree_add_51_79_groupi_n_7552, csa_tree_add_51_79_groupi_n_7553, csa_tree_add_51_79_groupi_n_7554, csa_tree_add_51_79_groupi_n_7555, csa_tree_add_51_79_groupi_n_7556, csa_tree_add_51_79_groupi_n_7557, csa_tree_add_51_79_groupi_n_7558, csa_tree_add_51_79_groupi_n_7559;
  wire csa_tree_add_51_79_groupi_n_7560, csa_tree_add_51_79_groupi_n_7561, csa_tree_add_51_79_groupi_n_7562, csa_tree_add_51_79_groupi_n_7563, csa_tree_add_51_79_groupi_n_7564, csa_tree_add_51_79_groupi_n_7565, csa_tree_add_51_79_groupi_n_7566, csa_tree_add_51_79_groupi_n_7567;
  wire csa_tree_add_51_79_groupi_n_7568, csa_tree_add_51_79_groupi_n_7569, csa_tree_add_51_79_groupi_n_7570, csa_tree_add_51_79_groupi_n_7571, csa_tree_add_51_79_groupi_n_7572, csa_tree_add_51_79_groupi_n_7573, csa_tree_add_51_79_groupi_n_7574, csa_tree_add_51_79_groupi_n_7575;
  wire csa_tree_add_51_79_groupi_n_7576, csa_tree_add_51_79_groupi_n_7577, csa_tree_add_51_79_groupi_n_7578, csa_tree_add_51_79_groupi_n_7579, csa_tree_add_51_79_groupi_n_7580, csa_tree_add_51_79_groupi_n_7581, csa_tree_add_51_79_groupi_n_7582, csa_tree_add_51_79_groupi_n_7583;
  wire csa_tree_add_51_79_groupi_n_7584, csa_tree_add_51_79_groupi_n_7585, csa_tree_add_51_79_groupi_n_7586, csa_tree_add_51_79_groupi_n_7587, csa_tree_add_51_79_groupi_n_7588, csa_tree_add_51_79_groupi_n_7589, csa_tree_add_51_79_groupi_n_7590, csa_tree_add_51_79_groupi_n_7591;
  wire csa_tree_add_51_79_groupi_n_7592, csa_tree_add_51_79_groupi_n_7593, csa_tree_add_51_79_groupi_n_7594, csa_tree_add_51_79_groupi_n_7595, csa_tree_add_51_79_groupi_n_7596, csa_tree_add_51_79_groupi_n_7597, csa_tree_add_51_79_groupi_n_7598, csa_tree_add_51_79_groupi_n_7599;
  wire csa_tree_add_51_79_groupi_n_7600, csa_tree_add_51_79_groupi_n_7601, csa_tree_add_51_79_groupi_n_7602, csa_tree_add_51_79_groupi_n_7603, csa_tree_add_51_79_groupi_n_7604, csa_tree_add_51_79_groupi_n_7605, csa_tree_add_51_79_groupi_n_7606, csa_tree_add_51_79_groupi_n_7607;
  wire csa_tree_add_51_79_groupi_n_7608, csa_tree_add_51_79_groupi_n_7609, csa_tree_add_51_79_groupi_n_7610, csa_tree_add_51_79_groupi_n_7611, csa_tree_add_51_79_groupi_n_7612, csa_tree_add_51_79_groupi_n_7613, csa_tree_add_51_79_groupi_n_7614, csa_tree_add_51_79_groupi_n_7615;
  wire csa_tree_add_51_79_groupi_n_7616, csa_tree_add_51_79_groupi_n_7617, csa_tree_add_51_79_groupi_n_7618, csa_tree_add_51_79_groupi_n_7619, csa_tree_add_51_79_groupi_n_7620, csa_tree_add_51_79_groupi_n_7621, csa_tree_add_51_79_groupi_n_7622, csa_tree_add_51_79_groupi_n_7623;
  wire csa_tree_add_51_79_groupi_n_7624, csa_tree_add_51_79_groupi_n_7625, csa_tree_add_51_79_groupi_n_7626, csa_tree_add_51_79_groupi_n_7627, csa_tree_add_51_79_groupi_n_7628, csa_tree_add_51_79_groupi_n_7629, csa_tree_add_51_79_groupi_n_7630, csa_tree_add_51_79_groupi_n_7631;
  wire csa_tree_add_51_79_groupi_n_7632, csa_tree_add_51_79_groupi_n_7633, csa_tree_add_51_79_groupi_n_7634, csa_tree_add_51_79_groupi_n_7635, csa_tree_add_51_79_groupi_n_7636, csa_tree_add_51_79_groupi_n_7637, csa_tree_add_51_79_groupi_n_7638, csa_tree_add_51_79_groupi_n_7639;
  wire csa_tree_add_51_79_groupi_n_7640, csa_tree_add_51_79_groupi_n_7641, csa_tree_add_51_79_groupi_n_7642, csa_tree_add_51_79_groupi_n_7643, csa_tree_add_51_79_groupi_n_7644, csa_tree_add_51_79_groupi_n_7645, csa_tree_add_51_79_groupi_n_7646, csa_tree_add_51_79_groupi_n_7647;
  wire csa_tree_add_51_79_groupi_n_7648, csa_tree_add_51_79_groupi_n_7649, csa_tree_add_51_79_groupi_n_7650, csa_tree_add_51_79_groupi_n_7651, csa_tree_add_51_79_groupi_n_7652, csa_tree_add_51_79_groupi_n_7653, csa_tree_add_51_79_groupi_n_7654, csa_tree_add_51_79_groupi_n_7655;
  wire csa_tree_add_51_79_groupi_n_7656, csa_tree_add_51_79_groupi_n_7657, csa_tree_add_51_79_groupi_n_7658, csa_tree_add_51_79_groupi_n_7659, csa_tree_add_51_79_groupi_n_7660, csa_tree_add_51_79_groupi_n_7661, csa_tree_add_51_79_groupi_n_7662, csa_tree_add_51_79_groupi_n_7663;
  wire csa_tree_add_51_79_groupi_n_7664, csa_tree_add_51_79_groupi_n_7665, csa_tree_add_51_79_groupi_n_7666, csa_tree_add_51_79_groupi_n_7667, csa_tree_add_51_79_groupi_n_7668, csa_tree_add_51_79_groupi_n_7669, csa_tree_add_51_79_groupi_n_7670, csa_tree_add_51_79_groupi_n_7671;
  wire csa_tree_add_51_79_groupi_n_7672, csa_tree_add_51_79_groupi_n_7673, csa_tree_add_51_79_groupi_n_7674, csa_tree_add_51_79_groupi_n_7675, csa_tree_add_51_79_groupi_n_7676, csa_tree_add_51_79_groupi_n_7677, csa_tree_add_51_79_groupi_n_7678, csa_tree_add_51_79_groupi_n_7679;
  wire csa_tree_add_51_79_groupi_n_7680, csa_tree_add_51_79_groupi_n_7681, csa_tree_add_51_79_groupi_n_7682, csa_tree_add_51_79_groupi_n_7683, csa_tree_add_51_79_groupi_n_7684, csa_tree_add_51_79_groupi_n_7685, csa_tree_add_51_79_groupi_n_7686, csa_tree_add_51_79_groupi_n_7687;
  wire csa_tree_add_51_79_groupi_n_7688, csa_tree_add_51_79_groupi_n_7689, csa_tree_add_51_79_groupi_n_7690, csa_tree_add_51_79_groupi_n_7691, csa_tree_add_51_79_groupi_n_7692, csa_tree_add_51_79_groupi_n_7693, csa_tree_add_51_79_groupi_n_7694, csa_tree_add_51_79_groupi_n_7695;
  wire csa_tree_add_51_79_groupi_n_7696, csa_tree_add_51_79_groupi_n_7697, csa_tree_add_51_79_groupi_n_7698, csa_tree_add_51_79_groupi_n_7699, csa_tree_add_51_79_groupi_n_7700, csa_tree_add_51_79_groupi_n_7701, csa_tree_add_51_79_groupi_n_7702, csa_tree_add_51_79_groupi_n_7703;
  wire csa_tree_add_51_79_groupi_n_7704, csa_tree_add_51_79_groupi_n_7705, csa_tree_add_51_79_groupi_n_7706, csa_tree_add_51_79_groupi_n_7707, csa_tree_add_51_79_groupi_n_7708, csa_tree_add_51_79_groupi_n_7709, csa_tree_add_51_79_groupi_n_7710, csa_tree_add_51_79_groupi_n_7711;
  wire csa_tree_add_51_79_groupi_n_7712, csa_tree_add_51_79_groupi_n_7713, csa_tree_add_51_79_groupi_n_7714, csa_tree_add_51_79_groupi_n_7715, csa_tree_add_51_79_groupi_n_7716, csa_tree_add_51_79_groupi_n_7717, csa_tree_add_51_79_groupi_n_7718, csa_tree_add_51_79_groupi_n_7719;
  wire csa_tree_add_51_79_groupi_n_7720, csa_tree_add_51_79_groupi_n_7721, csa_tree_add_51_79_groupi_n_7722, csa_tree_add_51_79_groupi_n_7723, csa_tree_add_51_79_groupi_n_7724, csa_tree_add_51_79_groupi_n_7725, csa_tree_add_51_79_groupi_n_7726, csa_tree_add_51_79_groupi_n_7727;
  wire csa_tree_add_51_79_groupi_n_7728, csa_tree_add_51_79_groupi_n_7729, csa_tree_add_51_79_groupi_n_7730, csa_tree_add_51_79_groupi_n_7731, csa_tree_add_51_79_groupi_n_7732, csa_tree_add_51_79_groupi_n_7733, csa_tree_add_51_79_groupi_n_7734, csa_tree_add_51_79_groupi_n_7735;
  wire csa_tree_add_51_79_groupi_n_7736, csa_tree_add_51_79_groupi_n_7737, csa_tree_add_51_79_groupi_n_7738, csa_tree_add_51_79_groupi_n_7739, csa_tree_add_51_79_groupi_n_7740, csa_tree_add_51_79_groupi_n_7741, csa_tree_add_51_79_groupi_n_7742, csa_tree_add_51_79_groupi_n_7743;
  wire csa_tree_add_51_79_groupi_n_7744, csa_tree_add_51_79_groupi_n_7745, csa_tree_add_51_79_groupi_n_7746, csa_tree_add_51_79_groupi_n_7747, csa_tree_add_51_79_groupi_n_7748, csa_tree_add_51_79_groupi_n_7749, csa_tree_add_51_79_groupi_n_7750, csa_tree_add_51_79_groupi_n_7751;
  wire csa_tree_add_51_79_groupi_n_7752, csa_tree_add_51_79_groupi_n_7753, csa_tree_add_51_79_groupi_n_7754, csa_tree_add_51_79_groupi_n_7755, csa_tree_add_51_79_groupi_n_7756, csa_tree_add_51_79_groupi_n_7757, csa_tree_add_51_79_groupi_n_7758, csa_tree_add_51_79_groupi_n_7759;
  wire csa_tree_add_51_79_groupi_n_7760, csa_tree_add_51_79_groupi_n_7761, csa_tree_add_51_79_groupi_n_7762, csa_tree_add_51_79_groupi_n_7763, csa_tree_add_51_79_groupi_n_7764, csa_tree_add_51_79_groupi_n_7765, csa_tree_add_51_79_groupi_n_7766, csa_tree_add_51_79_groupi_n_7767;
  wire csa_tree_add_51_79_groupi_n_7768, csa_tree_add_51_79_groupi_n_7769, csa_tree_add_51_79_groupi_n_7770, csa_tree_add_51_79_groupi_n_7771, csa_tree_add_51_79_groupi_n_7772, csa_tree_add_51_79_groupi_n_7773, csa_tree_add_51_79_groupi_n_7774, csa_tree_add_51_79_groupi_n_7775;
  wire csa_tree_add_51_79_groupi_n_7776, csa_tree_add_51_79_groupi_n_7777, csa_tree_add_51_79_groupi_n_7778, csa_tree_add_51_79_groupi_n_7779, csa_tree_add_51_79_groupi_n_7780, csa_tree_add_51_79_groupi_n_7781, csa_tree_add_51_79_groupi_n_7782, csa_tree_add_51_79_groupi_n_7783;
  wire csa_tree_add_51_79_groupi_n_7784, csa_tree_add_51_79_groupi_n_7785, csa_tree_add_51_79_groupi_n_7786, csa_tree_add_51_79_groupi_n_7787, csa_tree_add_51_79_groupi_n_7788, csa_tree_add_51_79_groupi_n_7789, csa_tree_add_51_79_groupi_n_7790, csa_tree_add_51_79_groupi_n_7791;
  wire csa_tree_add_51_79_groupi_n_7792, csa_tree_add_51_79_groupi_n_7793, csa_tree_add_51_79_groupi_n_7794, csa_tree_add_51_79_groupi_n_7795, csa_tree_add_51_79_groupi_n_7796, csa_tree_add_51_79_groupi_n_7797, csa_tree_add_51_79_groupi_n_7798, csa_tree_add_51_79_groupi_n_7799;
  wire csa_tree_add_51_79_groupi_n_7800, csa_tree_add_51_79_groupi_n_7801, csa_tree_add_51_79_groupi_n_7802, csa_tree_add_51_79_groupi_n_7803, csa_tree_add_51_79_groupi_n_7804, csa_tree_add_51_79_groupi_n_7805, csa_tree_add_51_79_groupi_n_7806, csa_tree_add_51_79_groupi_n_7807;
  wire csa_tree_add_51_79_groupi_n_7808, csa_tree_add_51_79_groupi_n_7809, csa_tree_add_51_79_groupi_n_7810, csa_tree_add_51_79_groupi_n_7811, csa_tree_add_51_79_groupi_n_7812, csa_tree_add_51_79_groupi_n_7813, csa_tree_add_51_79_groupi_n_7814, csa_tree_add_51_79_groupi_n_7815;
  wire csa_tree_add_51_79_groupi_n_7816, csa_tree_add_51_79_groupi_n_7817, csa_tree_add_51_79_groupi_n_7818, csa_tree_add_51_79_groupi_n_7819, csa_tree_add_51_79_groupi_n_7820, csa_tree_add_51_79_groupi_n_7821, csa_tree_add_51_79_groupi_n_7822, csa_tree_add_51_79_groupi_n_7823;
  wire csa_tree_add_51_79_groupi_n_7824, csa_tree_add_51_79_groupi_n_7825, csa_tree_add_51_79_groupi_n_7826, csa_tree_add_51_79_groupi_n_7827, csa_tree_add_51_79_groupi_n_7828, csa_tree_add_51_79_groupi_n_7829, csa_tree_add_51_79_groupi_n_7830, csa_tree_add_51_79_groupi_n_7831;
  wire csa_tree_add_51_79_groupi_n_7832, csa_tree_add_51_79_groupi_n_7833, csa_tree_add_51_79_groupi_n_7834, csa_tree_add_51_79_groupi_n_7835, csa_tree_add_51_79_groupi_n_7836, csa_tree_add_51_79_groupi_n_7837, csa_tree_add_51_79_groupi_n_7838, csa_tree_add_51_79_groupi_n_7839;
  wire csa_tree_add_51_79_groupi_n_7840, csa_tree_add_51_79_groupi_n_7841, csa_tree_add_51_79_groupi_n_7842, csa_tree_add_51_79_groupi_n_7843, csa_tree_add_51_79_groupi_n_7844, csa_tree_add_51_79_groupi_n_7845, csa_tree_add_51_79_groupi_n_7846, csa_tree_add_51_79_groupi_n_7847;
  wire csa_tree_add_51_79_groupi_n_7848, csa_tree_add_51_79_groupi_n_7849, csa_tree_add_51_79_groupi_n_7850, csa_tree_add_51_79_groupi_n_7851, csa_tree_add_51_79_groupi_n_7852, csa_tree_add_51_79_groupi_n_7853, csa_tree_add_51_79_groupi_n_7854, csa_tree_add_51_79_groupi_n_7855;
  wire csa_tree_add_51_79_groupi_n_7856, csa_tree_add_51_79_groupi_n_7857, csa_tree_add_51_79_groupi_n_7858, csa_tree_add_51_79_groupi_n_7859, csa_tree_add_51_79_groupi_n_7860, csa_tree_add_51_79_groupi_n_7861, csa_tree_add_51_79_groupi_n_7862, csa_tree_add_51_79_groupi_n_7863;
  wire csa_tree_add_51_79_groupi_n_7864, csa_tree_add_51_79_groupi_n_7865, csa_tree_add_51_79_groupi_n_7866, csa_tree_add_51_79_groupi_n_7867, csa_tree_add_51_79_groupi_n_7868, csa_tree_add_51_79_groupi_n_7869, csa_tree_add_51_79_groupi_n_7870, csa_tree_add_51_79_groupi_n_7871;
  wire csa_tree_add_51_79_groupi_n_7872, csa_tree_add_51_79_groupi_n_7873, csa_tree_add_51_79_groupi_n_7874, csa_tree_add_51_79_groupi_n_7875, csa_tree_add_51_79_groupi_n_7876, csa_tree_add_51_79_groupi_n_7877, csa_tree_add_51_79_groupi_n_7878, csa_tree_add_51_79_groupi_n_7879;
  wire csa_tree_add_51_79_groupi_n_7880, csa_tree_add_51_79_groupi_n_7881, csa_tree_add_51_79_groupi_n_7882, csa_tree_add_51_79_groupi_n_7883, csa_tree_add_51_79_groupi_n_7884, csa_tree_add_51_79_groupi_n_7885, csa_tree_add_51_79_groupi_n_7886, csa_tree_add_51_79_groupi_n_7887;
  wire csa_tree_add_51_79_groupi_n_7888, csa_tree_add_51_79_groupi_n_7889, csa_tree_add_51_79_groupi_n_7890, csa_tree_add_51_79_groupi_n_7891, csa_tree_add_51_79_groupi_n_7892, csa_tree_add_51_79_groupi_n_7893, csa_tree_add_51_79_groupi_n_7894, csa_tree_add_51_79_groupi_n_7895;
  wire csa_tree_add_51_79_groupi_n_7896, csa_tree_add_51_79_groupi_n_7897, csa_tree_add_51_79_groupi_n_7898, csa_tree_add_51_79_groupi_n_7899, csa_tree_add_51_79_groupi_n_7900, csa_tree_add_51_79_groupi_n_7901, csa_tree_add_51_79_groupi_n_7902, csa_tree_add_51_79_groupi_n_7903;
  wire csa_tree_add_51_79_groupi_n_7904, csa_tree_add_51_79_groupi_n_7905, csa_tree_add_51_79_groupi_n_7906, csa_tree_add_51_79_groupi_n_7907, csa_tree_add_51_79_groupi_n_7908, csa_tree_add_51_79_groupi_n_7909, csa_tree_add_51_79_groupi_n_7910, csa_tree_add_51_79_groupi_n_7911;
  wire csa_tree_add_51_79_groupi_n_7912, csa_tree_add_51_79_groupi_n_7913, csa_tree_add_51_79_groupi_n_7914, csa_tree_add_51_79_groupi_n_7915, csa_tree_add_51_79_groupi_n_7916, csa_tree_add_51_79_groupi_n_7917, csa_tree_add_51_79_groupi_n_7918, csa_tree_add_51_79_groupi_n_7919;
  wire csa_tree_add_51_79_groupi_n_7920, csa_tree_add_51_79_groupi_n_7921, csa_tree_add_51_79_groupi_n_7922, csa_tree_add_51_79_groupi_n_7923, csa_tree_add_51_79_groupi_n_7924, csa_tree_add_51_79_groupi_n_7925, csa_tree_add_51_79_groupi_n_7926, csa_tree_add_51_79_groupi_n_7927;
  wire csa_tree_add_51_79_groupi_n_7928, csa_tree_add_51_79_groupi_n_7929, csa_tree_add_51_79_groupi_n_7930, csa_tree_add_51_79_groupi_n_7931, csa_tree_add_51_79_groupi_n_7932, csa_tree_add_51_79_groupi_n_7933, csa_tree_add_51_79_groupi_n_7934, csa_tree_add_51_79_groupi_n_7935;
  wire csa_tree_add_51_79_groupi_n_7936, csa_tree_add_51_79_groupi_n_7937, csa_tree_add_51_79_groupi_n_7938, csa_tree_add_51_79_groupi_n_7939, csa_tree_add_51_79_groupi_n_7940, csa_tree_add_51_79_groupi_n_7941, csa_tree_add_51_79_groupi_n_7942, csa_tree_add_51_79_groupi_n_7943;
  wire csa_tree_add_51_79_groupi_n_7944, csa_tree_add_51_79_groupi_n_7945, csa_tree_add_51_79_groupi_n_7946, csa_tree_add_51_79_groupi_n_7947, csa_tree_add_51_79_groupi_n_7948, csa_tree_add_51_79_groupi_n_7949, csa_tree_add_51_79_groupi_n_7950, csa_tree_add_51_79_groupi_n_7951;
  wire csa_tree_add_51_79_groupi_n_7952, csa_tree_add_51_79_groupi_n_7953, csa_tree_add_51_79_groupi_n_7954, csa_tree_add_51_79_groupi_n_7955, csa_tree_add_51_79_groupi_n_7956, csa_tree_add_51_79_groupi_n_7957, csa_tree_add_51_79_groupi_n_7958, csa_tree_add_51_79_groupi_n_7959;
  wire csa_tree_add_51_79_groupi_n_7960, csa_tree_add_51_79_groupi_n_7961, csa_tree_add_51_79_groupi_n_7962, csa_tree_add_51_79_groupi_n_7963, csa_tree_add_51_79_groupi_n_7964, csa_tree_add_51_79_groupi_n_7965, csa_tree_add_51_79_groupi_n_7966, csa_tree_add_51_79_groupi_n_7967;
  wire csa_tree_add_51_79_groupi_n_7968, csa_tree_add_51_79_groupi_n_7969, csa_tree_add_51_79_groupi_n_7970, csa_tree_add_51_79_groupi_n_7971, csa_tree_add_51_79_groupi_n_7972, csa_tree_add_51_79_groupi_n_7973, csa_tree_add_51_79_groupi_n_7974, csa_tree_add_51_79_groupi_n_7975;
  wire csa_tree_add_51_79_groupi_n_7976, csa_tree_add_51_79_groupi_n_7977, csa_tree_add_51_79_groupi_n_7978, csa_tree_add_51_79_groupi_n_7979, csa_tree_add_51_79_groupi_n_7980, csa_tree_add_51_79_groupi_n_7981, csa_tree_add_51_79_groupi_n_7982, csa_tree_add_51_79_groupi_n_7983;
  wire csa_tree_add_51_79_groupi_n_7984, csa_tree_add_51_79_groupi_n_7985, csa_tree_add_51_79_groupi_n_7986, csa_tree_add_51_79_groupi_n_7987, csa_tree_add_51_79_groupi_n_7988, csa_tree_add_51_79_groupi_n_7989, csa_tree_add_51_79_groupi_n_7990, csa_tree_add_51_79_groupi_n_7991;
  wire csa_tree_add_51_79_groupi_n_7992, csa_tree_add_51_79_groupi_n_7993, csa_tree_add_51_79_groupi_n_7994, csa_tree_add_51_79_groupi_n_7995, csa_tree_add_51_79_groupi_n_7996, csa_tree_add_51_79_groupi_n_7997, csa_tree_add_51_79_groupi_n_7998, csa_tree_add_51_79_groupi_n_7999;
  wire csa_tree_add_51_79_groupi_n_8000, csa_tree_add_51_79_groupi_n_8001, csa_tree_add_51_79_groupi_n_8002, csa_tree_add_51_79_groupi_n_8003, csa_tree_add_51_79_groupi_n_8004, csa_tree_add_51_79_groupi_n_8005, csa_tree_add_51_79_groupi_n_8006, csa_tree_add_51_79_groupi_n_8007;
  wire csa_tree_add_51_79_groupi_n_8008, csa_tree_add_51_79_groupi_n_8009, csa_tree_add_51_79_groupi_n_8010, csa_tree_add_51_79_groupi_n_8011, csa_tree_add_51_79_groupi_n_8012, csa_tree_add_51_79_groupi_n_8013, csa_tree_add_51_79_groupi_n_8014, csa_tree_add_51_79_groupi_n_8015;
  wire csa_tree_add_51_79_groupi_n_8016, csa_tree_add_51_79_groupi_n_8017, csa_tree_add_51_79_groupi_n_8018, csa_tree_add_51_79_groupi_n_8019, csa_tree_add_51_79_groupi_n_8020, csa_tree_add_51_79_groupi_n_8021, csa_tree_add_51_79_groupi_n_8022, csa_tree_add_51_79_groupi_n_8023;
  wire csa_tree_add_51_79_groupi_n_8024, csa_tree_add_51_79_groupi_n_8025, csa_tree_add_51_79_groupi_n_8026, csa_tree_add_51_79_groupi_n_8027, csa_tree_add_51_79_groupi_n_8028, csa_tree_add_51_79_groupi_n_8029, csa_tree_add_51_79_groupi_n_8030, csa_tree_add_51_79_groupi_n_8031;
  wire csa_tree_add_51_79_groupi_n_8032, csa_tree_add_51_79_groupi_n_8033, csa_tree_add_51_79_groupi_n_8034, csa_tree_add_51_79_groupi_n_8035, csa_tree_add_51_79_groupi_n_8036, csa_tree_add_51_79_groupi_n_8037, csa_tree_add_51_79_groupi_n_8038, csa_tree_add_51_79_groupi_n_8039;
  wire csa_tree_add_51_79_groupi_n_8040, csa_tree_add_51_79_groupi_n_8041, csa_tree_add_51_79_groupi_n_8042, csa_tree_add_51_79_groupi_n_8043, csa_tree_add_51_79_groupi_n_8044, csa_tree_add_51_79_groupi_n_8045, csa_tree_add_51_79_groupi_n_8046, csa_tree_add_51_79_groupi_n_8047;
  wire csa_tree_add_51_79_groupi_n_8048, csa_tree_add_51_79_groupi_n_8049, csa_tree_add_51_79_groupi_n_8050, csa_tree_add_51_79_groupi_n_8051, csa_tree_add_51_79_groupi_n_8052, csa_tree_add_51_79_groupi_n_8053, csa_tree_add_51_79_groupi_n_8054, csa_tree_add_51_79_groupi_n_8055;
  wire csa_tree_add_51_79_groupi_n_8056, csa_tree_add_51_79_groupi_n_8057, csa_tree_add_51_79_groupi_n_8058, csa_tree_add_51_79_groupi_n_8059, csa_tree_add_51_79_groupi_n_8060, csa_tree_add_51_79_groupi_n_8061, csa_tree_add_51_79_groupi_n_8062, csa_tree_add_51_79_groupi_n_8063;
  wire csa_tree_add_51_79_groupi_n_8064, csa_tree_add_51_79_groupi_n_8065, csa_tree_add_51_79_groupi_n_8066, csa_tree_add_51_79_groupi_n_8067, csa_tree_add_51_79_groupi_n_8068, csa_tree_add_51_79_groupi_n_8069, csa_tree_add_51_79_groupi_n_8070, csa_tree_add_51_79_groupi_n_8071;
  wire csa_tree_add_51_79_groupi_n_8072, csa_tree_add_51_79_groupi_n_8073, csa_tree_add_51_79_groupi_n_8074, csa_tree_add_51_79_groupi_n_8075, csa_tree_add_51_79_groupi_n_8076, csa_tree_add_51_79_groupi_n_8077, csa_tree_add_51_79_groupi_n_8078, csa_tree_add_51_79_groupi_n_8079;
  wire csa_tree_add_51_79_groupi_n_8080, csa_tree_add_51_79_groupi_n_8081, csa_tree_add_51_79_groupi_n_8082, csa_tree_add_51_79_groupi_n_8083, csa_tree_add_51_79_groupi_n_8084, csa_tree_add_51_79_groupi_n_8085, csa_tree_add_51_79_groupi_n_8086, csa_tree_add_51_79_groupi_n_8087;
  wire csa_tree_add_51_79_groupi_n_8088, csa_tree_add_51_79_groupi_n_8089, csa_tree_add_51_79_groupi_n_8090, csa_tree_add_51_79_groupi_n_8091, csa_tree_add_51_79_groupi_n_8092, csa_tree_add_51_79_groupi_n_8093, csa_tree_add_51_79_groupi_n_8094, csa_tree_add_51_79_groupi_n_8095;
  wire csa_tree_add_51_79_groupi_n_8096, csa_tree_add_51_79_groupi_n_8097, csa_tree_add_51_79_groupi_n_8098, csa_tree_add_51_79_groupi_n_8099, csa_tree_add_51_79_groupi_n_8100, csa_tree_add_51_79_groupi_n_8101, csa_tree_add_51_79_groupi_n_8102, csa_tree_add_51_79_groupi_n_8103;
  wire csa_tree_add_51_79_groupi_n_8104, csa_tree_add_51_79_groupi_n_8105, csa_tree_add_51_79_groupi_n_8106, csa_tree_add_51_79_groupi_n_8107, csa_tree_add_51_79_groupi_n_8108, csa_tree_add_51_79_groupi_n_8109, csa_tree_add_51_79_groupi_n_8110, csa_tree_add_51_79_groupi_n_8111;
  wire csa_tree_add_51_79_groupi_n_8112, csa_tree_add_51_79_groupi_n_8113, csa_tree_add_51_79_groupi_n_8114, csa_tree_add_51_79_groupi_n_8115, csa_tree_add_51_79_groupi_n_8116, csa_tree_add_51_79_groupi_n_8117, csa_tree_add_51_79_groupi_n_8118, csa_tree_add_51_79_groupi_n_8119;
  wire csa_tree_add_51_79_groupi_n_8120, csa_tree_add_51_79_groupi_n_8121, csa_tree_add_51_79_groupi_n_8122, csa_tree_add_51_79_groupi_n_8123, csa_tree_add_51_79_groupi_n_8124, csa_tree_add_51_79_groupi_n_8125, csa_tree_add_51_79_groupi_n_8126, csa_tree_add_51_79_groupi_n_8127;
  wire csa_tree_add_51_79_groupi_n_8128, csa_tree_add_51_79_groupi_n_8129, csa_tree_add_51_79_groupi_n_8130, csa_tree_add_51_79_groupi_n_8131, csa_tree_add_51_79_groupi_n_8132, csa_tree_add_51_79_groupi_n_8133, csa_tree_add_51_79_groupi_n_8134, csa_tree_add_51_79_groupi_n_8135;
  wire csa_tree_add_51_79_groupi_n_8136, csa_tree_add_51_79_groupi_n_8137, csa_tree_add_51_79_groupi_n_8138, csa_tree_add_51_79_groupi_n_8140, csa_tree_add_51_79_groupi_n_8141, csa_tree_add_51_79_groupi_n_8142, csa_tree_add_51_79_groupi_n_8143, csa_tree_add_51_79_groupi_n_8144;
  wire csa_tree_add_51_79_groupi_n_8145, csa_tree_add_51_79_groupi_n_8146, csa_tree_add_51_79_groupi_n_8147, csa_tree_add_51_79_groupi_n_8148, csa_tree_add_51_79_groupi_n_8149, csa_tree_add_51_79_groupi_n_8150, csa_tree_add_51_79_groupi_n_8151, csa_tree_add_51_79_groupi_n_8152;
  wire csa_tree_add_51_79_groupi_n_8153, csa_tree_add_51_79_groupi_n_8154, csa_tree_add_51_79_groupi_n_8155, csa_tree_add_51_79_groupi_n_8156, csa_tree_add_51_79_groupi_n_8157, csa_tree_add_51_79_groupi_n_8158, csa_tree_add_51_79_groupi_n_8159, csa_tree_add_51_79_groupi_n_8160;
  wire csa_tree_add_51_79_groupi_n_8161, csa_tree_add_51_79_groupi_n_8162, csa_tree_add_51_79_groupi_n_8163, csa_tree_add_51_79_groupi_n_8164, csa_tree_add_51_79_groupi_n_8165, csa_tree_add_51_79_groupi_n_8166, csa_tree_add_51_79_groupi_n_8167, csa_tree_add_51_79_groupi_n_8168;
  wire csa_tree_add_51_79_groupi_n_8169, csa_tree_add_51_79_groupi_n_8170, csa_tree_add_51_79_groupi_n_8171, csa_tree_add_51_79_groupi_n_8172, csa_tree_add_51_79_groupi_n_8173, csa_tree_add_51_79_groupi_n_8174, csa_tree_add_51_79_groupi_n_8175, csa_tree_add_51_79_groupi_n_8176;
  wire csa_tree_add_51_79_groupi_n_8177, csa_tree_add_51_79_groupi_n_8178, csa_tree_add_51_79_groupi_n_8179, csa_tree_add_51_79_groupi_n_8180, csa_tree_add_51_79_groupi_n_8181, csa_tree_add_51_79_groupi_n_8182, csa_tree_add_51_79_groupi_n_8183, csa_tree_add_51_79_groupi_n_8184;
  wire csa_tree_add_51_79_groupi_n_8185, csa_tree_add_51_79_groupi_n_8186, csa_tree_add_51_79_groupi_n_8187, csa_tree_add_51_79_groupi_n_8188, csa_tree_add_51_79_groupi_n_8189, csa_tree_add_51_79_groupi_n_8190, csa_tree_add_51_79_groupi_n_8191, csa_tree_add_51_79_groupi_n_8192;
  wire csa_tree_add_51_79_groupi_n_8193, csa_tree_add_51_79_groupi_n_8194, csa_tree_add_51_79_groupi_n_8195, csa_tree_add_51_79_groupi_n_8196, csa_tree_add_51_79_groupi_n_8197, csa_tree_add_51_79_groupi_n_8198, csa_tree_add_51_79_groupi_n_8199, csa_tree_add_51_79_groupi_n_8200;
  wire csa_tree_add_51_79_groupi_n_8201, csa_tree_add_51_79_groupi_n_8202, csa_tree_add_51_79_groupi_n_8203, csa_tree_add_51_79_groupi_n_8204, csa_tree_add_51_79_groupi_n_8205, csa_tree_add_51_79_groupi_n_8206, csa_tree_add_51_79_groupi_n_8207, csa_tree_add_51_79_groupi_n_8208;
  wire csa_tree_add_51_79_groupi_n_8209, csa_tree_add_51_79_groupi_n_8210, csa_tree_add_51_79_groupi_n_8211, csa_tree_add_51_79_groupi_n_8212, csa_tree_add_51_79_groupi_n_8213, csa_tree_add_51_79_groupi_n_8214, csa_tree_add_51_79_groupi_n_8215, csa_tree_add_51_79_groupi_n_8216;
  wire csa_tree_add_51_79_groupi_n_8217, csa_tree_add_51_79_groupi_n_8218, csa_tree_add_51_79_groupi_n_8219, csa_tree_add_51_79_groupi_n_8220, csa_tree_add_51_79_groupi_n_8221, csa_tree_add_51_79_groupi_n_8222, csa_tree_add_51_79_groupi_n_8223, csa_tree_add_51_79_groupi_n_8224;
  wire csa_tree_add_51_79_groupi_n_8225, csa_tree_add_51_79_groupi_n_8226, csa_tree_add_51_79_groupi_n_8227, csa_tree_add_51_79_groupi_n_8228, csa_tree_add_51_79_groupi_n_8229, csa_tree_add_51_79_groupi_n_8230, csa_tree_add_51_79_groupi_n_8231, csa_tree_add_51_79_groupi_n_8232;
  wire csa_tree_add_51_79_groupi_n_8233, csa_tree_add_51_79_groupi_n_8234, csa_tree_add_51_79_groupi_n_8235, csa_tree_add_51_79_groupi_n_8236, csa_tree_add_51_79_groupi_n_8237, csa_tree_add_51_79_groupi_n_8238, csa_tree_add_51_79_groupi_n_8239, csa_tree_add_51_79_groupi_n_8240;
  wire csa_tree_add_51_79_groupi_n_8241, csa_tree_add_51_79_groupi_n_8242, csa_tree_add_51_79_groupi_n_8243, csa_tree_add_51_79_groupi_n_8244, csa_tree_add_51_79_groupi_n_8245, csa_tree_add_51_79_groupi_n_8246, csa_tree_add_51_79_groupi_n_8247, csa_tree_add_51_79_groupi_n_8248;
  wire csa_tree_add_51_79_groupi_n_8249, csa_tree_add_51_79_groupi_n_8250, csa_tree_add_51_79_groupi_n_8251, csa_tree_add_51_79_groupi_n_8252, csa_tree_add_51_79_groupi_n_8253, csa_tree_add_51_79_groupi_n_8254, csa_tree_add_51_79_groupi_n_8255, csa_tree_add_51_79_groupi_n_8256;
  wire csa_tree_add_51_79_groupi_n_8257, csa_tree_add_51_79_groupi_n_8258, csa_tree_add_51_79_groupi_n_8259, csa_tree_add_51_79_groupi_n_8260, csa_tree_add_51_79_groupi_n_8261, csa_tree_add_51_79_groupi_n_8262, csa_tree_add_51_79_groupi_n_8263, csa_tree_add_51_79_groupi_n_8264;
  wire csa_tree_add_51_79_groupi_n_8265, csa_tree_add_51_79_groupi_n_8266, csa_tree_add_51_79_groupi_n_8267, csa_tree_add_51_79_groupi_n_8268, csa_tree_add_51_79_groupi_n_8269, csa_tree_add_51_79_groupi_n_8270, csa_tree_add_51_79_groupi_n_8271, csa_tree_add_51_79_groupi_n_8272;
  wire csa_tree_add_51_79_groupi_n_8273, csa_tree_add_51_79_groupi_n_8274, csa_tree_add_51_79_groupi_n_8275, csa_tree_add_51_79_groupi_n_8276, csa_tree_add_51_79_groupi_n_8277, csa_tree_add_51_79_groupi_n_8278, csa_tree_add_51_79_groupi_n_8279, csa_tree_add_51_79_groupi_n_8280;
  wire csa_tree_add_51_79_groupi_n_8281, csa_tree_add_51_79_groupi_n_8282, csa_tree_add_51_79_groupi_n_8283, csa_tree_add_51_79_groupi_n_8284, csa_tree_add_51_79_groupi_n_8285, csa_tree_add_51_79_groupi_n_8286, csa_tree_add_51_79_groupi_n_8287, csa_tree_add_51_79_groupi_n_8288;
  wire csa_tree_add_51_79_groupi_n_8289, csa_tree_add_51_79_groupi_n_8290, csa_tree_add_51_79_groupi_n_8291, csa_tree_add_51_79_groupi_n_8292, csa_tree_add_51_79_groupi_n_8293, csa_tree_add_51_79_groupi_n_8294, csa_tree_add_51_79_groupi_n_8295, csa_tree_add_51_79_groupi_n_8296;
  wire csa_tree_add_51_79_groupi_n_8297, csa_tree_add_51_79_groupi_n_8298, csa_tree_add_51_79_groupi_n_8299, csa_tree_add_51_79_groupi_n_8300, csa_tree_add_51_79_groupi_n_8301, csa_tree_add_51_79_groupi_n_8302, csa_tree_add_51_79_groupi_n_8303, csa_tree_add_51_79_groupi_n_8304;
  wire csa_tree_add_51_79_groupi_n_8305, csa_tree_add_51_79_groupi_n_8306, csa_tree_add_51_79_groupi_n_8307, csa_tree_add_51_79_groupi_n_8308, csa_tree_add_51_79_groupi_n_8309, csa_tree_add_51_79_groupi_n_8310, csa_tree_add_51_79_groupi_n_8311, csa_tree_add_51_79_groupi_n_8312;
  wire csa_tree_add_51_79_groupi_n_8313, csa_tree_add_51_79_groupi_n_8314, csa_tree_add_51_79_groupi_n_8315, csa_tree_add_51_79_groupi_n_8316, csa_tree_add_51_79_groupi_n_8317, csa_tree_add_51_79_groupi_n_8318, csa_tree_add_51_79_groupi_n_8319, csa_tree_add_51_79_groupi_n_8320;
  wire csa_tree_add_51_79_groupi_n_8321, csa_tree_add_51_79_groupi_n_8322, csa_tree_add_51_79_groupi_n_8323, csa_tree_add_51_79_groupi_n_8324, csa_tree_add_51_79_groupi_n_8325, csa_tree_add_51_79_groupi_n_8326, csa_tree_add_51_79_groupi_n_8327, csa_tree_add_51_79_groupi_n_8328;
  wire csa_tree_add_51_79_groupi_n_8329, csa_tree_add_51_79_groupi_n_8330, csa_tree_add_51_79_groupi_n_8331, csa_tree_add_51_79_groupi_n_8332, csa_tree_add_51_79_groupi_n_8333, csa_tree_add_51_79_groupi_n_8334, csa_tree_add_51_79_groupi_n_8335, csa_tree_add_51_79_groupi_n_8336;
  wire csa_tree_add_51_79_groupi_n_8337, csa_tree_add_51_79_groupi_n_8338, csa_tree_add_51_79_groupi_n_8339, csa_tree_add_51_79_groupi_n_8340, csa_tree_add_51_79_groupi_n_8341, csa_tree_add_51_79_groupi_n_8342, csa_tree_add_51_79_groupi_n_8343, csa_tree_add_51_79_groupi_n_8344;
  wire csa_tree_add_51_79_groupi_n_8345, csa_tree_add_51_79_groupi_n_8346, csa_tree_add_51_79_groupi_n_8347, csa_tree_add_51_79_groupi_n_8348, csa_tree_add_51_79_groupi_n_8349, csa_tree_add_51_79_groupi_n_8350, csa_tree_add_51_79_groupi_n_8351, csa_tree_add_51_79_groupi_n_8352;
  wire csa_tree_add_51_79_groupi_n_8353, csa_tree_add_51_79_groupi_n_8354, csa_tree_add_51_79_groupi_n_8355, csa_tree_add_51_79_groupi_n_8356, csa_tree_add_51_79_groupi_n_8357, csa_tree_add_51_79_groupi_n_8358, csa_tree_add_51_79_groupi_n_8359, csa_tree_add_51_79_groupi_n_8360;
  wire csa_tree_add_51_79_groupi_n_8361, csa_tree_add_51_79_groupi_n_8362, csa_tree_add_51_79_groupi_n_8363, csa_tree_add_51_79_groupi_n_8364, csa_tree_add_51_79_groupi_n_8365, csa_tree_add_51_79_groupi_n_8366, csa_tree_add_51_79_groupi_n_8367, csa_tree_add_51_79_groupi_n_8368;
  wire csa_tree_add_51_79_groupi_n_8369, csa_tree_add_51_79_groupi_n_8370, csa_tree_add_51_79_groupi_n_8371, csa_tree_add_51_79_groupi_n_8372, csa_tree_add_51_79_groupi_n_8373, csa_tree_add_51_79_groupi_n_8374, csa_tree_add_51_79_groupi_n_8375, csa_tree_add_51_79_groupi_n_8376;
  wire csa_tree_add_51_79_groupi_n_8377, csa_tree_add_51_79_groupi_n_8378, csa_tree_add_51_79_groupi_n_8379, csa_tree_add_51_79_groupi_n_8380, csa_tree_add_51_79_groupi_n_8381, csa_tree_add_51_79_groupi_n_8382, csa_tree_add_51_79_groupi_n_8383, csa_tree_add_51_79_groupi_n_8384;
  wire csa_tree_add_51_79_groupi_n_8385, csa_tree_add_51_79_groupi_n_8386, csa_tree_add_51_79_groupi_n_8387, csa_tree_add_51_79_groupi_n_8388, csa_tree_add_51_79_groupi_n_8389, csa_tree_add_51_79_groupi_n_8390, csa_tree_add_51_79_groupi_n_8391, csa_tree_add_51_79_groupi_n_8392;
  wire csa_tree_add_51_79_groupi_n_8393, csa_tree_add_51_79_groupi_n_8394, csa_tree_add_51_79_groupi_n_8395, csa_tree_add_51_79_groupi_n_8396, csa_tree_add_51_79_groupi_n_8397, csa_tree_add_51_79_groupi_n_8398, csa_tree_add_51_79_groupi_n_8399, csa_tree_add_51_79_groupi_n_8400;
  wire csa_tree_add_51_79_groupi_n_8401, csa_tree_add_51_79_groupi_n_8402, csa_tree_add_51_79_groupi_n_8403, csa_tree_add_51_79_groupi_n_8404, csa_tree_add_51_79_groupi_n_8405, csa_tree_add_51_79_groupi_n_8406, csa_tree_add_51_79_groupi_n_8407, csa_tree_add_51_79_groupi_n_8408;
  wire csa_tree_add_51_79_groupi_n_8409, csa_tree_add_51_79_groupi_n_8410, csa_tree_add_51_79_groupi_n_8411, csa_tree_add_51_79_groupi_n_8412, csa_tree_add_51_79_groupi_n_8413, csa_tree_add_51_79_groupi_n_8414, csa_tree_add_51_79_groupi_n_8415, csa_tree_add_51_79_groupi_n_8416;
  wire csa_tree_add_51_79_groupi_n_8417, csa_tree_add_51_79_groupi_n_8418, csa_tree_add_51_79_groupi_n_8419, csa_tree_add_51_79_groupi_n_8420, csa_tree_add_51_79_groupi_n_8421, csa_tree_add_51_79_groupi_n_8422, csa_tree_add_51_79_groupi_n_8423, csa_tree_add_51_79_groupi_n_8424;
  wire csa_tree_add_51_79_groupi_n_8425, csa_tree_add_51_79_groupi_n_8426, csa_tree_add_51_79_groupi_n_8427, csa_tree_add_51_79_groupi_n_8428, csa_tree_add_51_79_groupi_n_8429, csa_tree_add_51_79_groupi_n_8430, csa_tree_add_51_79_groupi_n_8431, csa_tree_add_51_79_groupi_n_8432;
  wire csa_tree_add_51_79_groupi_n_8433, csa_tree_add_51_79_groupi_n_8434, csa_tree_add_51_79_groupi_n_8435, csa_tree_add_51_79_groupi_n_8436, csa_tree_add_51_79_groupi_n_8437, csa_tree_add_51_79_groupi_n_8438, csa_tree_add_51_79_groupi_n_8439, csa_tree_add_51_79_groupi_n_8440;
  wire csa_tree_add_51_79_groupi_n_8441, csa_tree_add_51_79_groupi_n_8442, csa_tree_add_51_79_groupi_n_8443, csa_tree_add_51_79_groupi_n_8444, csa_tree_add_51_79_groupi_n_8445, csa_tree_add_51_79_groupi_n_8446, csa_tree_add_51_79_groupi_n_8447, csa_tree_add_51_79_groupi_n_8448;
  wire csa_tree_add_51_79_groupi_n_8449, csa_tree_add_51_79_groupi_n_8450, csa_tree_add_51_79_groupi_n_8451, csa_tree_add_51_79_groupi_n_8452, csa_tree_add_51_79_groupi_n_8453, csa_tree_add_51_79_groupi_n_8454, csa_tree_add_51_79_groupi_n_8455, csa_tree_add_51_79_groupi_n_8456;
  wire csa_tree_add_51_79_groupi_n_8457, csa_tree_add_51_79_groupi_n_8458, csa_tree_add_51_79_groupi_n_8459, csa_tree_add_51_79_groupi_n_8460, csa_tree_add_51_79_groupi_n_8461, csa_tree_add_51_79_groupi_n_8462, csa_tree_add_51_79_groupi_n_8463, csa_tree_add_51_79_groupi_n_8464;
  wire csa_tree_add_51_79_groupi_n_8465, csa_tree_add_51_79_groupi_n_8466, csa_tree_add_51_79_groupi_n_8467, csa_tree_add_51_79_groupi_n_8468, csa_tree_add_51_79_groupi_n_8469, csa_tree_add_51_79_groupi_n_8470, csa_tree_add_51_79_groupi_n_8471, csa_tree_add_51_79_groupi_n_8472;
  wire csa_tree_add_51_79_groupi_n_8473, csa_tree_add_51_79_groupi_n_8474, csa_tree_add_51_79_groupi_n_8475, csa_tree_add_51_79_groupi_n_8476, csa_tree_add_51_79_groupi_n_8477, csa_tree_add_51_79_groupi_n_8478, csa_tree_add_51_79_groupi_n_8479, csa_tree_add_51_79_groupi_n_8480;
  wire csa_tree_add_51_79_groupi_n_8481, csa_tree_add_51_79_groupi_n_8482, csa_tree_add_51_79_groupi_n_8483, csa_tree_add_51_79_groupi_n_8484, csa_tree_add_51_79_groupi_n_8485, csa_tree_add_51_79_groupi_n_8486, csa_tree_add_51_79_groupi_n_8487, csa_tree_add_51_79_groupi_n_8488;
  wire csa_tree_add_51_79_groupi_n_8489, csa_tree_add_51_79_groupi_n_8490, csa_tree_add_51_79_groupi_n_8491, csa_tree_add_51_79_groupi_n_8492, csa_tree_add_51_79_groupi_n_8493, csa_tree_add_51_79_groupi_n_8494, csa_tree_add_51_79_groupi_n_8495, csa_tree_add_51_79_groupi_n_8496;
  wire csa_tree_add_51_79_groupi_n_8497, csa_tree_add_51_79_groupi_n_8498, csa_tree_add_51_79_groupi_n_8499, csa_tree_add_51_79_groupi_n_8500, csa_tree_add_51_79_groupi_n_8501, csa_tree_add_51_79_groupi_n_8502, csa_tree_add_51_79_groupi_n_8503, csa_tree_add_51_79_groupi_n_8504;
  wire csa_tree_add_51_79_groupi_n_8505, csa_tree_add_51_79_groupi_n_8506, csa_tree_add_51_79_groupi_n_8507, csa_tree_add_51_79_groupi_n_8508, csa_tree_add_51_79_groupi_n_8509, csa_tree_add_51_79_groupi_n_8510, csa_tree_add_51_79_groupi_n_8511, csa_tree_add_51_79_groupi_n_8512;
  wire csa_tree_add_51_79_groupi_n_8513, csa_tree_add_51_79_groupi_n_8514, csa_tree_add_51_79_groupi_n_8515, csa_tree_add_51_79_groupi_n_8516, csa_tree_add_51_79_groupi_n_8517, csa_tree_add_51_79_groupi_n_8518, csa_tree_add_51_79_groupi_n_8519, csa_tree_add_51_79_groupi_n_8520;
  wire csa_tree_add_51_79_groupi_n_8521, csa_tree_add_51_79_groupi_n_8522, csa_tree_add_51_79_groupi_n_8523, csa_tree_add_51_79_groupi_n_8524, csa_tree_add_51_79_groupi_n_8525, csa_tree_add_51_79_groupi_n_8526, csa_tree_add_51_79_groupi_n_8527, csa_tree_add_51_79_groupi_n_8528;
  wire csa_tree_add_51_79_groupi_n_8529, csa_tree_add_51_79_groupi_n_8530, csa_tree_add_51_79_groupi_n_8531, csa_tree_add_51_79_groupi_n_8532, csa_tree_add_51_79_groupi_n_8533, csa_tree_add_51_79_groupi_n_8534, csa_tree_add_51_79_groupi_n_8535, csa_tree_add_51_79_groupi_n_8536;
  wire csa_tree_add_51_79_groupi_n_8537, csa_tree_add_51_79_groupi_n_8538, csa_tree_add_51_79_groupi_n_8539, csa_tree_add_51_79_groupi_n_8540, csa_tree_add_51_79_groupi_n_8541, csa_tree_add_51_79_groupi_n_8542, csa_tree_add_51_79_groupi_n_8543, csa_tree_add_51_79_groupi_n_8544;
  wire csa_tree_add_51_79_groupi_n_8545, csa_tree_add_51_79_groupi_n_8546, csa_tree_add_51_79_groupi_n_8547, csa_tree_add_51_79_groupi_n_8548, csa_tree_add_51_79_groupi_n_8549, csa_tree_add_51_79_groupi_n_8550, csa_tree_add_51_79_groupi_n_8551, csa_tree_add_51_79_groupi_n_8552;
  wire csa_tree_add_51_79_groupi_n_8553, csa_tree_add_51_79_groupi_n_8554, csa_tree_add_51_79_groupi_n_8555, csa_tree_add_51_79_groupi_n_8556, csa_tree_add_51_79_groupi_n_8557, csa_tree_add_51_79_groupi_n_8558, csa_tree_add_51_79_groupi_n_8559, csa_tree_add_51_79_groupi_n_8560;
  wire csa_tree_add_51_79_groupi_n_8561, csa_tree_add_51_79_groupi_n_8562, csa_tree_add_51_79_groupi_n_8563, csa_tree_add_51_79_groupi_n_8564, csa_tree_add_51_79_groupi_n_8565, csa_tree_add_51_79_groupi_n_8566, csa_tree_add_51_79_groupi_n_8567, csa_tree_add_51_79_groupi_n_8568;
  wire csa_tree_add_51_79_groupi_n_8569, csa_tree_add_51_79_groupi_n_8570, csa_tree_add_51_79_groupi_n_8571, csa_tree_add_51_79_groupi_n_8572, csa_tree_add_51_79_groupi_n_8573, csa_tree_add_51_79_groupi_n_8574, csa_tree_add_51_79_groupi_n_8575, csa_tree_add_51_79_groupi_n_8576;
  wire csa_tree_add_51_79_groupi_n_8577, csa_tree_add_51_79_groupi_n_8578, csa_tree_add_51_79_groupi_n_8579, csa_tree_add_51_79_groupi_n_8580, csa_tree_add_51_79_groupi_n_8581, csa_tree_add_51_79_groupi_n_8582, csa_tree_add_51_79_groupi_n_8583, csa_tree_add_51_79_groupi_n_8584;
  wire csa_tree_add_51_79_groupi_n_8585, csa_tree_add_51_79_groupi_n_8586, csa_tree_add_51_79_groupi_n_8587, csa_tree_add_51_79_groupi_n_8588, csa_tree_add_51_79_groupi_n_8589, csa_tree_add_51_79_groupi_n_8590, csa_tree_add_51_79_groupi_n_8591, csa_tree_add_51_79_groupi_n_8592;
  wire csa_tree_add_51_79_groupi_n_8593, csa_tree_add_51_79_groupi_n_8594, csa_tree_add_51_79_groupi_n_8595, csa_tree_add_51_79_groupi_n_8596, csa_tree_add_51_79_groupi_n_8597, csa_tree_add_51_79_groupi_n_8598, csa_tree_add_51_79_groupi_n_8599, csa_tree_add_51_79_groupi_n_8600;
  wire csa_tree_add_51_79_groupi_n_8601, csa_tree_add_51_79_groupi_n_8602, csa_tree_add_51_79_groupi_n_8603, csa_tree_add_51_79_groupi_n_8604, csa_tree_add_51_79_groupi_n_8605, csa_tree_add_51_79_groupi_n_8606, csa_tree_add_51_79_groupi_n_8607, csa_tree_add_51_79_groupi_n_8608;
  wire csa_tree_add_51_79_groupi_n_8609, csa_tree_add_51_79_groupi_n_8610, csa_tree_add_51_79_groupi_n_8611, csa_tree_add_51_79_groupi_n_8612, csa_tree_add_51_79_groupi_n_8613, csa_tree_add_51_79_groupi_n_8614, csa_tree_add_51_79_groupi_n_8615, csa_tree_add_51_79_groupi_n_8616;
  wire csa_tree_add_51_79_groupi_n_8617, csa_tree_add_51_79_groupi_n_8618, csa_tree_add_51_79_groupi_n_8619, csa_tree_add_51_79_groupi_n_8620, csa_tree_add_51_79_groupi_n_8621, csa_tree_add_51_79_groupi_n_8622, csa_tree_add_51_79_groupi_n_8623, csa_tree_add_51_79_groupi_n_8624;
  wire csa_tree_add_51_79_groupi_n_8625, csa_tree_add_51_79_groupi_n_8626, csa_tree_add_51_79_groupi_n_8627, csa_tree_add_51_79_groupi_n_8628, csa_tree_add_51_79_groupi_n_8629, csa_tree_add_51_79_groupi_n_8630, csa_tree_add_51_79_groupi_n_8631, csa_tree_add_51_79_groupi_n_8632;
  wire csa_tree_add_51_79_groupi_n_8633, csa_tree_add_51_79_groupi_n_8634, csa_tree_add_51_79_groupi_n_8635, csa_tree_add_51_79_groupi_n_8636, csa_tree_add_51_79_groupi_n_8637, csa_tree_add_51_79_groupi_n_8638, csa_tree_add_51_79_groupi_n_8639, csa_tree_add_51_79_groupi_n_8640;
  wire csa_tree_add_51_79_groupi_n_8641, csa_tree_add_51_79_groupi_n_8642, csa_tree_add_51_79_groupi_n_8643, csa_tree_add_51_79_groupi_n_8644, csa_tree_add_51_79_groupi_n_8645, csa_tree_add_51_79_groupi_n_8646, csa_tree_add_51_79_groupi_n_8647, csa_tree_add_51_79_groupi_n_8648;
  wire csa_tree_add_51_79_groupi_n_8649, csa_tree_add_51_79_groupi_n_8650, csa_tree_add_51_79_groupi_n_8651, csa_tree_add_51_79_groupi_n_8652, csa_tree_add_51_79_groupi_n_8653, csa_tree_add_51_79_groupi_n_8654, csa_tree_add_51_79_groupi_n_8655, csa_tree_add_51_79_groupi_n_8656;
  wire csa_tree_add_51_79_groupi_n_8657, csa_tree_add_51_79_groupi_n_8658, csa_tree_add_51_79_groupi_n_8659, csa_tree_add_51_79_groupi_n_8660, csa_tree_add_51_79_groupi_n_8661, csa_tree_add_51_79_groupi_n_8662, csa_tree_add_51_79_groupi_n_8663, csa_tree_add_51_79_groupi_n_8664;
  wire csa_tree_add_51_79_groupi_n_8665, csa_tree_add_51_79_groupi_n_8666, csa_tree_add_51_79_groupi_n_8667, csa_tree_add_51_79_groupi_n_8668, csa_tree_add_51_79_groupi_n_8669, csa_tree_add_51_79_groupi_n_8670, csa_tree_add_51_79_groupi_n_8671, csa_tree_add_51_79_groupi_n_8672;
  wire csa_tree_add_51_79_groupi_n_8673, csa_tree_add_51_79_groupi_n_8674, csa_tree_add_51_79_groupi_n_8675, csa_tree_add_51_79_groupi_n_8676, csa_tree_add_51_79_groupi_n_8677, csa_tree_add_51_79_groupi_n_8678, csa_tree_add_51_79_groupi_n_8679, csa_tree_add_51_79_groupi_n_8680;
  wire csa_tree_add_51_79_groupi_n_8681, csa_tree_add_51_79_groupi_n_8682, csa_tree_add_51_79_groupi_n_8683, csa_tree_add_51_79_groupi_n_8684, csa_tree_add_51_79_groupi_n_8685, csa_tree_add_51_79_groupi_n_8686, csa_tree_add_51_79_groupi_n_8687, csa_tree_add_51_79_groupi_n_8688;
  wire csa_tree_add_51_79_groupi_n_8689, csa_tree_add_51_79_groupi_n_8690, csa_tree_add_51_79_groupi_n_8691, csa_tree_add_51_79_groupi_n_8692, csa_tree_add_51_79_groupi_n_8693, csa_tree_add_51_79_groupi_n_8694, csa_tree_add_51_79_groupi_n_8695, csa_tree_add_51_79_groupi_n_8696;
  wire csa_tree_add_51_79_groupi_n_8697, csa_tree_add_51_79_groupi_n_8698, csa_tree_add_51_79_groupi_n_8699, csa_tree_add_51_79_groupi_n_8700, csa_tree_add_51_79_groupi_n_8701, csa_tree_add_51_79_groupi_n_8702, csa_tree_add_51_79_groupi_n_8703, csa_tree_add_51_79_groupi_n_8704;
  wire csa_tree_add_51_79_groupi_n_8705, csa_tree_add_51_79_groupi_n_8706, csa_tree_add_51_79_groupi_n_8707, csa_tree_add_51_79_groupi_n_8708, csa_tree_add_51_79_groupi_n_8709, csa_tree_add_51_79_groupi_n_8710, csa_tree_add_51_79_groupi_n_8711, csa_tree_add_51_79_groupi_n_8712;
  wire csa_tree_add_51_79_groupi_n_8713, csa_tree_add_51_79_groupi_n_8714, csa_tree_add_51_79_groupi_n_8715, csa_tree_add_51_79_groupi_n_8716, csa_tree_add_51_79_groupi_n_8717, csa_tree_add_51_79_groupi_n_8718, csa_tree_add_51_79_groupi_n_8719, csa_tree_add_51_79_groupi_n_8720;
  wire csa_tree_add_51_79_groupi_n_8721, csa_tree_add_51_79_groupi_n_8722, csa_tree_add_51_79_groupi_n_8723, csa_tree_add_51_79_groupi_n_8724, csa_tree_add_51_79_groupi_n_8725, csa_tree_add_51_79_groupi_n_8726, csa_tree_add_51_79_groupi_n_8727, csa_tree_add_51_79_groupi_n_8728;
  wire csa_tree_add_51_79_groupi_n_8729, csa_tree_add_51_79_groupi_n_8730, csa_tree_add_51_79_groupi_n_8731, csa_tree_add_51_79_groupi_n_8732, csa_tree_add_51_79_groupi_n_8733, csa_tree_add_51_79_groupi_n_8734, csa_tree_add_51_79_groupi_n_8735, csa_tree_add_51_79_groupi_n_8736;
  wire csa_tree_add_51_79_groupi_n_8737, csa_tree_add_51_79_groupi_n_8738, csa_tree_add_51_79_groupi_n_8739, csa_tree_add_51_79_groupi_n_8740, csa_tree_add_51_79_groupi_n_8741, csa_tree_add_51_79_groupi_n_8742, csa_tree_add_51_79_groupi_n_8743, csa_tree_add_51_79_groupi_n_8744;
  wire csa_tree_add_51_79_groupi_n_8745, csa_tree_add_51_79_groupi_n_8746, csa_tree_add_51_79_groupi_n_8747, csa_tree_add_51_79_groupi_n_8748, csa_tree_add_51_79_groupi_n_8749, csa_tree_add_51_79_groupi_n_8750, csa_tree_add_51_79_groupi_n_8751, csa_tree_add_51_79_groupi_n_8752;
  wire csa_tree_add_51_79_groupi_n_8753, csa_tree_add_51_79_groupi_n_8754, csa_tree_add_51_79_groupi_n_8755, csa_tree_add_51_79_groupi_n_8756, csa_tree_add_51_79_groupi_n_8757, csa_tree_add_51_79_groupi_n_8758, csa_tree_add_51_79_groupi_n_8759, csa_tree_add_51_79_groupi_n_8760;
  wire csa_tree_add_51_79_groupi_n_8761, csa_tree_add_51_79_groupi_n_8762, csa_tree_add_51_79_groupi_n_8763, csa_tree_add_51_79_groupi_n_8764, csa_tree_add_51_79_groupi_n_8765, csa_tree_add_51_79_groupi_n_8766, csa_tree_add_51_79_groupi_n_8767, csa_tree_add_51_79_groupi_n_8768;
  wire csa_tree_add_51_79_groupi_n_8769, csa_tree_add_51_79_groupi_n_8770, csa_tree_add_51_79_groupi_n_8771, csa_tree_add_51_79_groupi_n_8772, csa_tree_add_51_79_groupi_n_8773, csa_tree_add_51_79_groupi_n_8774, csa_tree_add_51_79_groupi_n_8775, csa_tree_add_51_79_groupi_n_8776;
  wire csa_tree_add_51_79_groupi_n_8777, csa_tree_add_51_79_groupi_n_8778, csa_tree_add_51_79_groupi_n_8779, csa_tree_add_51_79_groupi_n_8780, csa_tree_add_51_79_groupi_n_8781, csa_tree_add_51_79_groupi_n_8782, csa_tree_add_51_79_groupi_n_8783, csa_tree_add_51_79_groupi_n_8784;
  wire csa_tree_add_51_79_groupi_n_8785, csa_tree_add_51_79_groupi_n_8786, csa_tree_add_51_79_groupi_n_8787, csa_tree_add_51_79_groupi_n_8788, csa_tree_add_51_79_groupi_n_8789, csa_tree_add_51_79_groupi_n_8790, csa_tree_add_51_79_groupi_n_8791, csa_tree_add_51_79_groupi_n_8792;
  wire csa_tree_add_51_79_groupi_n_8793, csa_tree_add_51_79_groupi_n_8794, csa_tree_add_51_79_groupi_n_8795, csa_tree_add_51_79_groupi_n_8796, csa_tree_add_51_79_groupi_n_8797, csa_tree_add_51_79_groupi_n_8798, csa_tree_add_51_79_groupi_n_8799, csa_tree_add_51_79_groupi_n_8800;
  wire csa_tree_add_51_79_groupi_n_8801, csa_tree_add_51_79_groupi_n_8802, csa_tree_add_51_79_groupi_n_8803, csa_tree_add_51_79_groupi_n_8804, csa_tree_add_51_79_groupi_n_8805, csa_tree_add_51_79_groupi_n_8806, csa_tree_add_51_79_groupi_n_8807, csa_tree_add_51_79_groupi_n_8808;
  wire csa_tree_add_51_79_groupi_n_8809, csa_tree_add_51_79_groupi_n_8810, csa_tree_add_51_79_groupi_n_8811, csa_tree_add_51_79_groupi_n_8812, csa_tree_add_51_79_groupi_n_8813, csa_tree_add_51_79_groupi_n_8814, csa_tree_add_51_79_groupi_n_8815, csa_tree_add_51_79_groupi_n_8816;
  wire csa_tree_add_51_79_groupi_n_8817, csa_tree_add_51_79_groupi_n_8818, csa_tree_add_51_79_groupi_n_8819, csa_tree_add_51_79_groupi_n_8820, csa_tree_add_51_79_groupi_n_8821, csa_tree_add_51_79_groupi_n_8822, csa_tree_add_51_79_groupi_n_8823, csa_tree_add_51_79_groupi_n_8824;
  wire csa_tree_add_51_79_groupi_n_8825, csa_tree_add_51_79_groupi_n_8826, csa_tree_add_51_79_groupi_n_8827, csa_tree_add_51_79_groupi_n_8828, csa_tree_add_51_79_groupi_n_8829, csa_tree_add_51_79_groupi_n_8830, csa_tree_add_51_79_groupi_n_8831, csa_tree_add_51_79_groupi_n_8832;
  wire csa_tree_add_51_79_groupi_n_8833, csa_tree_add_51_79_groupi_n_8834, csa_tree_add_51_79_groupi_n_8835, csa_tree_add_51_79_groupi_n_8836, csa_tree_add_51_79_groupi_n_8837, csa_tree_add_51_79_groupi_n_8838, csa_tree_add_51_79_groupi_n_8839, csa_tree_add_51_79_groupi_n_8840;
  wire csa_tree_add_51_79_groupi_n_8841, csa_tree_add_51_79_groupi_n_8842, csa_tree_add_51_79_groupi_n_8843, csa_tree_add_51_79_groupi_n_8844, csa_tree_add_51_79_groupi_n_8845, csa_tree_add_51_79_groupi_n_8846, csa_tree_add_51_79_groupi_n_8847, csa_tree_add_51_79_groupi_n_8848;
  wire csa_tree_add_51_79_groupi_n_8849, csa_tree_add_51_79_groupi_n_8850, csa_tree_add_51_79_groupi_n_8851, csa_tree_add_51_79_groupi_n_8852, csa_tree_add_51_79_groupi_n_8853, csa_tree_add_51_79_groupi_n_8854, csa_tree_add_51_79_groupi_n_8855, csa_tree_add_51_79_groupi_n_8856;
  wire csa_tree_add_51_79_groupi_n_8857, csa_tree_add_51_79_groupi_n_8858, csa_tree_add_51_79_groupi_n_8859, csa_tree_add_51_79_groupi_n_8860, csa_tree_add_51_79_groupi_n_8861, csa_tree_add_51_79_groupi_n_8862, csa_tree_add_51_79_groupi_n_8863, csa_tree_add_51_79_groupi_n_8864;
  wire csa_tree_add_51_79_groupi_n_8865, csa_tree_add_51_79_groupi_n_8866, csa_tree_add_51_79_groupi_n_8867, csa_tree_add_51_79_groupi_n_8868, csa_tree_add_51_79_groupi_n_8869, csa_tree_add_51_79_groupi_n_8870, csa_tree_add_51_79_groupi_n_8871, csa_tree_add_51_79_groupi_n_8872;
  wire csa_tree_add_51_79_groupi_n_8873, csa_tree_add_51_79_groupi_n_8874, csa_tree_add_51_79_groupi_n_8875, csa_tree_add_51_79_groupi_n_8876, csa_tree_add_51_79_groupi_n_8877, csa_tree_add_51_79_groupi_n_8878, csa_tree_add_51_79_groupi_n_8879, csa_tree_add_51_79_groupi_n_8880;
  wire csa_tree_add_51_79_groupi_n_8881, csa_tree_add_51_79_groupi_n_8882, csa_tree_add_51_79_groupi_n_8883, csa_tree_add_51_79_groupi_n_8884, csa_tree_add_51_79_groupi_n_8885, csa_tree_add_51_79_groupi_n_8886, csa_tree_add_51_79_groupi_n_8887, csa_tree_add_51_79_groupi_n_8888;
  wire csa_tree_add_51_79_groupi_n_8889, csa_tree_add_51_79_groupi_n_8890, csa_tree_add_51_79_groupi_n_8891, csa_tree_add_51_79_groupi_n_8892, csa_tree_add_51_79_groupi_n_8893, csa_tree_add_51_79_groupi_n_8894, csa_tree_add_51_79_groupi_n_8895, csa_tree_add_51_79_groupi_n_8896;
  wire csa_tree_add_51_79_groupi_n_8897, csa_tree_add_51_79_groupi_n_8898, csa_tree_add_51_79_groupi_n_8899, csa_tree_add_51_79_groupi_n_8900, csa_tree_add_51_79_groupi_n_8901, csa_tree_add_51_79_groupi_n_8902, csa_tree_add_51_79_groupi_n_8903, csa_tree_add_51_79_groupi_n_8904;
  wire csa_tree_add_51_79_groupi_n_8905, csa_tree_add_51_79_groupi_n_8906, csa_tree_add_51_79_groupi_n_8907, csa_tree_add_51_79_groupi_n_8908, csa_tree_add_51_79_groupi_n_8909, csa_tree_add_51_79_groupi_n_8910, csa_tree_add_51_79_groupi_n_8911, csa_tree_add_51_79_groupi_n_8912;
  wire csa_tree_add_51_79_groupi_n_8913, csa_tree_add_51_79_groupi_n_8914, csa_tree_add_51_79_groupi_n_8915, csa_tree_add_51_79_groupi_n_8916, csa_tree_add_51_79_groupi_n_8917, csa_tree_add_51_79_groupi_n_8918, csa_tree_add_51_79_groupi_n_8919, csa_tree_add_51_79_groupi_n_8920;
  wire csa_tree_add_51_79_groupi_n_8921, csa_tree_add_51_79_groupi_n_8922, csa_tree_add_51_79_groupi_n_8923, csa_tree_add_51_79_groupi_n_8924, csa_tree_add_51_79_groupi_n_8925, csa_tree_add_51_79_groupi_n_8926, csa_tree_add_51_79_groupi_n_8927, csa_tree_add_51_79_groupi_n_8928;
  wire csa_tree_add_51_79_groupi_n_8929, csa_tree_add_51_79_groupi_n_8930, csa_tree_add_51_79_groupi_n_8931, csa_tree_add_51_79_groupi_n_8932, csa_tree_add_51_79_groupi_n_8933, csa_tree_add_51_79_groupi_n_8934, csa_tree_add_51_79_groupi_n_8935, csa_tree_add_51_79_groupi_n_8936;
  wire csa_tree_add_51_79_groupi_n_8937, csa_tree_add_51_79_groupi_n_8938, csa_tree_add_51_79_groupi_n_8939, csa_tree_add_51_79_groupi_n_8940, csa_tree_add_51_79_groupi_n_8941, csa_tree_add_51_79_groupi_n_8942, csa_tree_add_51_79_groupi_n_8943, csa_tree_add_51_79_groupi_n_8944;
  wire csa_tree_add_51_79_groupi_n_8945, csa_tree_add_51_79_groupi_n_8946, csa_tree_add_51_79_groupi_n_8947, csa_tree_add_51_79_groupi_n_8948, csa_tree_add_51_79_groupi_n_8949, csa_tree_add_51_79_groupi_n_8950, csa_tree_add_51_79_groupi_n_8951, csa_tree_add_51_79_groupi_n_8952;
  wire csa_tree_add_51_79_groupi_n_8953, csa_tree_add_51_79_groupi_n_8954, csa_tree_add_51_79_groupi_n_8955, csa_tree_add_51_79_groupi_n_8956, csa_tree_add_51_79_groupi_n_8957, csa_tree_add_51_79_groupi_n_8958, csa_tree_add_51_79_groupi_n_8959, csa_tree_add_51_79_groupi_n_8960;
  wire csa_tree_add_51_79_groupi_n_8961, csa_tree_add_51_79_groupi_n_8962, csa_tree_add_51_79_groupi_n_8963, csa_tree_add_51_79_groupi_n_8964, csa_tree_add_51_79_groupi_n_8965, csa_tree_add_51_79_groupi_n_8966, csa_tree_add_51_79_groupi_n_8967, csa_tree_add_51_79_groupi_n_8968;
  wire csa_tree_add_51_79_groupi_n_8969, csa_tree_add_51_79_groupi_n_8970, csa_tree_add_51_79_groupi_n_8971, csa_tree_add_51_79_groupi_n_8972, csa_tree_add_51_79_groupi_n_8973, csa_tree_add_51_79_groupi_n_8974, csa_tree_add_51_79_groupi_n_8975, csa_tree_add_51_79_groupi_n_8976;
  wire csa_tree_add_51_79_groupi_n_8977, csa_tree_add_51_79_groupi_n_8978, csa_tree_add_51_79_groupi_n_8979, csa_tree_add_51_79_groupi_n_8980, csa_tree_add_51_79_groupi_n_8981, csa_tree_add_51_79_groupi_n_8982, csa_tree_add_51_79_groupi_n_8983, csa_tree_add_51_79_groupi_n_8984;
  wire csa_tree_add_51_79_groupi_n_8985, csa_tree_add_51_79_groupi_n_8986, csa_tree_add_51_79_groupi_n_8987, csa_tree_add_51_79_groupi_n_8988, csa_tree_add_51_79_groupi_n_8989, csa_tree_add_51_79_groupi_n_8990, csa_tree_add_51_79_groupi_n_8991, csa_tree_add_51_79_groupi_n_8992;
  wire csa_tree_add_51_79_groupi_n_8993, csa_tree_add_51_79_groupi_n_8994, csa_tree_add_51_79_groupi_n_8995, csa_tree_add_51_79_groupi_n_8996, csa_tree_add_51_79_groupi_n_8997, csa_tree_add_51_79_groupi_n_8998, csa_tree_add_51_79_groupi_n_8999, csa_tree_add_51_79_groupi_n_9000;
  wire csa_tree_add_51_79_groupi_n_9001, csa_tree_add_51_79_groupi_n_9002, csa_tree_add_51_79_groupi_n_9003, csa_tree_add_51_79_groupi_n_9004, csa_tree_add_51_79_groupi_n_9005, csa_tree_add_51_79_groupi_n_9006, csa_tree_add_51_79_groupi_n_9007, csa_tree_add_51_79_groupi_n_9008;
  wire csa_tree_add_51_79_groupi_n_9009, csa_tree_add_51_79_groupi_n_9010, csa_tree_add_51_79_groupi_n_9011, csa_tree_add_51_79_groupi_n_9012, csa_tree_add_51_79_groupi_n_9013, csa_tree_add_51_79_groupi_n_9014, csa_tree_add_51_79_groupi_n_9015, csa_tree_add_51_79_groupi_n_9016;
  wire csa_tree_add_51_79_groupi_n_9017, csa_tree_add_51_79_groupi_n_9018, csa_tree_add_51_79_groupi_n_9019, csa_tree_add_51_79_groupi_n_9020, csa_tree_add_51_79_groupi_n_9021, csa_tree_add_51_79_groupi_n_9022, csa_tree_add_51_79_groupi_n_9023, csa_tree_add_51_79_groupi_n_9024;
  wire csa_tree_add_51_79_groupi_n_9025, csa_tree_add_51_79_groupi_n_9026, csa_tree_add_51_79_groupi_n_9027, csa_tree_add_51_79_groupi_n_9028, csa_tree_add_51_79_groupi_n_9029, csa_tree_add_51_79_groupi_n_9030, csa_tree_add_51_79_groupi_n_9031, csa_tree_add_51_79_groupi_n_9032;
  wire csa_tree_add_51_79_groupi_n_9033, csa_tree_add_51_79_groupi_n_9034, csa_tree_add_51_79_groupi_n_9035, csa_tree_add_51_79_groupi_n_9036, csa_tree_add_51_79_groupi_n_9037, csa_tree_add_51_79_groupi_n_9038, csa_tree_add_51_79_groupi_n_9039, csa_tree_add_51_79_groupi_n_9040;
  wire csa_tree_add_51_79_groupi_n_9041, csa_tree_add_51_79_groupi_n_9042, csa_tree_add_51_79_groupi_n_9043, csa_tree_add_51_79_groupi_n_9044, csa_tree_add_51_79_groupi_n_9045, csa_tree_add_51_79_groupi_n_9046, csa_tree_add_51_79_groupi_n_9047, csa_tree_add_51_79_groupi_n_9048;
  wire csa_tree_add_51_79_groupi_n_9049, csa_tree_add_51_79_groupi_n_9050, csa_tree_add_51_79_groupi_n_9051, csa_tree_add_51_79_groupi_n_9052, csa_tree_add_51_79_groupi_n_9053, csa_tree_add_51_79_groupi_n_9054, csa_tree_add_51_79_groupi_n_9055, csa_tree_add_51_79_groupi_n_9056;
  wire csa_tree_add_51_79_groupi_n_9057, csa_tree_add_51_79_groupi_n_9058, csa_tree_add_51_79_groupi_n_9059, csa_tree_add_51_79_groupi_n_9060, csa_tree_add_51_79_groupi_n_9061, csa_tree_add_51_79_groupi_n_9062, csa_tree_add_51_79_groupi_n_9063, csa_tree_add_51_79_groupi_n_9064;
  wire csa_tree_add_51_79_groupi_n_9065, csa_tree_add_51_79_groupi_n_9066, csa_tree_add_51_79_groupi_n_9067, csa_tree_add_51_79_groupi_n_9068, csa_tree_add_51_79_groupi_n_9069, csa_tree_add_51_79_groupi_n_9070, csa_tree_add_51_79_groupi_n_9071, csa_tree_add_51_79_groupi_n_9072;
  wire csa_tree_add_51_79_groupi_n_9073, csa_tree_add_51_79_groupi_n_9074, csa_tree_add_51_79_groupi_n_9075, csa_tree_add_51_79_groupi_n_9076, csa_tree_add_51_79_groupi_n_9077, csa_tree_add_51_79_groupi_n_9078, csa_tree_add_51_79_groupi_n_9079, csa_tree_add_51_79_groupi_n_9080;
  wire csa_tree_add_51_79_groupi_n_9081, csa_tree_add_51_79_groupi_n_9082, csa_tree_add_51_79_groupi_n_9083, csa_tree_add_51_79_groupi_n_9084, csa_tree_add_51_79_groupi_n_9085, csa_tree_add_51_79_groupi_n_9086, csa_tree_add_51_79_groupi_n_9087, csa_tree_add_51_79_groupi_n_9088;
  wire csa_tree_add_51_79_groupi_n_9089, csa_tree_add_51_79_groupi_n_9090, csa_tree_add_51_79_groupi_n_9091, csa_tree_add_51_79_groupi_n_9092, csa_tree_add_51_79_groupi_n_9093, csa_tree_add_51_79_groupi_n_9094, csa_tree_add_51_79_groupi_n_9095, csa_tree_add_51_79_groupi_n_9096;
  wire csa_tree_add_51_79_groupi_n_9097, csa_tree_add_51_79_groupi_n_9098, csa_tree_add_51_79_groupi_n_9099, csa_tree_add_51_79_groupi_n_9100, csa_tree_add_51_79_groupi_n_9101, csa_tree_add_51_79_groupi_n_9102, csa_tree_add_51_79_groupi_n_9103, csa_tree_add_51_79_groupi_n_9104;
  wire csa_tree_add_51_79_groupi_n_9105, csa_tree_add_51_79_groupi_n_9106, csa_tree_add_51_79_groupi_n_9107, csa_tree_add_51_79_groupi_n_9108, csa_tree_add_51_79_groupi_n_9109, csa_tree_add_51_79_groupi_n_9110, csa_tree_add_51_79_groupi_n_9111, csa_tree_add_51_79_groupi_n_9112;
  wire csa_tree_add_51_79_groupi_n_9113, csa_tree_add_51_79_groupi_n_9114, csa_tree_add_51_79_groupi_n_9115, csa_tree_add_51_79_groupi_n_9116, csa_tree_add_51_79_groupi_n_9117, csa_tree_add_51_79_groupi_n_9118, csa_tree_add_51_79_groupi_n_9119, csa_tree_add_51_79_groupi_n_9120;
  wire csa_tree_add_51_79_groupi_n_9121, csa_tree_add_51_79_groupi_n_9122, csa_tree_add_51_79_groupi_n_9123, csa_tree_add_51_79_groupi_n_9124, csa_tree_add_51_79_groupi_n_9125, csa_tree_add_51_79_groupi_n_9126, csa_tree_add_51_79_groupi_n_9127, csa_tree_add_51_79_groupi_n_9128;
  wire csa_tree_add_51_79_groupi_n_9129, csa_tree_add_51_79_groupi_n_9130, csa_tree_add_51_79_groupi_n_9131, csa_tree_add_51_79_groupi_n_9132, csa_tree_add_51_79_groupi_n_9133, csa_tree_add_51_79_groupi_n_9134, csa_tree_add_51_79_groupi_n_9135, csa_tree_add_51_79_groupi_n_9136;
  wire csa_tree_add_51_79_groupi_n_9137, csa_tree_add_51_79_groupi_n_9138, csa_tree_add_51_79_groupi_n_9139, csa_tree_add_51_79_groupi_n_9140, csa_tree_add_51_79_groupi_n_9141, csa_tree_add_51_79_groupi_n_9142, csa_tree_add_51_79_groupi_n_9143, csa_tree_add_51_79_groupi_n_9144;
  wire csa_tree_add_51_79_groupi_n_9145, csa_tree_add_51_79_groupi_n_9146, csa_tree_add_51_79_groupi_n_9147, csa_tree_add_51_79_groupi_n_9148, csa_tree_add_51_79_groupi_n_9149, csa_tree_add_51_79_groupi_n_9150, csa_tree_add_51_79_groupi_n_9151, csa_tree_add_51_79_groupi_n_9152;
  wire csa_tree_add_51_79_groupi_n_9153, csa_tree_add_51_79_groupi_n_9154, csa_tree_add_51_79_groupi_n_9155, csa_tree_add_51_79_groupi_n_9156, csa_tree_add_51_79_groupi_n_9157, csa_tree_add_51_79_groupi_n_9158, csa_tree_add_51_79_groupi_n_9159, csa_tree_add_51_79_groupi_n_9160;
  wire csa_tree_add_51_79_groupi_n_9161, csa_tree_add_51_79_groupi_n_9162, csa_tree_add_51_79_groupi_n_9163, csa_tree_add_51_79_groupi_n_9164, csa_tree_add_51_79_groupi_n_9165, csa_tree_add_51_79_groupi_n_9166, csa_tree_add_51_79_groupi_n_9167, csa_tree_add_51_79_groupi_n_9168;
  wire csa_tree_add_51_79_groupi_n_9169, csa_tree_add_51_79_groupi_n_9170, csa_tree_add_51_79_groupi_n_9171, csa_tree_add_51_79_groupi_n_9172, csa_tree_add_51_79_groupi_n_9173, csa_tree_add_51_79_groupi_n_9174, csa_tree_add_51_79_groupi_n_9175, csa_tree_add_51_79_groupi_n_9176;
  wire csa_tree_add_51_79_groupi_n_9177, csa_tree_add_51_79_groupi_n_9178, csa_tree_add_51_79_groupi_n_9179, csa_tree_add_51_79_groupi_n_9180, csa_tree_add_51_79_groupi_n_9181, csa_tree_add_51_79_groupi_n_9182, csa_tree_add_51_79_groupi_n_9183, csa_tree_add_51_79_groupi_n_9184;
  wire csa_tree_add_51_79_groupi_n_9185, csa_tree_add_51_79_groupi_n_9186, csa_tree_add_51_79_groupi_n_9187, csa_tree_add_51_79_groupi_n_9188, csa_tree_add_51_79_groupi_n_9189, csa_tree_add_51_79_groupi_n_9190, csa_tree_add_51_79_groupi_n_9191, csa_tree_add_51_79_groupi_n_9192;
  wire csa_tree_add_51_79_groupi_n_9193, csa_tree_add_51_79_groupi_n_9194, csa_tree_add_51_79_groupi_n_9195, csa_tree_add_51_79_groupi_n_9196, csa_tree_add_51_79_groupi_n_9197, csa_tree_add_51_79_groupi_n_9198, csa_tree_add_51_79_groupi_n_9199, csa_tree_add_51_79_groupi_n_9200;
  wire csa_tree_add_51_79_groupi_n_9201, csa_tree_add_51_79_groupi_n_9202, csa_tree_add_51_79_groupi_n_9203, csa_tree_add_51_79_groupi_n_9204, csa_tree_add_51_79_groupi_n_9205, csa_tree_add_51_79_groupi_n_9206, csa_tree_add_51_79_groupi_n_9207, csa_tree_add_51_79_groupi_n_9208;
  wire csa_tree_add_51_79_groupi_n_9209, csa_tree_add_51_79_groupi_n_9210, csa_tree_add_51_79_groupi_n_9211, csa_tree_add_51_79_groupi_n_9212, csa_tree_add_51_79_groupi_n_9213, csa_tree_add_51_79_groupi_n_9214, csa_tree_add_51_79_groupi_n_9215, csa_tree_add_51_79_groupi_n_9216;
  wire csa_tree_add_51_79_groupi_n_9217, csa_tree_add_51_79_groupi_n_9218, csa_tree_add_51_79_groupi_n_9219, csa_tree_add_51_79_groupi_n_9220, csa_tree_add_51_79_groupi_n_9221, csa_tree_add_51_79_groupi_n_9222, csa_tree_add_51_79_groupi_n_9223, csa_tree_add_51_79_groupi_n_9224;
  wire csa_tree_add_51_79_groupi_n_9225, csa_tree_add_51_79_groupi_n_9226, csa_tree_add_51_79_groupi_n_9227, csa_tree_add_51_79_groupi_n_9228, csa_tree_add_51_79_groupi_n_9229, csa_tree_add_51_79_groupi_n_9230, csa_tree_add_51_79_groupi_n_9231, csa_tree_add_51_79_groupi_n_9232;
  wire csa_tree_add_51_79_groupi_n_9233, csa_tree_add_51_79_groupi_n_9234, csa_tree_add_51_79_groupi_n_9235, csa_tree_add_51_79_groupi_n_9236, csa_tree_add_51_79_groupi_n_9237, csa_tree_add_51_79_groupi_n_9238, csa_tree_add_51_79_groupi_n_9239, csa_tree_add_51_79_groupi_n_9240;
  wire csa_tree_add_51_79_groupi_n_9241, csa_tree_add_51_79_groupi_n_9242, csa_tree_add_51_79_groupi_n_9243, csa_tree_add_51_79_groupi_n_9244, csa_tree_add_51_79_groupi_n_9245, csa_tree_add_51_79_groupi_n_9246, csa_tree_add_51_79_groupi_n_9247, csa_tree_add_51_79_groupi_n_9248;
  wire csa_tree_add_51_79_groupi_n_9249, csa_tree_add_51_79_groupi_n_9250, csa_tree_add_51_79_groupi_n_9251, csa_tree_add_51_79_groupi_n_9252, csa_tree_add_51_79_groupi_n_9253, csa_tree_add_51_79_groupi_n_9254, csa_tree_add_51_79_groupi_n_9255, csa_tree_add_51_79_groupi_n_9256;
  wire csa_tree_add_51_79_groupi_n_9257, csa_tree_add_51_79_groupi_n_9258, csa_tree_add_51_79_groupi_n_9259, csa_tree_add_51_79_groupi_n_9260, csa_tree_add_51_79_groupi_n_9261, csa_tree_add_51_79_groupi_n_9262, csa_tree_add_51_79_groupi_n_9263, csa_tree_add_51_79_groupi_n_9264;
  wire csa_tree_add_51_79_groupi_n_9265, csa_tree_add_51_79_groupi_n_9266, csa_tree_add_51_79_groupi_n_9267, csa_tree_add_51_79_groupi_n_9268, csa_tree_add_51_79_groupi_n_9269, csa_tree_add_51_79_groupi_n_9270, csa_tree_add_51_79_groupi_n_9271, csa_tree_add_51_79_groupi_n_9272;
  wire csa_tree_add_51_79_groupi_n_9273, csa_tree_add_51_79_groupi_n_9274, csa_tree_add_51_79_groupi_n_9275, csa_tree_add_51_79_groupi_n_9276, csa_tree_add_51_79_groupi_n_9277, csa_tree_add_51_79_groupi_n_9278, csa_tree_add_51_79_groupi_n_9279, csa_tree_add_51_79_groupi_n_9280;
  wire csa_tree_add_51_79_groupi_n_9281, csa_tree_add_51_79_groupi_n_9282, csa_tree_add_51_79_groupi_n_9283, csa_tree_add_51_79_groupi_n_9284, csa_tree_add_51_79_groupi_n_9285, csa_tree_add_51_79_groupi_n_9286, csa_tree_add_51_79_groupi_n_9287, csa_tree_add_51_79_groupi_n_9288;
  wire csa_tree_add_51_79_groupi_n_9289, csa_tree_add_51_79_groupi_n_9290, csa_tree_add_51_79_groupi_n_9291, csa_tree_add_51_79_groupi_n_9292, csa_tree_add_51_79_groupi_n_9293, csa_tree_add_51_79_groupi_n_9294, csa_tree_add_51_79_groupi_n_9295, csa_tree_add_51_79_groupi_n_9296;
  wire csa_tree_add_51_79_groupi_n_9297, csa_tree_add_51_79_groupi_n_9298, csa_tree_add_51_79_groupi_n_9299, csa_tree_add_51_79_groupi_n_9300, csa_tree_add_51_79_groupi_n_9301, csa_tree_add_51_79_groupi_n_9302, csa_tree_add_51_79_groupi_n_9303, csa_tree_add_51_79_groupi_n_9304;
  wire csa_tree_add_51_79_groupi_n_9305, csa_tree_add_51_79_groupi_n_9306, csa_tree_add_51_79_groupi_n_9307, csa_tree_add_51_79_groupi_n_9308, csa_tree_add_51_79_groupi_n_9309, csa_tree_add_51_79_groupi_n_9310, csa_tree_add_51_79_groupi_n_9311, csa_tree_add_51_79_groupi_n_9312;
  wire csa_tree_add_51_79_groupi_n_9313, csa_tree_add_51_79_groupi_n_9314, csa_tree_add_51_79_groupi_n_9315, csa_tree_add_51_79_groupi_n_9316, csa_tree_add_51_79_groupi_n_9317, csa_tree_add_51_79_groupi_n_9318, csa_tree_add_51_79_groupi_n_9319, csa_tree_add_51_79_groupi_n_9320;
  wire csa_tree_add_51_79_groupi_n_9321, csa_tree_add_51_79_groupi_n_9322, csa_tree_add_51_79_groupi_n_9323, csa_tree_add_51_79_groupi_n_9324, csa_tree_add_51_79_groupi_n_9325, csa_tree_add_51_79_groupi_n_9326, csa_tree_add_51_79_groupi_n_9327, csa_tree_add_51_79_groupi_n_9328;
  wire csa_tree_add_51_79_groupi_n_9329, csa_tree_add_51_79_groupi_n_9330, csa_tree_add_51_79_groupi_n_9331, csa_tree_add_51_79_groupi_n_9332, csa_tree_add_51_79_groupi_n_9333, csa_tree_add_51_79_groupi_n_9334, csa_tree_add_51_79_groupi_n_9335, csa_tree_add_51_79_groupi_n_9336;
  wire csa_tree_add_51_79_groupi_n_9337, csa_tree_add_51_79_groupi_n_9338, csa_tree_add_51_79_groupi_n_9339, csa_tree_add_51_79_groupi_n_9340, csa_tree_add_51_79_groupi_n_9341, csa_tree_add_51_79_groupi_n_9342, csa_tree_add_51_79_groupi_n_9343, csa_tree_add_51_79_groupi_n_9344;
  wire csa_tree_add_51_79_groupi_n_9345, csa_tree_add_51_79_groupi_n_9346, csa_tree_add_51_79_groupi_n_9347, csa_tree_add_51_79_groupi_n_9348, csa_tree_add_51_79_groupi_n_9349, csa_tree_add_51_79_groupi_n_9350, csa_tree_add_51_79_groupi_n_9351, csa_tree_add_51_79_groupi_n_9352;
  wire csa_tree_add_51_79_groupi_n_9353, csa_tree_add_51_79_groupi_n_9354, csa_tree_add_51_79_groupi_n_9355, csa_tree_add_51_79_groupi_n_9356, csa_tree_add_51_79_groupi_n_9357, csa_tree_add_51_79_groupi_n_9358, csa_tree_add_51_79_groupi_n_9359, csa_tree_add_51_79_groupi_n_9360;
  wire csa_tree_add_51_79_groupi_n_9361, csa_tree_add_51_79_groupi_n_9362, csa_tree_add_51_79_groupi_n_9363, csa_tree_add_51_79_groupi_n_9364, csa_tree_add_51_79_groupi_n_9365, csa_tree_add_51_79_groupi_n_9366, csa_tree_add_51_79_groupi_n_9367, csa_tree_add_51_79_groupi_n_9368;
  wire csa_tree_add_51_79_groupi_n_9369, csa_tree_add_51_79_groupi_n_9370, csa_tree_add_51_79_groupi_n_9371, csa_tree_add_51_79_groupi_n_9372, csa_tree_add_51_79_groupi_n_9373, csa_tree_add_51_79_groupi_n_9374, csa_tree_add_51_79_groupi_n_9375, csa_tree_add_51_79_groupi_n_9376;
  wire csa_tree_add_51_79_groupi_n_9377, csa_tree_add_51_79_groupi_n_9378, csa_tree_add_51_79_groupi_n_9379, csa_tree_add_51_79_groupi_n_9380, csa_tree_add_51_79_groupi_n_9381, csa_tree_add_51_79_groupi_n_9382, csa_tree_add_51_79_groupi_n_9383, csa_tree_add_51_79_groupi_n_9384;
  wire csa_tree_add_51_79_groupi_n_9385, csa_tree_add_51_79_groupi_n_9386, csa_tree_add_51_79_groupi_n_9387, csa_tree_add_51_79_groupi_n_9388, csa_tree_add_51_79_groupi_n_9389, csa_tree_add_51_79_groupi_n_9390, csa_tree_add_51_79_groupi_n_9391, csa_tree_add_51_79_groupi_n_9392;
  wire csa_tree_add_51_79_groupi_n_9393, csa_tree_add_51_79_groupi_n_9394, csa_tree_add_51_79_groupi_n_9395, csa_tree_add_51_79_groupi_n_9396, csa_tree_add_51_79_groupi_n_9397, csa_tree_add_51_79_groupi_n_9398, csa_tree_add_51_79_groupi_n_9399, csa_tree_add_51_79_groupi_n_9400;
  wire csa_tree_add_51_79_groupi_n_9401, csa_tree_add_51_79_groupi_n_9402, csa_tree_add_51_79_groupi_n_9403, csa_tree_add_51_79_groupi_n_9404, csa_tree_add_51_79_groupi_n_9405, csa_tree_add_51_79_groupi_n_9406, csa_tree_add_51_79_groupi_n_9407, csa_tree_add_51_79_groupi_n_9408;
  wire csa_tree_add_51_79_groupi_n_9409, csa_tree_add_51_79_groupi_n_9410, csa_tree_add_51_79_groupi_n_9411, csa_tree_add_51_79_groupi_n_9412, csa_tree_add_51_79_groupi_n_9413, csa_tree_add_51_79_groupi_n_9414, csa_tree_add_51_79_groupi_n_9415, csa_tree_add_51_79_groupi_n_9416;
  wire csa_tree_add_51_79_groupi_n_9417, csa_tree_add_51_79_groupi_n_9418, csa_tree_add_51_79_groupi_n_9419, csa_tree_add_51_79_groupi_n_9420, csa_tree_add_51_79_groupi_n_9421, csa_tree_add_51_79_groupi_n_9422, csa_tree_add_51_79_groupi_n_9423, csa_tree_add_51_79_groupi_n_9424;
  wire csa_tree_add_51_79_groupi_n_9425, csa_tree_add_51_79_groupi_n_9426, csa_tree_add_51_79_groupi_n_9427, csa_tree_add_51_79_groupi_n_9428, csa_tree_add_51_79_groupi_n_9429, csa_tree_add_51_79_groupi_n_9430, csa_tree_add_51_79_groupi_n_9431, csa_tree_add_51_79_groupi_n_9432;
  wire csa_tree_add_51_79_groupi_n_9433, csa_tree_add_51_79_groupi_n_9434, csa_tree_add_51_79_groupi_n_9435, csa_tree_add_51_79_groupi_n_9436, csa_tree_add_51_79_groupi_n_9437, csa_tree_add_51_79_groupi_n_9438, csa_tree_add_51_79_groupi_n_9439, csa_tree_add_51_79_groupi_n_9440;
  wire csa_tree_add_51_79_groupi_n_9441, csa_tree_add_51_79_groupi_n_9442, csa_tree_add_51_79_groupi_n_9443, csa_tree_add_51_79_groupi_n_9444, csa_tree_add_51_79_groupi_n_9445, csa_tree_add_51_79_groupi_n_9446, csa_tree_add_51_79_groupi_n_9447, csa_tree_add_51_79_groupi_n_9448;
  wire csa_tree_add_51_79_groupi_n_9449, csa_tree_add_51_79_groupi_n_9450, csa_tree_add_51_79_groupi_n_9451, csa_tree_add_51_79_groupi_n_9452, csa_tree_add_51_79_groupi_n_9453, csa_tree_add_51_79_groupi_n_9454, csa_tree_add_51_79_groupi_n_9455, csa_tree_add_51_79_groupi_n_9456;
  wire csa_tree_add_51_79_groupi_n_9457, csa_tree_add_51_79_groupi_n_9458, csa_tree_add_51_79_groupi_n_9459, csa_tree_add_51_79_groupi_n_9460, csa_tree_add_51_79_groupi_n_9461, csa_tree_add_51_79_groupi_n_9462, csa_tree_add_51_79_groupi_n_9463, csa_tree_add_51_79_groupi_n_9464;
  wire csa_tree_add_51_79_groupi_n_9465, csa_tree_add_51_79_groupi_n_9466, csa_tree_add_51_79_groupi_n_9467, csa_tree_add_51_79_groupi_n_9468, csa_tree_add_51_79_groupi_n_9469, csa_tree_add_51_79_groupi_n_9470, csa_tree_add_51_79_groupi_n_9471, csa_tree_add_51_79_groupi_n_9472;
  wire csa_tree_add_51_79_groupi_n_9473, csa_tree_add_51_79_groupi_n_9474, csa_tree_add_51_79_groupi_n_9475, csa_tree_add_51_79_groupi_n_9476, csa_tree_add_51_79_groupi_n_9477, csa_tree_add_51_79_groupi_n_9478, csa_tree_add_51_79_groupi_n_9479, csa_tree_add_51_79_groupi_n_9480;
  wire csa_tree_add_51_79_groupi_n_9481, csa_tree_add_51_79_groupi_n_9482, csa_tree_add_51_79_groupi_n_9483, csa_tree_add_51_79_groupi_n_9484, csa_tree_add_51_79_groupi_n_9485, csa_tree_add_51_79_groupi_n_9486, csa_tree_add_51_79_groupi_n_9487, csa_tree_add_51_79_groupi_n_9488;
  wire csa_tree_add_51_79_groupi_n_9489, csa_tree_add_51_79_groupi_n_9490, csa_tree_add_51_79_groupi_n_9491, csa_tree_add_51_79_groupi_n_9492, csa_tree_add_51_79_groupi_n_9493, csa_tree_add_51_79_groupi_n_9494, csa_tree_add_51_79_groupi_n_9495, csa_tree_add_51_79_groupi_n_9496;
  wire csa_tree_add_51_79_groupi_n_9497, csa_tree_add_51_79_groupi_n_9498, csa_tree_add_51_79_groupi_n_9499, csa_tree_add_51_79_groupi_n_9500, csa_tree_add_51_79_groupi_n_9501, csa_tree_add_51_79_groupi_n_9502, csa_tree_add_51_79_groupi_n_9503, csa_tree_add_51_79_groupi_n_9504;
  wire csa_tree_add_51_79_groupi_n_9505, csa_tree_add_51_79_groupi_n_9506, csa_tree_add_51_79_groupi_n_9507, csa_tree_add_51_79_groupi_n_9508, csa_tree_add_51_79_groupi_n_9509, csa_tree_add_51_79_groupi_n_9510, csa_tree_add_51_79_groupi_n_9511, csa_tree_add_51_79_groupi_n_9512;
  wire csa_tree_add_51_79_groupi_n_9513, csa_tree_add_51_79_groupi_n_9514, csa_tree_add_51_79_groupi_n_9515, csa_tree_add_51_79_groupi_n_9516, csa_tree_add_51_79_groupi_n_9517, csa_tree_add_51_79_groupi_n_9518, csa_tree_add_51_79_groupi_n_9519, csa_tree_add_51_79_groupi_n_9520;
  wire csa_tree_add_51_79_groupi_n_9521, csa_tree_add_51_79_groupi_n_9522, csa_tree_add_51_79_groupi_n_9523, csa_tree_add_51_79_groupi_n_9524, csa_tree_add_51_79_groupi_n_9525, csa_tree_add_51_79_groupi_n_9526, csa_tree_add_51_79_groupi_n_9527, csa_tree_add_51_79_groupi_n_9528;
  wire csa_tree_add_51_79_groupi_n_9529, csa_tree_add_51_79_groupi_n_9530, csa_tree_add_51_79_groupi_n_9531, csa_tree_add_51_79_groupi_n_9532, csa_tree_add_51_79_groupi_n_9533, csa_tree_add_51_79_groupi_n_9534, csa_tree_add_51_79_groupi_n_9535, csa_tree_add_51_79_groupi_n_9536;
  wire csa_tree_add_51_79_groupi_n_9537, csa_tree_add_51_79_groupi_n_9538, csa_tree_add_51_79_groupi_n_9539, csa_tree_add_51_79_groupi_n_9540, csa_tree_add_51_79_groupi_n_9541, csa_tree_add_51_79_groupi_n_9542, csa_tree_add_51_79_groupi_n_9543, csa_tree_add_51_79_groupi_n_9544;
  wire csa_tree_add_51_79_groupi_n_9545, csa_tree_add_51_79_groupi_n_9546, csa_tree_add_51_79_groupi_n_9547, csa_tree_add_51_79_groupi_n_9548, csa_tree_add_51_79_groupi_n_9549, csa_tree_add_51_79_groupi_n_9550, csa_tree_add_51_79_groupi_n_9551, csa_tree_add_51_79_groupi_n_9552;
  wire csa_tree_add_51_79_groupi_n_9553, csa_tree_add_51_79_groupi_n_9554, csa_tree_add_51_79_groupi_n_9555, csa_tree_add_51_79_groupi_n_9556, csa_tree_add_51_79_groupi_n_9557, csa_tree_add_51_79_groupi_n_9558, csa_tree_add_51_79_groupi_n_9559, csa_tree_add_51_79_groupi_n_9560;
  wire csa_tree_add_51_79_groupi_n_9561, csa_tree_add_51_79_groupi_n_9562, csa_tree_add_51_79_groupi_n_9563, csa_tree_add_51_79_groupi_n_9564, csa_tree_add_51_79_groupi_n_9565, csa_tree_add_51_79_groupi_n_9566, csa_tree_add_51_79_groupi_n_9567, csa_tree_add_51_79_groupi_n_9568;
  wire csa_tree_add_51_79_groupi_n_9569, csa_tree_add_51_79_groupi_n_9570, csa_tree_add_51_79_groupi_n_9571, csa_tree_add_51_79_groupi_n_9572, csa_tree_add_51_79_groupi_n_9573, csa_tree_add_51_79_groupi_n_9574, csa_tree_add_51_79_groupi_n_9575, csa_tree_add_51_79_groupi_n_9576;
  wire csa_tree_add_51_79_groupi_n_9577, csa_tree_add_51_79_groupi_n_9578, csa_tree_add_51_79_groupi_n_9579, csa_tree_add_51_79_groupi_n_9580, csa_tree_add_51_79_groupi_n_9581, csa_tree_add_51_79_groupi_n_9582, csa_tree_add_51_79_groupi_n_9583, csa_tree_add_51_79_groupi_n_9584;
  wire csa_tree_add_51_79_groupi_n_9585, csa_tree_add_51_79_groupi_n_9586, csa_tree_add_51_79_groupi_n_9587, csa_tree_add_51_79_groupi_n_9588, csa_tree_add_51_79_groupi_n_9589, csa_tree_add_51_79_groupi_n_9590, csa_tree_add_51_79_groupi_n_9591, csa_tree_add_51_79_groupi_n_9592;
  wire csa_tree_add_51_79_groupi_n_9593, csa_tree_add_51_79_groupi_n_9594, csa_tree_add_51_79_groupi_n_9595, csa_tree_add_51_79_groupi_n_9596, csa_tree_add_51_79_groupi_n_9597, csa_tree_add_51_79_groupi_n_9598, csa_tree_add_51_79_groupi_n_9599, csa_tree_add_51_79_groupi_n_9600;
  wire csa_tree_add_51_79_groupi_n_9601, csa_tree_add_51_79_groupi_n_9602, csa_tree_add_51_79_groupi_n_9603, csa_tree_add_51_79_groupi_n_9604, csa_tree_add_51_79_groupi_n_9605, csa_tree_add_51_79_groupi_n_9606, csa_tree_add_51_79_groupi_n_9607, csa_tree_add_51_79_groupi_n_9608;
  wire csa_tree_add_51_79_groupi_n_9609, csa_tree_add_51_79_groupi_n_9610, csa_tree_add_51_79_groupi_n_9611, csa_tree_add_51_79_groupi_n_9612, csa_tree_add_51_79_groupi_n_9613, csa_tree_add_51_79_groupi_n_9614, csa_tree_add_51_79_groupi_n_9615, csa_tree_add_51_79_groupi_n_9616;
  wire csa_tree_add_51_79_groupi_n_9617, csa_tree_add_51_79_groupi_n_9618, csa_tree_add_51_79_groupi_n_9619, csa_tree_add_51_79_groupi_n_9620, csa_tree_add_51_79_groupi_n_9621, csa_tree_add_51_79_groupi_n_9622, csa_tree_add_51_79_groupi_n_9623, csa_tree_add_51_79_groupi_n_9624;
  wire csa_tree_add_51_79_groupi_n_9625, csa_tree_add_51_79_groupi_n_9626, csa_tree_add_51_79_groupi_n_9627, csa_tree_add_51_79_groupi_n_9628, csa_tree_add_51_79_groupi_n_9629, csa_tree_add_51_79_groupi_n_9630, csa_tree_add_51_79_groupi_n_9631, csa_tree_add_51_79_groupi_n_9632;
  wire csa_tree_add_51_79_groupi_n_9633, csa_tree_add_51_79_groupi_n_9634, csa_tree_add_51_79_groupi_n_9635, csa_tree_add_51_79_groupi_n_9636, csa_tree_add_51_79_groupi_n_9637, csa_tree_add_51_79_groupi_n_9638, csa_tree_add_51_79_groupi_n_9639, csa_tree_add_51_79_groupi_n_9640;
  wire csa_tree_add_51_79_groupi_n_9641, csa_tree_add_51_79_groupi_n_9642, csa_tree_add_51_79_groupi_n_9643, csa_tree_add_51_79_groupi_n_9644, csa_tree_add_51_79_groupi_n_9645, csa_tree_add_51_79_groupi_n_9646, csa_tree_add_51_79_groupi_n_9647, csa_tree_add_51_79_groupi_n_9648;
  wire csa_tree_add_51_79_groupi_n_9649, csa_tree_add_51_79_groupi_n_9650, csa_tree_add_51_79_groupi_n_9651, csa_tree_add_51_79_groupi_n_9652, csa_tree_add_51_79_groupi_n_9653, csa_tree_add_51_79_groupi_n_9654, csa_tree_add_51_79_groupi_n_9655, csa_tree_add_51_79_groupi_n_9656;
  wire csa_tree_add_51_79_groupi_n_9657, csa_tree_add_51_79_groupi_n_9658, csa_tree_add_51_79_groupi_n_9659, csa_tree_add_51_79_groupi_n_9660, csa_tree_add_51_79_groupi_n_9661, csa_tree_add_51_79_groupi_n_9662, csa_tree_add_51_79_groupi_n_9663, csa_tree_add_51_79_groupi_n_9664;
  wire csa_tree_add_51_79_groupi_n_9665, csa_tree_add_51_79_groupi_n_9666, csa_tree_add_51_79_groupi_n_9667, csa_tree_add_51_79_groupi_n_9668, csa_tree_add_51_79_groupi_n_9669, csa_tree_add_51_79_groupi_n_9670, csa_tree_add_51_79_groupi_n_9671, csa_tree_add_51_79_groupi_n_9672;
  wire csa_tree_add_51_79_groupi_n_9673, csa_tree_add_51_79_groupi_n_9674, csa_tree_add_51_79_groupi_n_9675, csa_tree_add_51_79_groupi_n_9676, csa_tree_add_51_79_groupi_n_9677, csa_tree_add_51_79_groupi_n_9678, csa_tree_add_51_79_groupi_n_9679, csa_tree_add_51_79_groupi_n_9680;
  wire csa_tree_add_51_79_groupi_n_9681, csa_tree_add_51_79_groupi_n_9682, csa_tree_add_51_79_groupi_n_9683, csa_tree_add_51_79_groupi_n_9684, csa_tree_add_51_79_groupi_n_9685, csa_tree_add_51_79_groupi_n_9686, csa_tree_add_51_79_groupi_n_9687, csa_tree_add_51_79_groupi_n_9688;
  wire csa_tree_add_51_79_groupi_n_9689, csa_tree_add_51_79_groupi_n_9690, csa_tree_add_51_79_groupi_n_9691, csa_tree_add_51_79_groupi_n_9692, csa_tree_add_51_79_groupi_n_9693, csa_tree_add_51_79_groupi_n_9694, csa_tree_add_51_79_groupi_n_9695, csa_tree_add_51_79_groupi_n_9696;
  wire csa_tree_add_51_79_groupi_n_9697, csa_tree_add_51_79_groupi_n_9698, csa_tree_add_51_79_groupi_n_9699, csa_tree_add_51_79_groupi_n_9700, csa_tree_add_51_79_groupi_n_9701, csa_tree_add_51_79_groupi_n_9702, csa_tree_add_51_79_groupi_n_9703, csa_tree_add_51_79_groupi_n_9704;
  wire csa_tree_add_51_79_groupi_n_9705, csa_tree_add_51_79_groupi_n_9706, csa_tree_add_51_79_groupi_n_9707, csa_tree_add_51_79_groupi_n_9708, csa_tree_add_51_79_groupi_n_9709, csa_tree_add_51_79_groupi_n_9710, csa_tree_add_51_79_groupi_n_9711, csa_tree_add_51_79_groupi_n_9712;
  wire csa_tree_add_51_79_groupi_n_9713, csa_tree_add_51_79_groupi_n_9714, csa_tree_add_51_79_groupi_n_9715, csa_tree_add_51_79_groupi_n_9716, csa_tree_add_51_79_groupi_n_9717, csa_tree_add_51_79_groupi_n_9718, csa_tree_add_51_79_groupi_n_9719, csa_tree_add_51_79_groupi_n_9720;
  wire csa_tree_add_51_79_groupi_n_9721, csa_tree_add_51_79_groupi_n_9722, csa_tree_add_51_79_groupi_n_9723, csa_tree_add_51_79_groupi_n_9724, csa_tree_add_51_79_groupi_n_9725, csa_tree_add_51_79_groupi_n_9726, csa_tree_add_51_79_groupi_n_9727, csa_tree_add_51_79_groupi_n_9728;
  wire csa_tree_add_51_79_groupi_n_9729, csa_tree_add_51_79_groupi_n_9730, csa_tree_add_51_79_groupi_n_9731, csa_tree_add_51_79_groupi_n_9732, csa_tree_add_51_79_groupi_n_9733, csa_tree_add_51_79_groupi_n_9734, csa_tree_add_51_79_groupi_n_9735, csa_tree_add_51_79_groupi_n_9736;
  wire csa_tree_add_51_79_groupi_n_9737, csa_tree_add_51_79_groupi_n_9738, csa_tree_add_51_79_groupi_n_9739, csa_tree_add_51_79_groupi_n_9740, csa_tree_add_51_79_groupi_n_9741, csa_tree_add_51_79_groupi_n_9742, csa_tree_add_51_79_groupi_n_9743, csa_tree_add_51_79_groupi_n_9744;
  wire csa_tree_add_51_79_groupi_n_9745, csa_tree_add_51_79_groupi_n_9746, csa_tree_add_51_79_groupi_n_9747, csa_tree_add_51_79_groupi_n_9748, csa_tree_add_51_79_groupi_n_9749, csa_tree_add_51_79_groupi_n_9750, csa_tree_add_51_79_groupi_n_9751, csa_tree_add_51_79_groupi_n_9752;
  wire csa_tree_add_51_79_groupi_n_9753, csa_tree_add_51_79_groupi_n_9754, csa_tree_add_51_79_groupi_n_9755, csa_tree_add_51_79_groupi_n_9756, csa_tree_add_51_79_groupi_n_9757, csa_tree_add_51_79_groupi_n_9758, csa_tree_add_51_79_groupi_n_9759, csa_tree_add_51_79_groupi_n_9760;
  wire csa_tree_add_51_79_groupi_n_9761, csa_tree_add_51_79_groupi_n_9762, csa_tree_add_51_79_groupi_n_9763, csa_tree_add_51_79_groupi_n_9764, csa_tree_add_51_79_groupi_n_9765, csa_tree_add_51_79_groupi_n_9766, csa_tree_add_51_79_groupi_n_9767, csa_tree_add_51_79_groupi_n_9768;
  wire csa_tree_add_51_79_groupi_n_9769, csa_tree_add_51_79_groupi_n_9770, csa_tree_add_51_79_groupi_n_9771, csa_tree_add_51_79_groupi_n_9772, csa_tree_add_51_79_groupi_n_9773, csa_tree_add_51_79_groupi_n_9774, csa_tree_add_51_79_groupi_n_9775, csa_tree_add_51_79_groupi_n_9776;
  wire csa_tree_add_51_79_groupi_n_9777, csa_tree_add_51_79_groupi_n_9778, csa_tree_add_51_79_groupi_n_9779, csa_tree_add_51_79_groupi_n_9780, csa_tree_add_51_79_groupi_n_9781, csa_tree_add_51_79_groupi_n_9782, csa_tree_add_51_79_groupi_n_9783, csa_tree_add_51_79_groupi_n_9784;
  wire csa_tree_add_51_79_groupi_n_9785, csa_tree_add_51_79_groupi_n_9786, csa_tree_add_51_79_groupi_n_9787, csa_tree_add_51_79_groupi_n_9788, csa_tree_add_51_79_groupi_n_9789, csa_tree_add_51_79_groupi_n_9790, csa_tree_add_51_79_groupi_n_9791, csa_tree_add_51_79_groupi_n_9792;
  wire csa_tree_add_51_79_groupi_n_9793, csa_tree_add_51_79_groupi_n_9794, csa_tree_add_51_79_groupi_n_9795, csa_tree_add_51_79_groupi_n_9796, csa_tree_add_51_79_groupi_n_9797, csa_tree_add_51_79_groupi_n_9798, csa_tree_add_51_79_groupi_n_9799, csa_tree_add_51_79_groupi_n_9800;
  wire csa_tree_add_51_79_groupi_n_9801, csa_tree_add_51_79_groupi_n_9802, csa_tree_add_51_79_groupi_n_9803, csa_tree_add_51_79_groupi_n_9804, csa_tree_add_51_79_groupi_n_9805, csa_tree_add_51_79_groupi_n_9806, csa_tree_add_51_79_groupi_n_9807, csa_tree_add_51_79_groupi_n_9808;
  wire csa_tree_add_51_79_groupi_n_9809, csa_tree_add_51_79_groupi_n_9810, csa_tree_add_51_79_groupi_n_9811, csa_tree_add_51_79_groupi_n_9812, csa_tree_add_51_79_groupi_n_9813, csa_tree_add_51_79_groupi_n_9814, csa_tree_add_51_79_groupi_n_9815, csa_tree_add_51_79_groupi_n_9816;
  wire csa_tree_add_51_79_groupi_n_9817, csa_tree_add_51_79_groupi_n_9818, csa_tree_add_51_79_groupi_n_9819, csa_tree_add_51_79_groupi_n_9820, csa_tree_add_51_79_groupi_n_9821, csa_tree_add_51_79_groupi_n_9822, csa_tree_add_51_79_groupi_n_9823, csa_tree_add_51_79_groupi_n_9824;
  wire csa_tree_add_51_79_groupi_n_9825, csa_tree_add_51_79_groupi_n_9826, csa_tree_add_51_79_groupi_n_9827, csa_tree_add_51_79_groupi_n_9828, csa_tree_add_51_79_groupi_n_9829, csa_tree_add_51_79_groupi_n_9830, csa_tree_add_51_79_groupi_n_9831, csa_tree_add_51_79_groupi_n_9832;
  wire csa_tree_add_51_79_groupi_n_9833, csa_tree_add_51_79_groupi_n_9834, csa_tree_add_51_79_groupi_n_9835, csa_tree_add_51_79_groupi_n_9836, csa_tree_add_51_79_groupi_n_9837, csa_tree_add_51_79_groupi_n_9838, csa_tree_add_51_79_groupi_n_9839, csa_tree_add_51_79_groupi_n_9840;
  wire csa_tree_add_51_79_groupi_n_9841, csa_tree_add_51_79_groupi_n_9842, csa_tree_add_51_79_groupi_n_9843, csa_tree_add_51_79_groupi_n_9844, csa_tree_add_51_79_groupi_n_9845, csa_tree_add_51_79_groupi_n_9846, csa_tree_add_51_79_groupi_n_9847, csa_tree_add_51_79_groupi_n_9848;
  wire csa_tree_add_51_79_groupi_n_9849, csa_tree_add_51_79_groupi_n_9850, csa_tree_add_51_79_groupi_n_9851, csa_tree_add_51_79_groupi_n_9852, csa_tree_add_51_79_groupi_n_9853, csa_tree_add_51_79_groupi_n_9854, csa_tree_add_51_79_groupi_n_9855, csa_tree_add_51_79_groupi_n_9856;
  wire csa_tree_add_51_79_groupi_n_9857, csa_tree_add_51_79_groupi_n_9858, csa_tree_add_51_79_groupi_n_9859, csa_tree_add_51_79_groupi_n_9860, csa_tree_add_51_79_groupi_n_9861, csa_tree_add_51_79_groupi_n_9862, csa_tree_add_51_79_groupi_n_9863, csa_tree_add_51_79_groupi_n_9864;
  wire csa_tree_add_51_79_groupi_n_9865, csa_tree_add_51_79_groupi_n_9866, csa_tree_add_51_79_groupi_n_9867, csa_tree_add_51_79_groupi_n_9868, csa_tree_add_51_79_groupi_n_9869, csa_tree_add_51_79_groupi_n_9870, csa_tree_add_51_79_groupi_n_9871, csa_tree_add_51_79_groupi_n_9872;
  wire csa_tree_add_51_79_groupi_n_9873, csa_tree_add_51_79_groupi_n_9874, csa_tree_add_51_79_groupi_n_9875, csa_tree_add_51_79_groupi_n_9876, csa_tree_add_51_79_groupi_n_9877, csa_tree_add_51_79_groupi_n_9878, csa_tree_add_51_79_groupi_n_9879, csa_tree_add_51_79_groupi_n_9880;
  wire csa_tree_add_51_79_groupi_n_9881, csa_tree_add_51_79_groupi_n_9882, csa_tree_add_51_79_groupi_n_9883, csa_tree_add_51_79_groupi_n_9884, csa_tree_add_51_79_groupi_n_9885, csa_tree_add_51_79_groupi_n_9886, csa_tree_add_51_79_groupi_n_9887, csa_tree_add_51_79_groupi_n_9888;
  wire csa_tree_add_51_79_groupi_n_9889, csa_tree_add_51_79_groupi_n_9890, csa_tree_add_51_79_groupi_n_9891, csa_tree_add_51_79_groupi_n_9892, csa_tree_add_51_79_groupi_n_9893, csa_tree_add_51_79_groupi_n_9894, csa_tree_add_51_79_groupi_n_9895, csa_tree_add_51_79_groupi_n_9896;
  wire csa_tree_add_51_79_groupi_n_9897, csa_tree_add_51_79_groupi_n_9898, csa_tree_add_51_79_groupi_n_9899, csa_tree_add_51_79_groupi_n_9900, csa_tree_add_51_79_groupi_n_9901, csa_tree_add_51_79_groupi_n_9902, csa_tree_add_51_79_groupi_n_9903, csa_tree_add_51_79_groupi_n_9904;
  wire csa_tree_add_51_79_groupi_n_9905, csa_tree_add_51_79_groupi_n_9906, csa_tree_add_51_79_groupi_n_9907, csa_tree_add_51_79_groupi_n_9908, csa_tree_add_51_79_groupi_n_9909, csa_tree_add_51_79_groupi_n_9910, csa_tree_add_51_79_groupi_n_9911, csa_tree_add_51_79_groupi_n_9912;
  wire csa_tree_add_51_79_groupi_n_9913, csa_tree_add_51_79_groupi_n_9914, csa_tree_add_51_79_groupi_n_9915, csa_tree_add_51_79_groupi_n_9916, csa_tree_add_51_79_groupi_n_9917, csa_tree_add_51_79_groupi_n_9918, csa_tree_add_51_79_groupi_n_9919, csa_tree_add_51_79_groupi_n_9920;
  wire csa_tree_add_51_79_groupi_n_9921, csa_tree_add_51_79_groupi_n_9922, csa_tree_add_51_79_groupi_n_9923, csa_tree_add_51_79_groupi_n_9924, csa_tree_add_51_79_groupi_n_9925, csa_tree_add_51_79_groupi_n_9926, csa_tree_add_51_79_groupi_n_9927, csa_tree_add_51_79_groupi_n_9928;
  wire csa_tree_add_51_79_groupi_n_9929, csa_tree_add_51_79_groupi_n_9930, csa_tree_add_51_79_groupi_n_9931, csa_tree_add_51_79_groupi_n_9932, csa_tree_add_51_79_groupi_n_9933, csa_tree_add_51_79_groupi_n_9934, csa_tree_add_51_79_groupi_n_9935, csa_tree_add_51_79_groupi_n_9936;
  wire csa_tree_add_51_79_groupi_n_9937, csa_tree_add_51_79_groupi_n_9938, csa_tree_add_51_79_groupi_n_9939, csa_tree_add_51_79_groupi_n_9940, csa_tree_add_51_79_groupi_n_9941, csa_tree_add_51_79_groupi_n_9942, csa_tree_add_51_79_groupi_n_9943, csa_tree_add_51_79_groupi_n_9944;
  wire csa_tree_add_51_79_groupi_n_9945, csa_tree_add_51_79_groupi_n_9946, csa_tree_add_51_79_groupi_n_9947, csa_tree_add_51_79_groupi_n_9948, csa_tree_add_51_79_groupi_n_9949, csa_tree_add_51_79_groupi_n_9950, csa_tree_add_51_79_groupi_n_9951, csa_tree_add_51_79_groupi_n_9952;
  wire csa_tree_add_51_79_groupi_n_9953, csa_tree_add_51_79_groupi_n_9954, csa_tree_add_51_79_groupi_n_9955, csa_tree_add_51_79_groupi_n_9956, csa_tree_add_51_79_groupi_n_9957, csa_tree_add_51_79_groupi_n_9958, csa_tree_add_51_79_groupi_n_9959, csa_tree_add_51_79_groupi_n_9960;
  wire csa_tree_add_51_79_groupi_n_9961, csa_tree_add_51_79_groupi_n_9962, csa_tree_add_51_79_groupi_n_9963, csa_tree_add_51_79_groupi_n_9964, csa_tree_add_51_79_groupi_n_9966, csa_tree_add_51_79_groupi_n_9967, csa_tree_add_51_79_groupi_n_9968, csa_tree_add_51_79_groupi_n_9969;
  wire csa_tree_add_51_79_groupi_n_9970, csa_tree_add_51_79_groupi_n_9971, csa_tree_add_51_79_groupi_n_9972, csa_tree_add_51_79_groupi_n_9973, csa_tree_add_51_79_groupi_n_9974, csa_tree_add_51_79_groupi_n_9975, csa_tree_add_51_79_groupi_n_9976, csa_tree_add_51_79_groupi_n_9977;
  wire csa_tree_add_51_79_groupi_n_9978, csa_tree_add_51_79_groupi_n_9979, csa_tree_add_51_79_groupi_n_9980, csa_tree_add_51_79_groupi_n_9981, csa_tree_add_51_79_groupi_n_9982, csa_tree_add_51_79_groupi_n_9983, csa_tree_add_51_79_groupi_n_9984, csa_tree_add_51_79_groupi_n_9985;
  wire csa_tree_add_51_79_groupi_n_9986, csa_tree_add_51_79_groupi_n_9987, csa_tree_add_51_79_groupi_n_9988, csa_tree_add_51_79_groupi_n_9989, csa_tree_add_51_79_groupi_n_9990, csa_tree_add_51_79_groupi_n_9991, csa_tree_add_51_79_groupi_n_9992, csa_tree_add_51_79_groupi_n_9993;
  wire csa_tree_add_51_79_groupi_n_9994, csa_tree_add_51_79_groupi_n_9995, csa_tree_add_51_79_groupi_n_9996, csa_tree_add_51_79_groupi_n_9997, csa_tree_add_51_79_groupi_n_9998, csa_tree_add_51_79_groupi_n_9999, csa_tree_add_51_79_groupi_n_10000, csa_tree_add_51_79_groupi_n_10001;
  wire csa_tree_add_51_79_groupi_n_10002, csa_tree_add_51_79_groupi_n_10003, csa_tree_add_51_79_groupi_n_10004, csa_tree_add_51_79_groupi_n_10005, csa_tree_add_51_79_groupi_n_10006, csa_tree_add_51_79_groupi_n_10007, csa_tree_add_51_79_groupi_n_10008, csa_tree_add_51_79_groupi_n_10009;
  wire csa_tree_add_51_79_groupi_n_10010, csa_tree_add_51_79_groupi_n_10011, csa_tree_add_51_79_groupi_n_10012, csa_tree_add_51_79_groupi_n_10013, csa_tree_add_51_79_groupi_n_10014, csa_tree_add_51_79_groupi_n_10015, csa_tree_add_51_79_groupi_n_10016, csa_tree_add_51_79_groupi_n_10017;
  wire csa_tree_add_51_79_groupi_n_10018, csa_tree_add_51_79_groupi_n_10019, csa_tree_add_51_79_groupi_n_10020, csa_tree_add_51_79_groupi_n_10021, csa_tree_add_51_79_groupi_n_10022, csa_tree_add_51_79_groupi_n_10023, csa_tree_add_51_79_groupi_n_10024, csa_tree_add_51_79_groupi_n_10025;
  wire csa_tree_add_51_79_groupi_n_10026, csa_tree_add_51_79_groupi_n_10027, csa_tree_add_51_79_groupi_n_10028, csa_tree_add_51_79_groupi_n_10029, csa_tree_add_51_79_groupi_n_10030, csa_tree_add_51_79_groupi_n_10031, csa_tree_add_51_79_groupi_n_10032, csa_tree_add_51_79_groupi_n_10033;
  wire csa_tree_add_51_79_groupi_n_10034, csa_tree_add_51_79_groupi_n_10035, csa_tree_add_51_79_groupi_n_10036, csa_tree_add_51_79_groupi_n_10037, csa_tree_add_51_79_groupi_n_10038, csa_tree_add_51_79_groupi_n_10039, csa_tree_add_51_79_groupi_n_10040, csa_tree_add_51_79_groupi_n_10041;
  wire csa_tree_add_51_79_groupi_n_10042, csa_tree_add_51_79_groupi_n_10043, csa_tree_add_51_79_groupi_n_10044, csa_tree_add_51_79_groupi_n_10045, csa_tree_add_51_79_groupi_n_10046, csa_tree_add_51_79_groupi_n_10047, csa_tree_add_51_79_groupi_n_10048, csa_tree_add_51_79_groupi_n_10049;
  wire csa_tree_add_51_79_groupi_n_10050, csa_tree_add_51_79_groupi_n_10051, csa_tree_add_51_79_groupi_n_10052, csa_tree_add_51_79_groupi_n_10053, csa_tree_add_51_79_groupi_n_10054, csa_tree_add_51_79_groupi_n_10055, csa_tree_add_51_79_groupi_n_10056, csa_tree_add_51_79_groupi_n_10057;
  wire csa_tree_add_51_79_groupi_n_10058, csa_tree_add_51_79_groupi_n_10059, csa_tree_add_51_79_groupi_n_10060, csa_tree_add_51_79_groupi_n_10061, csa_tree_add_51_79_groupi_n_10062, csa_tree_add_51_79_groupi_n_10063, csa_tree_add_51_79_groupi_n_10064, csa_tree_add_51_79_groupi_n_10065;
  wire csa_tree_add_51_79_groupi_n_10066, csa_tree_add_51_79_groupi_n_10067, csa_tree_add_51_79_groupi_n_10068, csa_tree_add_51_79_groupi_n_10069, csa_tree_add_51_79_groupi_n_10070, csa_tree_add_51_79_groupi_n_10071, csa_tree_add_51_79_groupi_n_10072, csa_tree_add_51_79_groupi_n_10073;
  wire csa_tree_add_51_79_groupi_n_10074, csa_tree_add_51_79_groupi_n_10075, csa_tree_add_51_79_groupi_n_10076, csa_tree_add_51_79_groupi_n_10077, csa_tree_add_51_79_groupi_n_10078, csa_tree_add_51_79_groupi_n_10079, csa_tree_add_51_79_groupi_n_10080, csa_tree_add_51_79_groupi_n_10081;
  wire csa_tree_add_51_79_groupi_n_10082, csa_tree_add_51_79_groupi_n_10083, csa_tree_add_51_79_groupi_n_10084, csa_tree_add_51_79_groupi_n_10085, csa_tree_add_51_79_groupi_n_10086, csa_tree_add_51_79_groupi_n_10087, csa_tree_add_51_79_groupi_n_10088, csa_tree_add_51_79_groupi_n_10089;
  wire csa_tree_add_51_79_groupi_n_10090, csa_tree_add_51_79_groupi_n_10091, csa_tree_add_51_79_groupi_n_10092, csa_tree_add_51_79_groupi_n_10093, csa_tree_add_51_79_groupi_n_10094, csa_tree_add_51_79_groupi_n_10095, csa_tree_add_51_79_groupi_n_10096, csa_tree_add_51_79_groupi_n_10097;
  wire csa_tree_add_51_79_groupi_n_10098, csa_tree_add_51_79_groupi_n_10099, csa_tree_add_51_79_groupi_n_10100, csa_tree_add_51_79_groupi_n_10101, csa_tree_add_51_79_groupi_n_10102, csa_tree_add_51_79_groupi_n_10103, csa_tree_add_51_79_groupi_n_10104, csa_tree_add_51_79_groupi_n_10105;
  wire csa_tree_add_51_79_groupi_n_10106, csa_tree_add_51_79_groupi_n_10107, csa_tree_add_51_79_groupi_n_10108, csa_tree_add_51_79_groupi_n_10109, csa_tree_add_51_79_groupi_n_10110, csa_tree_add_51_79_groupi_n_10111, csa_tree_add_51_79_groupi_n_10112, csa_tree_add_51_79_groupi_n_10113;
  wire csa_tree_add_51_79_groupi_n_10114, csa_tree_add_51_79_groupi_n_10115, csa_tree_add_51_79_groupi_n_10116, csa_tree_add_51_79_groupi_n_10117, csa_tree_add_51_79_groupi_n_10118, csa_tree_add_51_79_groupi_n_10119, csa_tree_add_51_79_groupi_n_10120, csa_tree_add_51_79_groupi_n_10121;
  wire csa_tree_add_51_79_groupi_n_10122, csa_tree_add_51_79_groupi_n_10123, csa_tree_add_51_79_groupi_n_10124, csa_tree_add_51_79_groupi_n_10125, csa_tree_add_51_79_groupi_n_10126, csa_tree_add_51_79_groupi_n_10127, csa_tree_add_51_79_groupi_n_10128, csa_tree_add_51_79_groupi_n_10129;
  wire csa_tree_add_51_79_groupi_n_10130, csa_tree_add_51_79_groupi_n_10131, csa_tree_add_51_79_groupi_n_10132, csa_tree_add_51_79_groupi_n_10133, csa_tree_add_51_79_groupi_n_10134, csa_tree_add_51_79_groupi_n_10135, csa_tree_add_51_79_groupi_n_10136, csa_tree_add_51_79_groupi_n_10137;
  wire csa_tree_add_51_79_groupi_n_10138, csa_tree_add_51_79_groupi_n_10139, csa_tree_add_51_79_groupi_n_10140, csa_tree_add_51_79_groupi_n_10141, csa_tree_add_51_79_groupi_n_10142, csa_tree_add_51_79_groupi_n_10143, csa_tree_add_51_79_groupi_n_10144, csa_tree_add_51_79_groupi_n_10145;
  wire csa_tree_add_51_79_groupi_n_10146, csa_tree_add_51_79_groupi_n_10147, csa_tree_add_51_79_groupi_n_10148, csa_tree_add_51_79_groupi_n_10149, csa_tree_add_51_79_groupi_n_10150, csa_tree_add_51_79_groupi_n_10151, csa_tree_add_51_79_groupi_n_10152, csa_tree_add_51_79_groupi_n_10153;
  wire csa_tree_add_51_79_groupi_n_10154, csa_tree_add_51_79_groupi_n_10155, csa_tree_add_51_79_groupi_n_10156, csa_tree_add_51_79_groupi_n_10157, csa_tree_add_51_79_groupi_n_10158, csa_tree_add_51_79_groupi_n_10159, csa_tree_add_51_79_groupi_n_10160, csa_tree_add_51_79_groupi_n_10161;
  wire csa_tree_add_51_79_groupi_n_10162, csa_tree_add_51_79_groupi_n_10163, csa_tree_add_51_79_groupi_n_10164, csa_tree_add_51_79_groupi_n_10165, csa_tree_add_51_79_groupi_n_10166, csa_tree_add_51_79_groupi_n_10167, csa_tree_add_51_79_groupi_n_10168, csa_tree_add_51_79_groupi_n_10169;
  wire csa_tree_add_51_79_groupi_n_10170, csa_tree_add_51_79_groupi_n_10171, csa_tree_add_51_79_groupi_n_10172, csa_tree_add_51_79_groupi_n_10173, csa_tree_add_51_79_groupi_n_10174, csa_tree_add_51_79_groupi_n_10175, csa_tree_add_51_79_groupi_n_10176, csa_tree_add_51_79_groupi_n_10177;
  wire csa_tree_add_51_79_groupi_n_10178, csa_tree_add_51_79_groupi_n_10179, csa_tree_add_51_79_groupi_n_10180, csa_tree_add_51_79_groupi_n_10181, csa_tree_add_51_79_groupi_n_10182, csa_tree_add_51_79_groupi_n_10183, csa_tree_add_51_79_groupi_n_10184, csa_tree_add_51_79_groupi_n_10185;
  wire csa_tree_add_51_79_groupi_n_10186, csa_tree_add_51_79_groupi_n_10187, csa_tree_add_51_79_groupi_n_10188, csa_tree_add_51_79_groupi_n_10189, csa_tree_add_51_79_groupi_n_10190, csa_tree_add_51_79_groupi_n_10191, csa_tree_add_51_79_groupi_n_10192, csa_tree_add_51_79_groupi_n_10193;
  wire csa_tree_add_51_79_groupi_n_10194, csa_tree_add_51_79_groupi_n_10195, csa_tree_add_51_79_groupi_n_10196, csa_tree_add_51_79_groupi_n_10197, csa_tree_add_51_79_groupi_n_10198, csa_tree_add_51_79_groupi_n_10199, csa_tree_add_51_79_groupi_n_10200, csa_tree_add_51_79_groupi_n_10201;
  wire csa_tree_add_51_79_groupi_n_10202, csa_tree_add_51_79_groupi_n_10203, csa_tree_add_51_79_groupi_n_10204, csa_tree_add_51_79_groupi_n_10205, csa_tree_add_51_79_groupi_n_10206, csa_tree_add_51_79_groupi_n_10207, csa_tree_add_51_79_groupi_n_10208, csa_tree_add_51_79_groupi_n_10209;
  wire csa_tree_add_51_79_groupi_n_10210, csa_tree_add_51_79_groupi_n_10211, csa_tree_add_51_79_groupi_n_10212, csa_tree_add_51_79_groupi_n_10213, csa_tree_add_51_79_groupi_n_10214, csa_tree_add_51_79_groupi_n_10215, csa_tree_add_51_79_groupi_n_10216, csa_tree_add_51_79_groupi_n_10217;
  wire csa_tree_add_51_79_groupi_n_10218, csa_tree_add_51_79_groupi_n_10219, csa_tree_add_51_79_groupi_n_10220, csa_tree_add_51_79_groupi_n_10221, csa_tree_add_51_79_groupi_n_10222, csa_tree_add_51_79_groupi_n_10223, csa_tree_add_51_79_groupi_n_10224, csa_tree_add_51_79_groupi_n_10225;
  wire csa_tree_add_51_79_groupi_n_10226, csa_tree_add_51_79_groupi_n_10227, csa_tree_add_51_79_groupi_n_10228, csa_tree_add_51_79_groupi_n_10229, csa_tree_add_51_79_groupi_n_10230, csa_tree_add_51_79_groupi_n_10231, csa_tree_add_51_79_groupi_n_10232, csa_tree_add_51_79_groupi_n_10233;
  wire csa_tree_add_51_79_groupi_n_10234, csa_tree_add_51_79_groupi_n_10235, csa_tree_add_51_79_groupi_n_10236, csa_tree_add_51_79_groupi_n_10237, csa_tree_add_51_79_groupi_n_10238, csa_tree_add_51_79_groupi_n_10239, csa_tree_add_51_79_groupi_n_10240, csa_tree_add_51_79_groupi_n_10241;
  wire csa_tree_add_51_79_groupi_n_10242, csa_tree_add_51_79_groupi_n_10243, csa_tree_add_51_79_groupi_n_10244, csa_tree_add_51_79_groupi_n_10245, csa_tree_add_51_79_groupi_n_10246, csa_tree_add_51_79_groupi_n_10247, csa_tree_add_51_79_groupi_n_10248, csa_tree_add_51_79_groupi_n_10249;
  wire csa_tree_add_51_79_groupi_n_10250, csa_tree_add_51_79_groupi_n_10251, csa_tree_add_51_79_groupi_n_10252, csa_tree_add_51_79_groupi_n_10253, csa_tree_add_51_79_groupi_n_10254, csa_tree_add_51_79_groupi_n_10255, csa_tree_add_51_79_groupi_n_10256, csa_tree_add_51_79_groupi_n_10257;
  wire csa_tree_add_51_79_groupi_n_10258, csa_tree_add_51_79_groupi_n_10259, csa_tree_add_51_79_groupi_n_10260, csa_tree_add_51_79_groupi_n_10261, csa_tree_add_51_79_groupi_n_10262, csa_tree_add_51_79_groupi_n_10263, csa_tree_add_51_79_groupi_n_10264, csa_tree_add_51_79_groupi_n_10265;
  wire csa_tree_add_51_79_groupi_n_10266, csa_tree_add_51_79_groupi_n_10267, csa_tree_add_51_79_groupi_n_10268, csa_tree_add_51_79_groupi_n_10269, csa_tree_add_51_79_groupi_n_10270, csa_tree_add_51_79_groupi_n_10271, csa_tree_add_51_79_groupi_n_10272, csa_tree_add_51_79_groupi_n_10273;
  wire csa_tree_add_51_79_groupi_n_10274, csa_tree_add_51_79_groupi_n_10275, csa_tree_add_51_79_groupi_n_10276, csa_tree_add_51_79_groupi_n_10277, csa_tree_add_51_79_groupi_n_10278, csa_tree_add_51_79_groupi_n_10279, csa_tree_add_51_79_groupi_n_10280, csa_tree_add_51_79_groupi_n_10281;
  wire csa_tree_add_51_79_groupi_n_10282, csa_tree_add_51_79_groupi_n_10283, csa_tree_add_51_79_groupi_n_10284, csa_tree_add_51_79_groupi_n_10285, csa_tree_add_51_79_groupi_n_10286, csa_tree_add_51_79_groupi_n_10287, csa_tree_add_51_79_groupi_n_10288, csa_tree_add_51_79_groupi_n_10289;
  wire csa_tree_add_51_79_groupi_n_10290, csa_tree_add_51_79_groupi_n_10291, csa_tree_add_51_79_groupi_n_10292, csa_tree_add_51_79_groupi_n_10293, csa_tree_add_51_79_groupi_n_10294, csa_tree_add_51_79_groupi_n_10295, csa_tree_add_51_79_groupi_n_10296, csa_tree_add_51_79_groupi_n_10297;
  wire csa_tree_add_51_79_groupi_n_10298, csa_tree_add_51_79_groupi_n_10299, csa_tree_add_51_79_groupi_n_10300, csa_tree_add_51_79_groupi_n_10301, csa_tree_add_51_79_groupi_n_10302, csa_tree_add_51_79_groupi_n_10303, csa_tree_add_51_79_groupi_n_10304, csa_tree_add_51_79_groupi_n_10305;
  wire csa_tree_add_51_79_groupi_n_10306, csa_tree_add_51_79_groupi_n_10307, csa_tree_add_51_79_groupi_n_10308, csa_tree_add_51_79_groupi_n_10309, csa_tree_add_51_79_groupi_n_10310, csa_tree_add_51_79_groupi_n_10311, csa_tree_add_51_79_groupi_n_10312, csa_tree_add_51_79_groupi_n_10313;
  wire csa_tree_add_51_79_groupi_n_10314, csa_tree_add_51_79_groupi_n_10315, csa_tree_add_51_79_groupi_n_10316, csa_tree_add_51_79_groupi_n_10317, csa_tree_add_51_79_groupi_n_10318, csa_tree_add_51_79_groupi_n_10319, csa_tree_add_51_79_groupi_n_10320, csa_tree_add_51_79_groupi_n_10321;
  wire csa_tree_add_51_79_groupi_n_10322, csa_tree_add_51_79_groupi_n_10323, csa_tree_add_51_79_groupi_n_10324, csa_tree_add_51_79_groupi_n_10325, csa_tree_add_51_79_groupi_n_10326, csa_tree_add_51_79_groupi_n_10327, csa_tree_add_51_79_groupi_n_10328, csa_tree_add_51_79_groupi_n_10329;
  wire csa_tree_add_51_79_groupi_n_10330, csa_tree_add_51_79_groupi_n_10331, csa_tree_add_51_79_groupi_n_10332, csa_tree_add_51_79_groupi_n_10333, csa_tree_add_51_79_groupi_n_10334, csa_tree_add_51_79_groupi_n_10335, csa_tree_add_51_79_groupi_n_10336, csa_tree_add_51_79_groupi_n_10337;
  wire csa_tree_add_51_79_groupi_n_10338, csa_tree_add_51_79_groupi_n_10339, csa_tree_add_51_79_groupi_n_10340, csa_tree_add_51_79_groupi_n_10341, csa_tree_add_51_79_groupi_n_10342, csa_tree_add_51_79_groupi_n_10343, csa_tree_add_51_79_groupi_n_10344, csa_tree_add_51_79_groupi_n_10345;
  wire csa_tree_add_51_79_groupi_n_10346, csa_tree_add_51_79_groupi_n_10347, csa_tree_add_51_79_groupi_n_10348, csa_tree_add_51_79_groupi_n_10349, csa_tree_add_51_79_groupi_n_10350, csa_tree_add_51_79_groupi_n_10351, csa_tree_add_51_79_groupi_n_10352, csa_tree_add_51_79_groupi_n_10353;
  wire csa_tree_add_51_79_groupi_n_10354, csa_tree_add_51_79_groupi_n_10355, csa_tree_add_51_79_groupi_n_10356, csa_tree_add_51_79_groupi_n_10357, csa_tree_add_51_79_groupi_n_10358, csa_tree_add_51_79_groupi_n_10359, csa_tree_add_51_79_groupi_n_10360, csa_tree_add_51_79_groupi_n_10361;
  wire csa_tree_add_51_79_groupi_n_10362, csa_tree_add_51_79_groupi_n_10363, csa_tree_add_51_79_groupi_n_10364, csa_tree_add_51_79_groupi_n_10365, csa_tree_add_51_79_groupi_n_10366, csa_tree_add_51_79_groupi_n_10367, csa_tree_add_51_79_groupi_n_10368, csa_tree_add_51_79_groupi_n_10369;
  wire csa_tree_add_51_79_groupi_n_10370, csa_tree_add_51_79_groupi_n_10371, csa_tree_add_51_79_groupi_n_10372, csa_tree_add_51_79_groupi_n_10373, csa_tree_add_51_79_groupi_n_10374, csa_tree_add_51_79_groupi_n_10375, csa_tree_add_51_79_groupi_n_10376, csa_tree_add_51_79_groupi_n_10377;
  wire csa_tree_add_51_79_groupi_n_10378, csa_tree_add_51_79_groupi_n_10379, csa_tree_add_51_79_groupi_n_10380, csa_tree_add_51_79_groupi_n_10381, csa_tree_add_51_79_groupi_n_10382, csa_tree_add_51_79_groupi_n_10383, csa_tree_add_51_79_groupi_n_10384, csa_tree_add_51_79_groupi_n_10385;
  wire csa_tree_add_51_79_groupi_n_10386, csa_tree_add_51_79_groupi_n_10387, csa_tree_add_51_79_groupi_n_10388, csa_tree_add_51_79_groupi_n_10389, csa_tree_add_51_79_groupi_n_10390, csa_tree_add_51_79_groupi_n_10391, csa_tree_add_51_79_groupi_n_10392, csa_tree_add_51_79_groupi_n_10393;
  wire csa_tree_add_51_79_groupi_n_10394, csa_tree_add_51_79_groupi_n_10395, csa_tree_add_51_79_groupi_n_10396, csa_tree_add_51_79_groupi_n_10397, csa_tree_add_51_79_groupi_n_10398, csa_tree_add_51_79_groupi_n_10399, csa_tree_add_51_79_groupi_n_10400, csa_tree_add_51_79_groupi_n_10401;
  wire csa_tree_add_51_79_groupi_n_10402, csa_tree_add_51_79_groupi_n_10403, csa_tree_add_51_79_groupi_n_10404, csa_tree_add_51_79_groupi_n_10405, csa_tree_add_51_79_groupi_n_10406, csa_tree_add_51_79_groupi_n_10407, csa_tree_add_51_79_groupi_n_10408, csa_tree_add_51_79_groupi_n_10409;
  wire csa_tree_add_51_79_groupi_n_10410, csa_tree_add_51_79_groupi_n_10411, csa_tree_add_51_79_groupi_n_10412, csa_tree_add_51_79_groupi_n_10413, csa_tree_add_51_79_groupi_n_10414, csa_tree_add_51_79_groupi_n_10415, csa_tree_add_51_79_groupi_n_10416, csa_tree_add_51_79_groupi_n_10417;
  wire csa_tree_add_51_79_groupi_n_10418, csa_tree_add_51_79_groupi_n_10419, csa_tree_add_51_79_groupi_n_10420, csa_tree_add_51_79_groupi_n_10421, csa_tree_add_51_79_groupi_n_10422, csa_tree_add_51_79_groupi_n_10423, csa_tree_add_51_79_groupi_n_10424, csa_tree_add_51_79_groupi_n_10425;
  wire csa_tree_add_51_79_groupi_n_10426, csa_tree_add_51_79_groupi_n_10427, csa_tree_add_51_79_groupi_n_10428, csa_tree_add_51_79_groupi_n_10429, csa_tree_add_51_79_groupi_n_10430, csa_tree_add_51_79_groupi_n_10431, csa_tree_add_51_79_groupi_n_10432, csa_tree_add_51_79_groupi_n_10433;
  wire csa_tree_add_51_79_groupi_n_10434, csa_tree_add_51_79_groupi_n_10435, csa_tree_add_51_79_groupi_n_10436, csa_tree_add_51_79_groupi_n_10437, csa_tree_add_51_79_groupi_n_10438, csa_tree_add_51_79_groupi_n_10439, csa_tree_add_51_79_groupi_n_10440, csa_tree_add_51_79_groupi_n_10441;
  wire csa_tree_add_51_79_groupi_n_10442, csa_tree_add_51_79_groupi_n_10443, csa_tree_add_51_79_groupi_n_10444, csa_tree_add_51_79_groupi_n_10445, csa_tree_add_51_79_groupi_n_10446, csa_tree_add_51_79_groupi_n_10447, csa_tree_add_51_79_groupi_n_10448, csa_tree_add_51_79_groupi_n_10449;
  wire csa_tree_add_51_79_groupi_n_10451, csa_tree_add_51_79_groupi_n_10452, csa_tree_add_51_79_groupi_n_10453, csa_tree_add_51_79_groupi_n_10454, csa_tree_add_51_79_groupi_n_10455, csa_tree_add_51_79_groupi_n_10456, csa_tree_add_51_79_groupi_n_10457, csa_tree_add_51_79_groupi_n_10458;
  wire csa_tree_add_51_79_groupi_n_10459, csa_tree_add_51_79_groupi_n_10460, csa_tree_add_51_79_groupi_n_10461, csa_tree_add_51_79_groupi_n_10462, csa_tree_add_51_79_groupi_n_10463, csa_tree_add_51_79_groupi_n_10464, csa_tree_add_51_79_groupi_n_10465, csa_tree_add_51_79_groupi_n_10466;
  wire csa_tree_add_51_79_groupi_n_10467, csa_tree_add_51_79_groupi_n_10468, csa_tree_add_51_79_groupi_n_10469, csa_tree_add_51_79_groupi_n_10470, csa_tree_add_51_79_groupi_n_10471, csa_tree_add_51_79_groupi_n_10472, csa_tree_add_51_79_groupi_n_10473, csa_tree_add_51_79_groupi_n_10474;
  wire csa_tree_add_51_79_groupi_n_10475, csa_tree_add_51_79_groupi_n_10476, csa_tree_add_51_79_groupi_n_10477, csa_tree_add_51_79_groupi_n_10478, csa_tree_add_51_79_groupi_n_10479, csa_tree_add_51_79_groupi_n_10480, csa_tree_add_51_79_groupi_n_10481, csa_tree_add_51_79_groupi_n_10482;
  wire csa_tree_add_51_79_groupi_n_10483, csa_tree_add_51_79_groupi_n_10484, csa_tree_add_51_79_groupi_n_10485, csa_tree_add_51_79_groupi_n_10486, csa_tree_add_51_79_groupi_n_10487, csa_tree_add_51_79_groupi_n_10488, csa_tree_add_51_79_groupi_n_10489, csa_tree_add_51_79_groupi_n_10490;
  wire csa_tree_add_51_79_groupi_n_10491, csa_tree_add_51_79_groupi_n_10492, csa_tree_add_51_79_groupi_n_10493, csa_tree_add_51_79_groupi_n_10494, csa_tree_add_51_79_groupi_n_10495, csa_tree_add_51_79_groupi_n_10496, csa_tree_add_51_79_groupi_n_10497, csa_tree_add_51_79_groupi_n_10498;
  wire csa_tree_add_51_79_groupi_n_10499, csa_tree_add_51_79_groupi_n_10500, csa_tree_add_51_79_groupi_n_10501, csa_tree_add_51_79_groupi_n_10502, csa_tree_add_51_79_groupi_n_10503, csa_tree_add_51_79_groupi_n_10504, csa_tree_add_51_79_groupi_n_10505, csa_tree_add_51_79_groupi_n_10506;
  wire csa_tree_add_51_79_groupi_n_10507, csa_tree_add_51_79_groupi_n_10508, csa_tree_add_51_79_groupi_n_10509, csa_tree_add_51_79_groupi_n_10510, csa_tree_add_51_79_groupi_n_10511, csa_tree_add_51_79_groupi_n_10512, csa_tree_add_51_79_groupi_n_10513, csa_tree_add_51_79_groupi_n_10514;
  wire csa_tree_add_51_79_groupi_n_10515, csa_tree_add_51_79_groupi_n_10516, csa_tree_add_51_79_groupi_n_10517, csa_tree_add_51_79_groupi_n_10518, csa_tree_add_51_79_groupi_n_10519, csa_tree_add_51_79_groupi_n_10520, csa_tree_add_51_79_groupi_n_10521, csa_tree_add_51_79_groupi_n_10522;
  wire csa_tree_add_51_79_groupi_n_10523, csa_tree_add_51_79_groupi_n_10524, csa_tree_add_51_79_groupi_n_10525, csa_tree_add_51_79_groupi_n_10526, csa_tree_add_51_79_groupi_n_10527, csa_tree_add_51_79_groupi_n_10528, csa_tree_add_51_79_groupi_n_10529, csa_tree_add_51_79_groupi_n_10530;
  wire csa_tree_add_51_79_groupi_n_10531, csa_tree_add_51_79_groupi_n_10532, csa_tree_add_51_79_groupi_n_10533, csa_tree_add_51_79_groupi_n_10534, csa_tree_add_51_79_groupi_n_10535, csa_tree_add_51_79_groupi_n_10536, csa_tree_add_51_79_groupi_n_10537, csa_tree_add_51_79_groupi_n_10538;
  wire csa_tree_add_51_79_groupi_n_10539, csa_tree_add_51_79_groupi_n_10540, csa_tree_add_51_79_groupi_n_10541, csa_tree_add_51_79_groupi_n_10542, csa_tree_add_51_79_groupi_n_10543, csa_tree_add_51_79_groupi_n_10544, csa_tree_add_51_79_groupi_n_10545, csa_tree_add_51_79_groupi_n_10546;
  wire csa_tree_add_51_79_groupi_n_10547, csa_tree_add_51_79_groupi_n_10548, csa_tree_add_51_79_groupi_n_10549, csa_tree_add_51_79_groupi_n_10550, csa_tree_add_51_79_groupi_n_10551, csa_tree_add_51_79_groupi_n_10552, csa_tree_add_51_79_groupi_n_10553, csa_tree_add_51_79_groupi_n_10554;
  wire csa_tree_add_51_79_groupi_n_10555, csa_tree_add_51_79_groupi_n_10556, csa_tree_add_51_79_groupi_n_10557, csa_tree_add_51_79_groupi_n_10558, csa_tree_add_51_79_groupi_n_10559, csa_tree_add_51_79_groupi_n_10560, csa_tree_add_51_79_groupi_n_10561, csa_tree_add_51_79_groupi_n_10562;
  wire csa_tree_add_51_79_groupi_n_10563, csa_tree_add_51_79_groupi_n_10564, csa_tree_add_51_79_groupi_n_10565, csa_tree_add_51_79_groupi_n_10566, csa_tree_add_51_79_groupi_n_10567, csa_tree_add_51_79_groupi_n_10568, csa_tree_add_51_79_groupi_n_10569, csa_tree_add_51_79_groupi_n_10570;
  wire csa_tree_add_51_79_groupi_n_10571, csa_tree_add_51_79_groupi_n_10572, csa_tree_add_51_79_groupi_n_10573, csa_tree_add_51_79_groupi_n_10574, csa_tree_add_51_79_groupi_n_10575, csa_tree_add_51_79_groupi_n_10576, csa_tree_add_51_79_groupi_n_10577, csa_tree_add_51_79_groupi_n_10578;
  wire csa_tree_add_51_79_groupi_n_10579, csa_tree_add_51_79_groupi_n_10580, csa_tree_add_51_79_groupi_n_10581, csa_tree_add_51_79_groupi_n_10582, csa_tree_add_51_79_groupi_n_10583, csa_tree_add_51_79_groupi_n_10584, csa_tree_add_51_79_groupi_n_10585, csa_tree_add_51_79_groupi_n_10586;
  wire csa_tree_add_51_79_groupi_n_10587, csa_tree_add_51_79_groupi_n_10588, csa_tree_add_51_79_groupi_n_10589, csa_tree_add_51_79_groupi_n_10590, csa_tree_add_51_79_groupi_n_10591, csa_tree_add_51_79_groupi_n_10592, csa_tree_add_51_79_groupi_n_10593, csa_tree_add_51_79_groupi_n_10594;
  wire csa_tree_add_51_79_groupi_n_10595, csa_tree_add_51_79_groupi_n_10596, csa_tree_add_51_79_groupi_n_10597, csa_tree_add_51_79_groupi_n_10598, csa_tree_add_51_79_groupi_n_10599, csa_tree_add_51_79_groupi_n_10600, csa_tree_add_51_79_groupi_n_10601, csa_tree_add_51_79_groupi_n_10602;
  wire csa_tree_add_51_79_groupi_n_10603, csa_tree_add_51_79_groupi_n_10604, csa_tree_add_51_79_groupi_n_10605, csa_tree_add_51_79_groupi_n_10606, csa_tree_add_51_79_groupi_n_10607, csa_tree_add_51_79_groupi_n_10608, csa_tree_add_51_79_groupi_n_10609, csa_tree_add_51_79_groupi_n_10610;
  wire csa_tree_add_51_79_groupi_n_10611, csa_tree_add_51_79_groupi_n_10612, csa_tree_add_51_79_groupi_n_10613, csa_tree_add_51_79_groupi_n_10614, csa_tree_add_51_79_groupi_n_10615, csa_tree_add_51_79_groupi_n_10616, csa_tree_add_51_79_groupi_n_10617, csa_tree_add_51_79_groupi_n_10618;
  wire csa_tree_add_51_79_groupi_n_10619, csa_tree_add_51_79_groupi_n_10620, csa_tree_add_51_79_groupi_n_10621, csa_tree_add_51_79_groupi_n_10622, csa_tree_add_51_79_groupi_n_10623, csa_tree_add_51_79_groupi_n_10624, csa_tree_add_51_79_groupi_n_10625, csa_tree_add_51_79_groupi_n_10626;
  wire csa_tree_add_51_79_groupi_n_10627, csa_tree_add_51_79_groupi_n_10628, csa_tree_add_51_79_groupi_n_10629, csa_tree_add_51_79_groupi_n_10630, csa_tree_add_51_79_groupi_n_10631, csa_tree_add_51_79_groupi_n_10632, csa_tree_add_51_79_groupi_n_10633, csa_tree_add_51_79_groupi_n_10634;
  wire csa_tree_add_51_79_groupi_n_10635, csa_tree_add_51_79_groupi_n_10636, csa_tree_add_51_79_groupi_n_10637, csa_tree_add_51_79_groupi_n_10638, csa_tree_add_51_79_groupi_n_10639, csa_tree_add_51_79_groupi_n_10640, csa_tree_add_51_79_groupi_n_10641, csa_tree_add_51_79_groupi_n_10642;
  wire csa_tree_add_51_79_groupi_n_10643, csa_tree_add_51_79_groupi_n_10644, csa_tree_add_51_79_groupi_n_10645, csa_tree_add_51_79_groupi_n_10646, csa_tree_add_51_79_groupi_n_10647, csa_tree_add_51_79_groupi_n_10648, csa_tree_add_51_79_groupi_n_10649, csa_tree_add_51_79_groupi_n_10650;
  wire csa_tree_add_51_79_groupi_n_10651, csa_tree_add_51_79_groupi_n_10652, csa_tree_add_51_79_groupi_n_10653, csa_tree_add_51_79_groupi_n_10654, csa_tree_add_51_79_groupi_n_10655, csa_tree_add_51_79_groupi_n_10656, csa_tree_add_51_79_groupi_n_10657, csa_tree_add_51_79_groupi_n_10658;
  wire csa_tree_add_51_79_groupi_n_10659, csa_tree_add_51_79_groupi_n_10660, csa_tree_add_51_79_groupi_n_10661, csa_tree_add_51_79_groupi_n_10662, csa_tree_add_51_79_groupi_n_10663, csa_tree_add_51_79_groupi_n_10664, csa_tree_add_51_79_groupi_n_10665, csa_tree_add_51_79_groupi_n_10666;
  wire csa_tree_add_51_79_groupi_n_10667, csa_tree_add_51_79_groupi_n_10668, csa_tree_add_51_79_groupi_n_10669, csa_tree_add_51_79_groupi_n_10670, csa_tree_add_51_79_groupi_n_10671, csa_tree_add_51_79_groupi_n_10672, csa_tree_add_51_79_groupi_n_10673, csa_tree_add_51_79_groupi_n_10674;
  wire csa_tree_add_51_79_groupi_n_10675, csa_tree_add_51_79_groupi_n_10676, csa_tree_add_51_79_groupi_n_10677, csa_tree_add_51_79_groupi_n_10678, csa_tree_add_51_79_groupi_n_10679, csa_tree_add_51_79_groupi_n_10680, csa_tree_add_51_79_groupi_n_10681, csa_tree_add_51_79_groupi_n_10682;
  wire csa_tree_add_51_79_groupi_n_10683, csa_tree_add_51_79_groupi_n_10684, csa_tree_add_51_79_groupi_n_10685, csa_tree_add_51_79_groupi_n_10686, csa_tree_add_51_79_groupi_n_10687, csa_tree_add_51_79_groupi_n_10688, csa_tree_add_51_79_groupi_n_10689, csa_tree_add_51_79_groupi_n_10690;
  wire csa_tree_add_51_79_groupi_n_10691, csa_tree_add_51_79_groupi_n_10692, csa_tree_add_51_79_groupi_n_10693, csa_tree_add_51_79_groupi_n_10694, csa_tree_add_51_79_groupi_n_10695, csa_tree_add_51_79_groupi_n_10696, csa_tree_add_51_79_groupi_n_10697, csa_tree_add_51_79_groupi_n_10698;
  wire csa_tree_add_51_79_groupi_n_10699, csa_tree_add_51_79_groupi_n_10700, csa_tree_add_51_79_groupi_n_10701, csa_tree_add_51_79_groupi_n_10702, csa_tree_add_51_79_groupi_n_10703, csa_tree_add_51_79_groupi_n_10704, csa_tree_add_51_79_groupi_n_10705, csa_tree_add_51_79_groupi_n_10706;
  wire csa_tree_add_51_79_groupi_n_10707, csa_tree_add_51_79_groupi_n_10708, csa_tree_add_51_79_groupi_n_10709, csa_tree_add_51_79_groupi_n_10711, csa_tree_add_51_79_groupi_n_10712, csa_tree_add_51_79_groupi_n_10713, csa_tree_add_51_79_groupi_n_10714, csa_tree_add_51_79_groupi_n_10715;
  wire csa_tree_add_51_79_groupi_n_10716, csa_tree_add_51_79_groupi_n_10717, csa_tree_add_51_79_groupi_n_10718, csa_tree_add_51_79_groupi_n_10719, csa_tree_add_51_79_groupi_n_10720, csa_tree_add_51_79_groupi_n_10721, csa_tree_add_51_79_groupi_n_10722, csa_tree_add_51_79_groupi_n_10723;
  wire csa_tree_add_51_79_groupi_n_10724, csa_tree_add_51_79_groupi_n_10725, csa_tree_add_51_79_groupi_n_10726, csa_tree_add_51_79_groupi_n_10727, csa_tree_add_51_79_groupi_n_10728, csa_tree_add_51_79_groupi_n_10729, csa_tree_add_51_79_groupi_n_10730, csa_tree_add_51_79_groupi_n_10731;
  wire csa_tree_add_51_79_groupi_n_10732, csa_tree_add_51_79_groupi_n_10733, csa_tree_add_51_79_groupi_n_10734, csa_tree_add_51_79_groupi_n_10735, csa_tree_add_51_79_groupi_n_10736, csa_tree_add_51_79_groupi_n_10737, csa_tree_add_51_79_groupi_n_10738, csa_tree_add_51_79_groupi_n_10739;
  wire csa_tree_add_51_79_groupi_n_10740, csa_tree_add_51_79_groupi_n_10741, csa_tree_add_51_79_groupi_n_10742, csa_tree_add_51_79_groupi_n_10743, csa_tree_add_51_79_groupi_n_10744, csa_tree_add_51_79_groupi_n_10745, csa_tree_add_51_79_groupi_n_10746, csa_tree_add_51_79_groupi_n_10747;
  wire csa_tree_add_51_79_groupi_n_10748, csa_tree_add_51_79_groupi_n_10749, csa_tree_add_51_79_groupi_n_10750, csa_tree_add_51_79_groupi_n_10751, csa_tree_add_51_79_groupi_n_10752, csa_tree_add_51_79_groupi_n_10753, csa_tree_add_51_79_groupi_n_10754, csa_tree_add_51_79_groupi_n_10755;
  wire csa_tree_add_51_79_groupi_n_10756, csa_tree_add_51_79_groupi_n_10757, csa_tree_add_51_79_groupi_n_10758, csa_tree_add_51_79_groupi_n_10759, csa_tree_add_51_79_groupi_n_10760, csa_tree_add_51_79_groupi_n_10761, csa_tree_add_51_79_groupi_n_10762, csa_tree_add_51_79_groupi_n_10763;
  wire csa_tree_add_51_79_groupi_n_10764, csa_tree_add_51_79_groupi_n_10765, csa_tree_add_51_79_groupi_n_10766, csa_tree_add_51_79_groupi_n_10767, csa_tree_add_51_79_groupi_n_10768, csa_tree_add_51_79_groupi_n_10769, csa_tree_add_51_79_groupi_n_10770, csa_tree_add_51_79_groupi_n_10771;
  wire csa_tree_add_51_79_groupi_n_10772, csa_tree_add_51_79_groupi_n_10773, csa_tree_add_51_79_groupi_n_10774, csa_tree_add_51_79_groupi_n_10775, csa_tree_add_51_79_groupi_n_10776, csa_tree_add_51_79_groupi_n_10777, csa_tree_add_51_79_groupi_n_10778, csa_tree_add_51_79_groupi_n_10779;
  wire csa_tree_add_51_79_groupi_n_10780, csa_tree_add_51_79_groupi_n_10781, csa_tree_add_51_79_groupi_n_10782, csa_tree_add_51_79_groupi_n_10783, csa_tree_add_51_79_groupi_n_10784, csa_tree_add_51_79_groupi_n_10785, csa_tree_add_51_79_groupi_n_10786, csa_tree_add_51_79_groupi_n_10787;
  wire csa_tree_add_51_79_groupi_n_10788, csa_tree_add_51_79_groupi_n_10789, csa_tree_add_51_79_groupi_n_10790, csa_tree_add_51_79_groupi_n_10791, csa_tree_add_51_79_groupi_n_10792, csa_tree_add_51_79_groupi_n_10793, csa_tree_add_51_79_groupi_n_10794, csa_tree_add_51_79_groupi_n_10795;
  wire csa_tree_add_51_79_groupi_n_10796, csa_tree_add_51_79_groupi_n_10797, csa_tree_add_51_79_groupi_n_10798, csa_tree_add_51_79_groupi_n_10799, csa_tree_add_51_79_groupi_n_10800, csa_tree_add_51_79_groupi_n_10801, csa_tree_add_51_79_groupi_n_10802, csa_tree_add_51_79_groupi_n_10803;
  wire csa_tree_add_51_79_groupi_n_10804, csa_tree_add_51_79_groupi_n_10805, csa_tree_add_51_79_groupi_n_10806, csa_tree_add_51_79_groupi_n_10807, csa_tree_add_51_79_groupi_n_10808, csa_tree_add_51_79_groupi_n_10809, csa_tree_add_51_79_groupi_n_10810, csa_tree_add_51_79_groupi_n_10811;
  wire csa_tree_add_51_79_groupi_n_10812, csa_tree_add_51_79_groupi_n_10813, csa_tree_add_51_79_groupi_n_10814, csa_tree_add_51_79_groupi_n_10815, csa_tree_add_51_79_groupi_n_10816, csa_tree_add_51_79_groupi_n_10817, csa_tree_add_51_79_groupi_n_10818, csa_tree_add_51_79_groupi_n_10819;
  wire csa_tree_add_51_79_groupi_n_10820, csa_tree_add_51_79_groupi_n_10821, csa_tree_add_51_79_groupi_n_10822, csa_tree_add_51_79_groupi_n_10823, csa_tree_add_51_79_groupi_n_10824, csa_tree_add_51_79_groupi_n_10825, csa_tree_add_51_79_groupi_n_10826, csa_tree_add_51_79_groupi_n_10827;
  wire csa_tree_add_51_79_groupi_n_10828, csa_tree_add_51_79_groupi_n_10829, csa_tree_add_51_79_groupi_n_10830, csa_tree_add_51_79_groupi_n_10831, csa_tree_add_51_79_groupi_n_10832, csa_tree_add_51_79_groupi_n_10833, csa_tree_add_51_79_groupi_n_10834, csa_tree_add_51_79_groupi_n_10835;
  wire csa_tree_add_51_79_groupi_n_10836, csa_tree_add_51_79_groupi_n_10837, csa_tree_add_51_79_groupi_n_10838, csa_tree_add_51_79_groupi_n_10839, csa_tree_add_51_79_groupi_n_10840, csa_tree_add_51_79_groupi_n_10841, csa_tree_add_51_79_groupi_n_10842, csa_tree_add_51_79_groupi_n_10843;
  wire csa_tree_add_51_79_groupi_n_10844, csa_tree_add_51_79_groupi_n_10845, csa_tree_add_51_79_groupi_n_10846, csa_tree_add_51_79_groupi_n_10847, csa_tree_add_51_79_groupi_n_10848, csa_tree_add_51_79_groupi_n_10849, csa_tree_add_51_79_groupi_n_10850, csa_tree_add_51_79_groupi_n_10851;
  wire csa_tree_add_51_79_groupi_n_10852, csa_tree_add_51_79_groupi_n_10853, csa_tree_add_51_79_groupi_n_10854, csa_tree_add_51_79_groupi_n_10855, csa_tree_add_51_79_groupi_n_10856, csa_tree_add_51_79_groupi_n_10857, csa_tree_add_51_79_groupi_n_10858, csa_tree_add_51_79_groupi_n_10859;
  wire csa_tree_add_51_79_groupi_n_10860, csa_tree_add_51_79_groupi_n_10861, csa_tree_add_51_79_groupi_n_10862, csa_tree_add_51_79_groupi_n_10863, csa_tree_add_51_79_groupi_n_10864, csa_tree_add_51_79_groupi_n_10865, csa_tree_add_51_79_groupi_n_10866, csa_tree_add_51_79_groupi_n_10867;
  wire csa_tree_add_51_79_groupi_n_10868, csa_tree_add_51_79_groupi_n_10869, csa_tree_add_51_79_groupi_n_10870, csa_tree_add_51_79_groupi_n_10871, csa_tree_add_51_79_groupi_n_10872, csa_tree_add_51_79_groupi_n_10873, csa_tree_add_51_79_groupi_n_10874, csa_tree_add_51_79_groupi_n_10875;
  wire csa_tree_add_51_79_groupi_n_10876, csa_tree_add_51_79_groupi_n_10877, csa_tree_add_51_79_groupi_n_10878, csa_tree_add_51_79_groupi_n_10879, csa_tree_add_51_79_groupi_n_10880, csa_tree_add_51_79_groupi_n_10881, csa_tree_add_51_79_groupi_n_10882, csa_tree_add_51_79_groupi_n_10883;
  wire csa_tree_add_51_79_groupi_n_10884, csa_tree_add_51_79_groupi_n_10885, csa_tree_add_51_79_groupi_n_10886, csa_tree_add_51_79_groupi_n_10887, csa_tree_add_51_79_groupi_n_10888, csa_tree_add_51_79_groupi_n_10889, csa_tree_add_51_79_groupi_n_10890, csa_tree_add_51_79_groupi_n_10891;
  wire csa_tree_add_51_79_groupi_n_10892, csa_tree_add_51_79_groupi_n_10893, csa_tree_add_51_79_groupi_n_10895, csa_tree_add_51_79_groupi_n_10896, csa_tree_add_51_79_groupi_n_10897, csa_tree_add_51_79_groupi_n_10898, csa_tree_add_51_79_groupi_n_10899, csa_tree_add_51_79_groupi_n_10900;
  wire csa_tree_add_51_79_groupi_n_10901, csa_tree_add_51_79_groupi_n_10902, csa_tree_add_51_79_groupi_n_10903, csa_tree_add_51_79_groupi_n_10904, csa_tree_add_51_79_groupi_n_10905, csa_tree_add_51_79_groupi_n_10906, csa_tree_add_51_79_groupi_n_10907, csa_tree_add_51_79_groupi_n_10908;
  wire csa_tree_add_51_79_groupi_n_10909, csa_tree_add_51_79_groupi_n_10910, csa_tree_add_51_79_groupi_n_10911, csa_tree_add_51_79_groupi_n_10912, csa_tree_add_51_79_groupi_n_10913, csa_tree_add_51_79_groupi_n_10914, csa_tree_add_51_79_groupi_n_10915, csa_tree_add_51_79_groupi_n_10916;
  wire csa_tree_add_51_79_groupi_n_10917, csa_tree_add_51_79_groupi_n_10918, csa_tree_add_51_79_groupi_n_10919, csa_tree_add_51_79_groupi_n_10920, csa_tree_add_51_79_groupi_n_10921, csa_tree_add_51_79_groupi_n_10922, csa_tree_add_51_79_groupi_n_10923, csa_tree_add_51_79_groupi_n_10924;
  wire csa_tree_add_51_79_groupi_n_10925, csa_tree_add_51_79_groupi_n_10926, csa_tree_add_51_79_groupi_n_10927, csa_tree_add_51_79_groupi_n_10928, csa_tree_add_51_79_groupi_n_10929, csa_tree_add_51_79_groupi_n_10930, csa_tree_add_51_79_groupi_n_10931, csa_tree_add_51_79_groupi_n_10932;
  wire csa_tree_add_51_79_groupi_n_10933, csa_tree_add_51_79_groupi_n_10934, csa_tree_add_51_79_groupi_n_10935, csa_tree_add_51_79_groupi_n_10936, csa_tree_add_51_79_groupi_n_10937, csa_tree_add_51_79_groupi_n_10938, csa_tree_add_51_79_groupi_n_10939, csa_tree_add_51_79_groupi_n_10940;
  wire csa_tree_add_51_79_groupi_n_10941, csa_tree_add_51_79_groupi_n_10942, csa_tree_add_51_79_groupi_n_10943, csa_tree_add_51_79_groupi_n_10944, csa_tree_add_51_79_groupi_n_10945, csa_tree_add_51_79_groupi_n_10946, csa_tree_add_51_79_groupi_n_10947, csa_tree_add_51_79_groupi_n_10948;
  wire csa_tree_add_51_79_groupi_n_10949, csa_tree_add_51_79_groupi_n_10950, csa_tree_add_51_79_groupi_n_10951, csa_tree_add_51_79_groupi_n_10952, csa_tree_add_51_79_groupi_n_10953, csa_tree_add_51_79_groupi_n_10954, csa_tree_add_51_79_groupi_n_10955, csa_tree_add_51_79_groupi_n_10956;
  wire csa_tree_add_51_79_groupi_n_10957, csa_tree_add_51_79_groupi_n_10958, csa_tree_add_51_79_groupi_n_10959, csa_tree_add_51_79_groupi_n_10960, csa_tree_add_51_79_groupi_n_10961, csa_tree_add_51_79_groupi_n_10962, csa_tree_add_51_79_groupi_n_10963, csa_tree_add_51_79_groupi_n_10964;
  wire csa_tree_add_51_79_groupi_n_10965, csa_tree_add_51_79_groupi_n_10966, csa_tree_add_51_79_groupi_n_10967, csa_tree_add_51_79_groupi_n_10968, csa_tree_add_51_79_groupi_n_10969, csa_tree_add_51_79_groupi_n_10970, csa_tree_add_51_79_groupi_n_10971, csa_tree_add_51_79_groupi_n_10972;
  wire csa_tree_add_51_79_groupi_n_10973, csa_tree_add_51_79_groupi_n_10974, csa_tree_add_51_79_groupi_n_10975, csa_tree_add_51_79_groupi_n_10976, csa_tree_add_51_79_groupi_n_10977, csa_tree_add_51_79_groupi_n_10978, csa_tree_add_51_79_groupi_n_10979, csa_tree_add_51_79_groupi_n_10980;
  wire csa_tree_add_51_79_groupi_n_10981, csa_tree_add_51_79_groupi_n_10982, csa_tree_add_51_79_groupi_n_10983, csa_tree_add_51_79_groupi_n_10984, csa_tree_add_51_79_groupi_n_10985, csa_tree_add_51_79_groupi_n_10986, csa_tree_add_51_79_groupi_n_10987, csa_tree_add_51_79_groupi_n_10988;
  wire csa_tree_add_51_79_groupi_n_10989, csa_tree_add_51_79_groupi_n_10990, csa_tree_add_51_79_groupi_n_10991, csa_tree_add_51_79_groupi_n_10992, csa_tree_add_51_79_groupi_n_10993, csa_tree_add_51_79_groupi_n_10994, csa_tree_add_51_79_groupi_n_10995, csa_tree_add_51_79_groupi_n_10996;
  wire csa_tree_add_51_79_groupi_n_10997, csa_tree_add_51_79_groupi_n_10998, csa_tree_add_51_79_groupi_n_10999, csa_tree_add_51_79_groupi_n_11000, csa_tree_add_51_79_groupi_n_11001, csa_tree_add_51_79_groupi_n_11002, csa_tree_add_51_79_groupi_n_11003, csa_tree_add_51_79_groupi_n_11004;
  wire csa_tree_add_51_79_groupi_n_11005, csa_tree_add_51_79_groupi_n_11006, csa_tree_add_51_79_groupi_n_11007, csa_tree_add_51_79_groupi_n_11008, csa_tree_add_51_79_groupi_n_11009, csa_tree_add_51_79_groupi_n_11010, csa_tree_add_51_79_groupi_n_11011, csa_tree_add_51_79_groupi_n_11012;
  wire csa_tree_add_51_79_groupi_n_11013, csa_tree_add_51_79_groupi_n_11014, csa_tree_add_51_79_groupi_n_11015, csa_tree_add_51_79_groupi_n_11016, csa_tree_add_51_79_groupi_n_11017, csa_tree_add_51_79_groupi_n_11018, csa_tree_add_51_79_groupi_n_11019, csa_tree_add_51_79_groupi_n_11020;
  wire csa_tree_add_51_79_groupi_n_11021, csa_tree_add_51_79_groupi_n_11022, csa_tree_add_51_79_groupi_n_11023, csa_tree_add_51_79_groupi_n_11024, csa_tree_add_51_79_groupi_n_11025, csa_tree_add_51_79_groupi_n_11026, csa_tree_add_51_79_groupi_n_11027, csa_tree_add_51_79_groupi_n_11028;
  wire csa_tree_add_51_79_groupi_n_11029, csa_tree_add_51_79_groupi_n_11030, csa_tree_add_51_79_groupi_n_11031, csa_tree_add_51_79_groupi_n_11032, csa_tree_add_51_79_groupi_n_11034, csa_tree_add_51_79_groupi_n_11035, csa_tree_add_51_79_groupi_n_11036, csa_tree_add_51_79_groupi_n_11037;
  wire csa_tree_add_51_79_groupi_n_11038, csa_tree_add_51_79_groupi_n_11039, csa_tree_add_51_79_groupi_n_11040, csa_tree_add_51_79_groupi_n_11041, csa_tree_add_51_79_groupi_n_11042, csa_tree_add_51_79_groupi_n_11043, csa_tree_add_51_79_groupi_n_11044, csa_tree_add_51_79_groupi_n_11045;
  wire csa_tree_add_51_79_groupi_n_11046, csa_tree_add_51_79_groupi_n_11047, csa_tree_add_51_79_groupi_n_11048, csa_tree_add_51_79_groupi_n_11049, csa_tree_add_51_79_groupi_n_11050, csa_tree_add_51_79_groupi_n_11051, csa_tree_add_51_79_groupi_n_11052, csa_tree_add_51_79_groupi_n_11053;
  wire csa_tree_add_51_79_groupi_n_11054, csa_tree_add_51_79_groupi_n_11055, csa_tree_add_51_79_groupi_n_11056, csa_tree_add_51_79_groupi_n_11057, csa_tree_add_51_79_groupi_n_11058, csa_tree_add_51_79_groupi_n_11059, csa_tree_add_51_79_groupi_n_11060, csa_tree_add_51_79_groupi_n_11061;
  wire csa_tree_add_51_79_groupi_n_11063, csa_tree_add_51_79_groupi_n_11064, csa_tree_add_51_79_groupi_n_11065, csa_tree_add_51_79_groupi_n_11066, csa_tree_add_51_79_groupi_n_11067, csa_tree_add_51_79_groupi_n_11068, csa_tree_add_51_79_groupi_n_11069, csa_tree_add_51_79_groupi_n_11070;
  wire csa_tree_add_51_79_groupi_n_11071, csa_tree_add_51_79_groupi_n_11072, csa_tree_add_51_79_groupi_n_11073, csa_tree_add_51_79_groupi_n_11074, csa_tree_add_51_79_groupi_n_11075, csa_tree_add_51_79_groupi_n_11076, csa_tree_add_51_79_groupi_n_11077, csa_tree_add_51_79_groupi_n_11078;
  wire csa_tree_add_51_79_groupi_n_11079, csa_tree_add_51_79_groupi_n_11080, csa_tree_add_51_79_groupi_n_11081, csa_tree_add_51_79_groupi_n_11082, csa_tree_add_51_79_groupi_n_11083, csa_tree_add_51_79_groupi_n_11084, csa_tree_add_51_79_groupi_n_11085, csa_tree_add_51_79_groupi_n_11086;
  wire csa_tree_add_51_79_groupi_n_11087, csa_tree_add_51_79_groupi_n_11088, csa_tree_add_51_79_groupi_n_11089, csa_tree_add_51_79_groupi_n_11090, csa_tree_add_51_79_groupi_n_11091, csa_tree_add_51_79_groupi_n_11092, csa_tree_add_51_79_groupi_n_11093, csa_tree_add_51_79_groupi_n_11094;
  wire csa_tree_add_51_79_groupi_n_11095, csa_tree_add_51_79_groupi_n_11096, csa_tree_add_51_79_groupi_n_11097, csa_tree_add_51_79_groupi_n_11098, csa_tree_add_51_79_groupi_n_11099, csa_tree_add_51_79_groupi_n_11100, csa_tree_add_51_79_groupi_n_11101, csa_tree_add_51_79_groupi_n_11102;
  wire csa_tree_add_51_79_groupi_n_11103, csa_tree_add_51_79_groupi_n_11104, csa_tree_add_51_79_groupi_n_11105, csa_tree_add_51_79_groupi_n_11106, csa_tree_add_51_79_groupi_n_11107, csa_tree_add_51_79_groupi_n_11108, csa_tree_add_51_79_groupi_n_11109, csa_tree_add_51_79_groupi_n_11110;
  wire csa_tree_add_51_79_groupi_n_11111, csa_tree_add_51_79_groupi_n_11112, csa_tree_add_51_79_groupi_n_11113, csa_tree_add_51_79_groupi_n_11114, csa_tree_add_51_79_groupi_n_11115, csa_tree_add_51_79_groupi_n_11116, csa_tree_add_51_79_groupi_n_11117, csa_tree_add_51_79_groupi_n_11119;
  wire csa_tree_add_51_79_groupi_n_11120, csa_tree_add_51_79_groupi_n_11121, csa_tree_add_51_79_groupi_n_11122, csa_tree_add_51_79_groupi_n_11123, csa_tree_add_51_79_groupi_n_11124, csa_tree_add_51_79_groupi_n_11125, csa_tree_add_51_79_groupi_n_11126, csa_tree_add_51_79_groupi_n_11127;
  wire csa_tree_add_51_79_groupi_n_11128, csa_tree_add_51_79_groupi_n_11129, csa_tree_add_51_79_groupi_n_11130, csa_tree_add_51_79_groupi_n_11131, csa_tree_add_51_79_groupi_n_11132, csa_tree_add_51_79_groupi_n_11133, csa_tree_add_51_79_groupi_n_11134, csa_tree_add_51_79_groupi_n_11135;
  wire csa_tree_add_51_79_groupi_n_11136, csa_tree_add_51_79_groupi_n_11137, csa_tree_add_51_79_groupi_n_11138, csa_tree_add_51_79_groupi_n_11139, csa_tree_add_51_79_groupi_n_11140, csa_tree_add_51_79_groupi_n_11141, csa_tree_add_51_79_groupi_n_11142, csa_tree_add_51_79_groupi_n_11143;
  wire csa_tree_add_51_79_groupi_n_11144, csa_tree_add_51_79_groupi_n_11145, csa_tree_add_51_79_groupi_n_11146, csa_tree_add_51_79_groupi_n_11147, csa_tree_add_51_79_groupi_n_11148, csa_tree_add_51_79_groupi_n_11149, csa_tree_add_51_79_groupi_n_11150, csa_tree_add_51_79_groupi_n_11151;
  wire csa_tree_add_51_79_groupi_n_11152, csa_tree_add_51_79_groupi_n_11153, csa_tree_add_51_79_groupi_n_11154, csa_tree_add_51_79_groupi_n_11155, csa_tree_add_51_79_groupi_n_11156, csa_tree_add_51_79_groupi_n_11158, csa_tree_add_51_79_groupi_n_11159, csa_tree_add_51_79_groupi_n_11160;
  wire csa_tree_add_51_79_groupi_n_11161, csa_tree_add_51_79_groupi_n_11162, csa_tree_add_51_79_groupi_n_11163, csa_tree_add_51_79_groupi_n_11164, csa_tree_add_51_79_groupi_n_11165, csa_tree_add_51_79_groupi_n_11166, csa_tree_add_51_79_groupi_n_11167, csa_tree_add_51_79_groupi_n_11168;
  wire csa_tree_add_51_79_groupi_n_11169, csa_tree_add_51_79_groupi_n_11170, csa_tree_add_51_79_groupi_n_11171, csa_tree_add_51_79_groupi_n_11172, csa_tree_add_51_79_groupi_n_11173, csa_tree_add_51_79_groupi_n_11174, csa_tree_add_51_79_groupi_n_11175, csa_tree_add_51_79_groupi_n_11176;
  wire csa_tree_add_51_79_groupi_n_11178, csa_tree_add_51_79_groupi_n_11179, csa_tree_add_51_79_groupi_n_11180, csa_tree_add_51_79_groupi_n_11181, csa_tree_add_51_79_groupi_n_11183, csa_tree_add_51_79_groupi_n_11184, csa_tree_add_51_79_groupi_n_11186, csa_tree_add_51_79_groupi_n_11187;
  wire csa_tree_add_51_79_groupi_n_11189, csa_tree_add_51_79_groupi_n_11190, csa_tree_add_51_79_groupi_n_11192, csa_tree_add_51_79_groupi_n_11193, csa_tree_add_51_79_groupi_n_11195, csa_tree_add_51_79_groupi_n_11196, csa_tree_add_51_79_groupi_n_11198, csa_tree_add_51_79_groupi_n_11199;
  wire csa_tree_add_51_79_groupi_n_11201, csa_tree_add_51_79_groupi_n_11202, csa_tree_add_51_79_groupi_n_11204, csa_tree_add_51_79_groupi_n_11205, csa_tree_add_51_79_groupi_n_11207, csa_tree_add_51_79_groupi_n_11208, csa_tree_add_51_79_groupi_n_11210, csa_tree_add_51_79_groupi_n_11211;
  wire csa_tree_add_51_79_groupi_n_11213, csa_tree_add_51_79_groupi_n_11214, csa_tree_add_51_79_groupi_n_11216, csa_tree_add_51_79_groupi_n_11217, csa_tree_add_51_79_groupi_n_11219, csa_tree_add_51_79_groupi_n_11220, csa_tree_add_51_79_groupi_n_11222, csa_tree_add_51_79_groupi_n_11223;
  wire csa_tree_add_51_79_groupi_n_11225;
  xnor csa_tree_add_51_79_groupi_g34832__2398(out1[25] ,csa_tree_add_51_79_groupi_n_11225 ,csa_tree_add_51_79_groupi_n_10164);
  nor csa_tree_add_51_79_groupi_g34833__5107(csa_tree_add_51_79_groupi_n_11225 ,csa_tree_add_51_79_groupi_n_10778 ,csa_tree_add_51_79_groupi_n_11223);
  xnor csa_tree_add_51_79_groupi_g34834__6260(out1[24] ,csa_tree_add_51_79_groupi_n_11222 ,csa_tree_add_51_79_groupi_n_10837);
  nor csa_tree_add_51_79_groupi_g34835__4319(csa_tree_add_51_79_groupi_n_11223 ,csa_tree_add_51_79_groupi_n_10813 ,csa_tree_add_51_79_groupi_n_11222);
  and csa_tree_add_51_79_groupi_g34836__8428(csa_tree_add_51_79_groupi_n_11222 ,csa_tree_add_51_79_groupi_n_10970 ,csa_tree_add_51_79_groupi_n_11220);
  xnor csa_tree_add_51_79_groupi_g34837__5526(out1[23] ,csa_tree_add_51_79_groupi_n_11219 ,csa_tree_add_51_79_groupi_n_38);
  or csa_tree_add_51_79_groupi_g34838__6783(csa_tree_add_51_79_groupi_n_11220 ,csa_tree_add_51_79_groupi_n_11219 ,csa_tree_add_51_79_groupi_n_10949);
  and csa_tree_add_51_79_groupi_g34839__3680(csa_tree_add_51_79_groupi_n_11219 ,csa_tree_add_51_79_groupi_n_10998 ,csa_tree_add_51_79_groupi_n_11217);
  xnor csa_tree_add_51_79_groupi_g34840__1617(out1[22] ,csa_tree_add_51_79_groupi_n_11216 ,csa_tree_add_51_79_groupi_n_11031);
  or csa_tree_add_51_79_groupi_g34841__2802(csa_tree_add_51_79_groupi_n_11217 ,csa_tree_add_51_79_groupi_n_11010 ,csa_tree_add_51_79_groupi_n_11216);
  and csa_tree_add_51_79_groupi_g34842__1705(csa_tree_add_51_79_groupi_n_11216 ,csa_tree_add_51_79_groupi_n_11078 ,csa_tree_add_51_79_groupi_n_11214);
  xnor csa_tree_add_51_79_groupi_g34843__5122(out1[21] ,csa_tree_add_51_79_groupi_n_11213 ,csa_tree_add_51_79_groupi_n_11088);
  or csa_tree_add_51_79_groupi_g34844__8246(csa_tree_add_51_79_groupi_n_11214 ,csa_tree_add_51_79_groupi_n_11073 ,csa_tree_add_51_79_groupi_n_11213);
  and csa_tree_add_51_79_groupi_g34845__7098(csa_tree_add_51_79_groupi_n_11213 ,csa_tree_add_51_79_groupi_n_11107 ,csa_tree_add_51_79_groupi_n_11211);
  xnor csa_tree_add_51_79_groupi_g34846__6131(out1[20] ,csa_tree_add_51_79_groupi_n_11210 ,csa_tree_add_51_79_groupi_n_11115);
  or csa_tree_add_51_79_groupi_g34847__1881(csa_tree_add_51_79_groupi_n_11211 ,csa_tree_add_51_79_groupi_n_11210 ,csa_tree_add_51_79_groupi_n_11091);
  and csa_tree_add_51_79_groupi_g34848__5115(csa_tree_add_51_79_groupi_n_11210 ,csa_tree_add_51_79_groupi_n_11208 ,csa_tree_add_51_79_groupi_n_11117);
  xnor csa_tree_add_51_79_groupi_g34849__7482(out1[19] ,csa_tree_add_51_79_groupi_n_11207 ,csa_tree_add_51_79_groupi_n_11135);
  or csa_tree_add_51_79_groupi_g34850__4733(csa_tree_add_51_79_groupi_n_11208 ,csa_tree_add_51_79_groupi_n_11127 ,csa_tree_add_51_79_groupi_n_11207);
  and csa_tree_add_51_79_groupi_g34851__6161(csa_tree_add_51_79_groupi_n_11207 ,csa_tree_add_51_79_groupi_n_11136 ,csa_tree_add_51_79_groupi_n_11205);
  xnor csa_tree_add_51_79_groupi_g34852__9315(out1[18] ,csa_tree_add_51_79_groupi_n_11204 ,csa_tree_add_51_79_groupi_n_11155);
  or csa_tree_add_51_79_groupi_g34853__9945(csa_tree_add_51_79_groupi_n_11205 ,csa_tree_add_51_79_groupi_n_11145 ,csa_tree_add_51_79_groupi_n_11204);
  and csa_tree_add_51_79_groupi_g34854__2883(csa_tree_add_51_79_groupi_n_11204 ,csa_tree_add_51_79_groupi_n_11202 ,csa_tree_add_51_79_groupi_n_11158);
  xnor csa_tree_add_51_79_groupi_g34855__2346(out1[17] ,csa_tree_add_51_79_groupi_n_11201 ,csa_tree_add_51_79_groupi_n_11171);
  or csa_tree_add_51_79_groupi_g34856__1666(csa_tree_add_51_79_groupi_n_11202 ,csa_tree_add_51_79_groupi_n_11164 ,csa_tree_add_51_79_groupi_n_11201);
  and csa_tree_add_51_79_groupi_g34857__7410(csa_tree_add_51_79_groupi_n_11201 ,csa_tree_add_51_79_groupi_n_11175 ,csa_tree_add_51_79_groupi_n_11199);
  xnor csa_tree_add_51_79_groupi_g34858__6417(out1[16] ,csa_tree_add_51_79_groupi_n_11198 ,csa_tree_add_51_79_groupi_n_11179);
  or csa_tree_add_51_79_groupi_g34859__5477(csa_tree_add_51_79_groupi_n_11199 ,csa_tree_add_51_79_groupi_n_11174 ,csa_tree_add_51_79_groupi_n_11198);
  and csa_tree_add_51_79_groupi_g34860__2398(csa_tree_add_51_79_groupi_n_11198 ,csa_tree_add_51_79_groupi_n_11196 ,csa_tree_add_51_79_groupi_n_11172);
  xnor csa_tree_add_51_79_groupi_g34861__5107(out1[15] ,csa_tree_add_51_79_groupi_n_11195 ,csa_tree_add_51_79_groupi_n_11178);
  or csa_tree_add_51_79_groupi_g34862__6260(csa_tree_add_51_79_groupi_n_11196 ,csa_tree_add_51_79_groupi_n_11195 ,csa_tree_add_51_79_groupi_n_11173);
  and csa_tree_add_51_79_groupi_g34863__4319(csa_tree_add_51_79_groupi_n_11195 ,csa_tree_add_51_79_groupi_n_11167 ,csa_tree_add_51_79_groupi_n_11193);
  xnor csa_tree_add_51_79_groupi_g34864__8428(out1[14] ,csa_tree_add_51_79_groupi_n_11192 ,csa_tree_add_51_79_groupi_n_11170);
  or csa_tree_add_51_79_groupi_g34865__5526(csa_tree_add_51_79_groupi_n_11193 ,csa_tree_add_51_79_groupi_n_11192 ,csa_tree_add_51_79_groupi_n_11165);
  and csa_tree_add_51_79_groupi_g34866__6783(csa_tree_add_51_79_groupi_n_11192 ,csa_tree_add_51_79_groupi_n_11190 ,csa_tree_add_51_79_groupi_n_11163);
  xnor csa_tree_add_51_79_groupi_g34867__3680(out1[13] ,csa_tree_add_51_79_groupi_n_11189 ,csa_tree_add_51_79_groupi_n_11169);
  or csa_tree_add_51_79_groupi_g34868__1617(csa_tree_add_51_79_groupi_n_11190 ,csa_tree_add_51_79_groupi_n_11189 ,csa_tree_add_51_79_groupi_n_11166);
  and csa_tree_add_51_79_groupi_g34869__2802(csa_tree_add_51_79_groupi_n_11189 ,csa_tree_add_51_79_groupi_n_11187 ,csa_tree_add_51_79_groupi_n_11137);
  xnor csa_tree_add_51_79_groupi_g34870__1705(out1[12] ,csa_tree_add_51_79_groupi_n_11186 ,csa_tree_add_51_79_groupi_n_11156);
  or csa_tree_add_51_79_groupi_g34871__5122(csa_tree_add_51_79_groupi_n_11187 ,csa_tree_add_51_79_groupi_n_11147 ,csa_tree_add_51_79_groupi_n_11186);
  and csa_tree_add_51_79_groupi_g34872__8246(csa_tree_add_51_79_groupi_n_11186 ,csa_tree_add_51_79_groupi_n_11184 ,csa_tree_add_51_79_groupi_n_11125);
  xnor csa_tree_add_51_79_groupi_g34873__7098(out1[11] ,csa_tree_add_51_79_groupi_n_11183 ,csa_tree_add_51_79_groupi_n_11134);
  or csa_tree_add_51_79_groupi_g34874__6131(csa_tree_add_51_79_groupi_n_11184 ,csa_tree_add_51_79_groupi_n_11183 ,csa_tree_add_51_79_groupi_n_11132);
  and csa_tree_add_51_79_groupi_g34875__1881(csa_tree_add_51_79_groupi_n_11183 ,csa_tree_add_51_79_groupi_n_11181 ,csa_tree_add_51_79_groupi_n_11100);
  xnor csa_tree_add_51_79_groupi_g34876__5115(out1[10] ,csa_tree_add_51_79_groupi_n_11180 ,csa_tree_add_51_79_groupi_n_11116);
  or csa_tree_add_51_79_groupi_g34877__7482(csa_tree_add_51_79_groupi_n_11181 ,csa_tree_add_51_79_groupi_n_11099 ,csa_tree_add_51_79_groupi_n_11180);
  and csa_tree_add_51_79_groupi_g34878__4733(csa_tree_add_51_79_groupi_n_11180 ,csa_tree_add_51_79_groupi_n_11074 ,csa_tree_add_51_79_groupi_n_11176);
  xnor csa_tree_add_51_79_groupi_g34879__6161(csa_tree_add_51_79_groupi_n_11179 ,csa_tree_add_51_79_groupi_n_11152 ,csa_tree_add_51_79_groupi_n_11159);
  xnor csa_tree_add_51_79_groupi_g34880__9315(csa_tree_add_51_79_groupi_n_11178 ,csa_tree_add_51_79_groupi_n_11162 ,csa_tree_add_51_79_groupi_n_11149);
  xnor csa_tree_add_51_79_groupi_g34881__9945(out1[9] ,csa_tree_add_51_79_groupi_n_11168 ,csa_tree_add_51_79_groupi_n_11087);
  or csa_tree_add_51_79_groupi_g34882__2883(csa_tree_add_51_79_groupi_n_11176 ,csa_tree_add_51_79_groupi_n_11077 ,csa_tree_add_51_79_groupi_n_11168);
  or csa_tree_add_51_79_groupi_g34883__2346(csa_tree_add_51_79_groupi_n_11175 ,csa_tree_add_51_79_groupi_n_11152 ,csa_tree_add_51_79_groupi_n_11160);
  and csa_tree_add_51_79_groupi_g34884__1666(csa_tree_add_51_79_groupi_n_11174 ,csa_tree_add_51_79_groupi_n_11152 ,csa_tree_add_51_79_groupi_n_11160);
  nor csa_tree_add_51_79_groupi_g34885__7410(csa_tree_add_51_79_groupi_n_11173 ,csa_tree_add_51_79_groupi_n_11161 ,csa_tree_add_51_79_groupi_n_11149);
  or csa_tree_add_51_79_groupi_g34886__6417(csa_tree_add_51_79_groupi_n_11172 ,csa_tree_add_51_79_groupi_n_11162 ,csa_tree_add_51_79_groupi_n_11148);
  xnor csa_tree_add_51_79_groupi_g34887__5477(csa_tree_add_51_79_groupi_n_11171 ,csa_tree_add_51_79_groupi_n_11138 ,csa_tree_add_51_79_groupi_n_11151);
  xnor csa_tree_add_51_79_groupi_g34888__2398(csa_tree_add_51_79_groupi_n_11170 ,csa_tree_add_51_79_groupi_n_11140 ,csa_tree_add_51_79_groupi_n_11154);
  xnor csa_tree_add_51_79_groupi_g34889__5107(csa_tree_add_51_79_groupi_n_11169 ,csa_tree_add_51_79_groupi_n_11142 ,csa_tree_add_51_79_groupi_n_11144);
  or csa_tree_add_51_79_groupi_g34890__6260(csa_tree_add_51_79_groupi_n_11167 ,csa_tree_add_51_79_groupi_n_11139 ,csa_tree_add_51_79_groupi_n_11154);
  nor csa_tree_add_51_79_groupi_g34891__4319(csa_tree_add_51_79_groupi_n_11166 ,csa_tree_add_51_79_groupi_n_11141 ,csa_tree_add_51_79_groupi_n_11144);
  nor csa_tree_add_51_79_groupi_g34892__8428(csa_tree_add_51_79_groupi_n_11165 ,csa_tree_add_51_79_groupi_n_11140 ,csa_tree_add_51_79_groupi_n_11153);
  nor csa_tree_add_51_79_groupi_g34893__5526(csa_tree_add_51_79_groupi_n_11164 ,csa_tree_add_51_79_groupi_n_43 ,csa_tree_add_51_79_groupi_n_11151);
  or csa_tree_add_51_79_groupi_g34894__6783(csa_tree_add_51_79_groupi_n_11163 ,csa_tree_add_51_79_groupi_n_11142 ,csa_tree_add_51_79_groupi_n_11143);
  and csa_tree_add_51_79_groupi_g34895__3680(csa_tree_add_51_79_groupi_n_11168 ,csa_tree_add_51_79_groupi_n_11146 ,csa_tree_add_51_79_groupi_n_11034);
  not csa_tree_add_51_79_groupi_g34896(csa_tree_add_51_79_groupi_n_11162 ,csa_tree_add_51_79_groupi_n_11161);
  not csa_tree_add_51_79_groupi_g34897(csa_tree_add_51_79_groupi_n_11160 ,csa_tree_add_51_79_groupi_n_11159);
  or csa_tree_add_51_79_groupi_g34898__1617(csa_tree_add_51_79_groupi_n_11158 ,csa_tree_add_51_79_groupi_n_11138 ,csa_tree_add_51_79_groupi_n_11150);
  xnor csa_tree_add_51_79_groupi_g34899__2802(out1[8] ,csa_tree_add_51_79_groupi_n_11133 ,csa_tree_add_51_79_groupi_n_11059);
  xnor csa_tree_add_51_79_groupi_g34900__1705(csa_tree_add_51_79_groupi_n_11156 ,csa_tree_add_51_79_groupi_n_11120 ,csa_tree_add_51_79_groupi_n_11112);
  xnor csa_tree_add_51_79_groupi_g34901__5122(csa_tree_add_51_79_groupi_n_11155 ,csa_tree_add_51_79_groupi_n_11124 ,csa_tree_add_51_79_groupi_n_11122);
  xnor csa_tree_add_51_79_groupi_g34902__8246(csa_tree_add_51_79_groupi_n_11161 ,csa_tree_add_51_79_groupi_n_11070 ,csa_tree_add_51_79_groupi_n_11114);
  xnor csa_tree_add_51_79_groupi_g34903__7098(csa_tree_add_51_79_groupi_n_11159 ,csa_tree_add_51_79_groupi_n_11056 ,csa_tree_add_51_79_groupi_n_11113);
  not csa_tree_add_51_79_groupi_g34904(csa_tree_add_51_79_groupi_n_11153 ,csa_tree_add_51_79_groupi_n_11154);
  not csa_tree_add_51_79_groupi_g34905(csa_tree_add_51_79_groupi_n_11151 ,csa_tree_add_51_79_groupi_n_11150);
  not csa_tree_add_51_79_groupi_g34906(csa_tree_add_51_79_groupi_n_11149 ,csa_tree_add_51_79_groupi_n_11148);
  nor csa_tree_add_51_79_groupi_g34907__6131(csa_tree_add_51_79_groupi_n_11147 ,csa_tree_add_51_79_groupi_n_11119 ,csa_tree_add_51_79_groupi_n_11112);
  or csa_tree_add_51_79_groupi_g34908__1881(csa_tree_add_51_79_groupi_n_11146 ,csa_tree_add_51_79_groupi_n_11133 ,csa_tree_add_51_79_groupi_n_11046);
  nor csa_tree_add_51_79_groupi_g34909__5115(csa_tree_add_51_79_groupi_n_11145 ,csa_tree_add_51_79_groupi_n_11123 ,csa_tree_add_51_79_groupi_n_11122);
  and csa_tree_add_51_79_groupi_g34910__7482(csa_tree_add_51_79_groupi_n_11154 ,csa_tree_add_51_79_groupi_n_11131 ,csa_tree_add_51_79_groupi_n_11101);
  and csa_tree_add_51_79_groupi_g34911__4733(csa_tree_add_51_79_groupi_n_11152 ,csa_tree_add_51_79_groupi_n_11128 ,csa_tree_add_51_79_groupi_n_11103);
  and csa_tree_add_51_79_groupi_g34912__6161(csa_tree_add_51_79_groupi_n_11150 ,csa_tree_add_51_79_groupi_n_11106 ,csa_tree_add_51_79_groupi_n_11129);
  and csa_tree_add_51_79_groupi_g34913__9315(csa_tree_add_51_79_groupi_n_11148 ,csa_tree_add_51_79_groupi_n_11130 ,csa_tree_add_51_79_groupi_n_11075);
  not csa_tree_add_51_79_groupi_g34914(csa_tree_add_51_79_groupi_n_11144 ,csa_tree_add_51_79_groupi_n_11143);
  not csa_tree_add_51_79_groupi_g34915(csa_tree_add_51_79_groupi_n_11142 ,csa_tree_add_51_79_groupi_n_11141);
  not csa_tree_add_51_79_groupi_g34916(csa_tree_add_51_79_groupi_n_11140 ,csa_tree_add_51_79_groupi_n_11139);
  not csa_tree_add_51_79_groupi_g34917(csa_tree_add_51_79_groupi_n_11138 ,csa_tree_add_51_79_groupi_n_43);
  or csa_tree_add_51_79_groupi_g34918__9945(csa_tree_add_51_79_groupi_n_11137 ,csa_tree_add_51_79_groupi_n_11120 ,csa_tree_add_51_79_groupi_n_11111);
  or csa_tree_add_51_79_groupi_g34919__2883(csa_tree_add_51_79_groupi_n_11136 ,csa_tree_add_51_79_groupi_n_11124 ,csa_tree_add_51_79_groupi_n_11121);
  xnor csa_tree_add_51_79_groupi_g34920__2346(csa_tree_add_51_79_groupi_n_11135 ,csa_tree_add_51_79_groupi_n_11110 ,csa_tree_add_51_79_groupi_n_11097);
  xnor csa_tree_add_51_79_groupi_g34921__1666(csa_tree_add_51_79_groupi_n_11134 ,csa_tree_add_51_79_groupi_n_11080 ,csa_tree_add_51_79_groupi_n_11095);
  and csa_tree_add_51_79_groupi_g34922__7410(csa_tree_add_51_79_groupi_n_11143 ,csa_tree_add_51_79_groupi_n_11093 ,csa_tree_add_51_79_groupi_n_11126);
  xnor csa_tree_add_51_79_groupi_g34923__6417(csa_tree_add_51_79_groupi_n_11141 ,csa_tree_add_51_79_groupi_n_11065 ,csa_tree_add_51_79_groupi_n_11086);
  xnor csa_tree_add_51_79_groupi_g34924__5477(csa_tree_add_51_79_groupi_n_11139 ,csa_tree_add_51_79_groupi_n_11098 ,csa_tree_add_51_79_groupi_n_11089);
  nor csa_tree_add_51_79_groupi_g34926__2398(csa_tree_add_51_79_groupi_n_11132 ,csa_tree_add_51_79_groupi_n_11079 ,csa_tree_add_51_79_groupi_n_11095);
  or csa_tree_add_51_79_groupi_g34927__5107(csa_tree_add_51_79_groupi_n_11131 ,csa_tree_add_51_79_groupi_n_11054 ,csa_tree_add_51_79_groupi_n_11108);
  or csa_tree_add_51_79_groupi_g34928__6260(csa_tree_add_51_79_groupi_n_11130 ,csa_tree_add_51_79_groupi_n_11098 ,csa_tree_add_51_79_groupi_n_11076);
  or csa_tree_add_51_79_groupi_g34929__4319(csa_tree_add_51_79_groupi_n_11129 ,csa_tree_add_51_79_groupi_n_11056 ,csa_tree_add_51_79_groupi_n_11105);
  or csa_tree_add_51_79_groupi_g34930__8428(csa_tree_add_51_79_groupi_n_11128 ,csa_tree_add_51_79_groupi_n_11070 ,csa_tree_add_51_79_groupi_n_11104);
  nor csa_tree_add_51_79_groupi_g34931__5526(csa_tree_add_51_79_groupi_n_11127 ,csa_tree_add_51_79_groupi_n_11109 ,csa_tree_add_51_79_groupi_n_11097);
  or csa_tree_add_51_79_groupi_g34932__6783(csa_tree_add_51_79_groupi_n_11126 ,csa_tree_add_51_79_groupi_n_11090 ,csa_tree_add_51_79_groupi_n_11026);
  or csa_tree_add_51_79_groupi_g34933__3680(csa_tree_add_51_79_groupi_n_11125 ,csa_tree_add_51_79_groupi_n_11080 ,csa_tree_add_51_79_groupi_n_11094);
  and csa_tree_add_51_79_groupi_g34934__1617(csa_tree_add_51_79_groupi_n_11133 ,csa_tree_add_51_79_groupi_n_10996 ,csa_tree_add_51_79_groupi_n_11102);
  not csa_tree_add_51_79_groupi_g34935(csa_tree_add_51_79_groupi_n_11123 ,csa_tree_add_51_79_groupi_n_11124);
  not csa_tree_add_51_79_groupi_g34936(csa_tree_add_51_79_groupi_n_11122 ,csa_tree_add_51_79_groupi_n_11121);
  not csa_tree_add_51_79_groupi_g34937(csa_tree_add_51_79_groupi_n_11120 ,csa_tree_add_51_79_groupi_n_11119);
  xnor csa_tree_add_51_79_groupi_g34938__2802(out1[7] ,csa_tree_add_51_79_groupi_n_11084 ,csa_tree_add_51_79_groupi_n_11032);
  or csa_tree_add_51_79_groupi_g34939__1705(csa_tree_add_51_79_groupi_n_11117 ,csa_tree_add_51_79_groupi_n_11110 ,csa_tree_add_51_79_groupi_n_11096);
  xnor csa_tree_add_51_79_groupi_g34940__5122(csa_tree_add_51_79_groupi_n_11116 ,csa_tree_add_51_79_groupi_n_11053 ,csa_tree_add_51_79_groupi_n_11067);
  xnor csa_tree_add_51_79_groupi_g34941__8246(csa_tree_add_51_79_groupi_n_11115 ,csa_tree_add_51_79_groupi_n_11083 ,csa_tree_add_51_79_groupi_n_41);
  xnor csa_tree_add_51_79_groupi_g34942__7098(csa_tree_add_51_79_groupi_n_11114 ,csa_tree_add_51_79_groupi_n_10985 ,csa_tree_add_51_79_groupi_n_11082);
  xnor csa_tree_add_51_79_groupi_g34943__6131(csa_tree_add_51_79_groupi_n_11113 ,csa_tree_add_51_79_groupi_n_11007 ,csa_tree_add_51_79_groupi_n_11063);
  and csa_tree_add_51_79_groupi_g34944__1881(csa_tree_add_51_79_groupi_n_11124 ,csa_tree_add_51_79_groupi_n_11060 ,csa_tree_add_51_79_groupi_n_11092);
  xnor csa_tree_add_51_79_groupi_g34945__5115(csa_tree_add_51_79_groupi_n_11121 ,csa_tree_add_51_79_groupi_n_11055 ,csa_tree_add_51_79_groupi_n_11057);
  xnor csa_tree_add_51_79_groupi_g34946__7482(csa_tree_add_51_79_groupi_n_11119 ,csa_tree_add_51_79_groupi_n_11069 ,csa_tree_add_51_79_groupi_n_11058);
  not csa_tree_add_51_79_groupi_g34947(csa_tree_add_51_79_groupi_n_11111 ,csa_tree_add_51_79_groupi_n_11112);
  not csa_tree_add_51_79_groupi_g34948(csa_tree_add_51_79_groupi_n_11109 ,csa_tree_add_51_79_groupi_n_11110);
  nor csa_tree_add_51_79_groupi_g34949__4733(csa_tree_add_51_79_groupi_n_11108 ,csa_tree_add_51_79_groupi_n_11040 ,csa_tree_add_51_79_groupi_n_11065);
  or csa_tree_add_51_79_groupi_g34950__6161(csa_tree_add_51_79_groupi_n_11107 ,csa_tree_add_51_79_groupi_n_11083 ,csa_tree_add_51_79_groupi_n_11068);
  or csa_tree_add_51_79_groupi_g34951__9315(csa_tree_add_51_79_groupi_n_11106 ,csa_tree_add_51_79_groupi_n_11007 ,csa_tree_add_51_79_groupi_n_42);
  nor csa_tree_add_51_79_groupi_g34952__9945(csa_tree_add_51_79_groupi_n_11105 ,csa_tree_add_51_79_groupi_n_11006 ,csa_tree_add_51_79_groupi_n_11063);
  nor csa_tree_add_51_79_groupi_g34953__2883(csa_tree_add_51_79_groupi_n_11104 ,csa_tree_add_51_79_groupi_n_10984 ,csa_tree_add_51_79_groupi_n_11082);
  or csa_tree_add_51_79_groupi_g34954__2346(csa_tree_add_51_79_groupi_n_11103 ,csa_tree_add_51_79_groupi_n_10985 ,csa_tree_add_51_79_groupi_n_11081);
  or csa_tree_add_51_79_groupi_g34955__1666(csa_tree_add_51_79_groupi_n_11102 ,csa_tree_add_51_79_groupi_n_10997 ,csa_tree_add_51_79_groupi_n_11084);
  or csa_tree_add_51_79_groupi_g34956__7410(csa_tree_add_51_79_groupi_n_11101 ,csa_tree_add_51_79_groupi_n_11041 ,csa_tree_add_51_79_groupi_n_11064);
  or csa_tree_add_51_79_groupi_g34957__6417(csa_tree_add_51_79_groupi_n_11100 ,csa_tree_add_51_79_groupi_n_11053 ,csa_tree_add_51_79_groupi_n_11066);
  nor csa_tree_add_51_79_groupi_g34958__5477(csa_tree_add_51_79_groupi_n_11099 ,csa_tree_add_51_79_groupi_n_11052 ,csa_tree_add_51_79_groupi_n_11067);
  or csa_tree_add_51_79_groupi_g34959__2398(csa_tree_add_51_79_groupi_n_11112 ,csa_tree_add_51_79_groupi_n_11011 ,csa_tree_add_51_79_groupi_n_11072);
  and csa_tree_add_51_79_groupi_g34960__5107(csa_tree_add_51_79_groupi_n_11110 ,csa_tree_add_51_79_groupi_n_11048 ,csa_tree_add_51_79_groupi_n_11071);
  not csa_tree_add_51_79_groupi_g34961(csa_tree_add_51_79_groupi_n_11097 ,csa_tree_add_51_79_groupi_n_11096);
  not csa_tree_add_51_79_groupi_g34962(csa_tree_add_51_79_groupi_n_11095 ,csa_tree_add_51_79_groupi_n_11094);
  or csa_tree_add_51_79_groupi_g34963__6260(csa_tree_add_51_79_groupi_n_11093 ,csa_tree_add_51_79_groupi_n_11069 ,csa_tree_add_51_79_groupi_n_10954);
  or csa_tree_add_51_79_groupi_g34964__4319(csa_tree_add_51_79_groupi_n_11092 ,csa_tree_add_51_79_groupi_n_11061 ,csa_tree_add_51_79_groupi_n_11042);
  and csa_tree_add_51_79_groupi_g34965__8428(csa_tree_add_51_79_groupi_n_11091 ,csa_tree_add_51_79_groupi_n_11083 ,csa_tree_add_51_79_groupi_n_11068);
  and csa_tree_add_51_79_groupi_g34966__5526(csa_tree_add_51_79_groupi_n_11090 ,csa_tree_add_51_79_groupi_n_11069 ,csa_tree_add_51_79_groupi_n_10954);
  xnor csa_tree_add_51_79_groupi_g34967__6783(csa_tree_add_51_79_groupi_n_11089 ,csa_tree_add_51_79_groupi_n_11051 ,csa_tree_add_51_79_groupi_n_11005);
  xnor csa_tree_add_51_79_groupi_g34968__3680(csa_tree_add_51_79_groupi_n_11088 ,csa_tree_add_51_79_groupi_n_11050 ,csa_tree_add_51_79_groupi_n_11002);
  xnor csa_tree_add_51_79_groupi_g34969__1617(csa_tree_add_51_79_groupi_n_11087 ,csa_tree_add_51_79_groupi_n_11037 ,csa_tree_add_51_79_groupi_n_11024);
  xnor csa_tree_add_51_79_groupi_g34970__2802(csa_tree_add_51_79_groupi_n_11086 ,csa_tree_add_51_79_groupi_n_11054 ,csa_tree_add_51_79_groupi_n_11041);
  xnor csa_tree_add_51_79_groupi_g34971__1705(csa_tree_add_51_79_groupi_n_11085 ,csa_tree_add_51_79_groupi_n_10953 ,csa_tree_add_51_79_groupi_n_11039);
  xnor csa_tree_add_51_79_groupi_g34972__5122(csa_tree_add_51_79_groupi_n_11098 ,csa_tree_add_51_79_groupi_n_10963 ,csa_tree_add_51_79_groupi_n_11029);
  xnor csa_tree_add_51_79_groupi_g34973__8246(csa_tree_add_51_79_groupi_n_11096 ,csa_tree_add_51_79_groupi_n_11025 ,csa_tree_add_51_79_groupi_n_11028);
  xnor csa_tree_add_51_79_groupi_g34974__7098(csa_tree_add_51_79_groupi_n_11094 ,csa_tree_add_51_79_groupi_n_39 ,csa_tree_add_51_79_groupi_n_11030);
  not csa_tree_add_51_79_groupi_g34975(csa_tree_add_51_79_groupi_n_11081 ,csa_tree_add_51_79_groupi_n_11082);
  not csa_tree_add_51_79_groupi_g34976(csa_tree_add_51_79_groupi_n_11079 ,csa_tree_add_51_79_groupi_n_11080);
  or csa_tree_add_51_79_groupi_g34977__6131(csa_tree_add_51_79_groupi_n_11078 ,csa_tree_add_51_79_groupi_n_11050 ,csa_tree_add_51_79_groupi_n_11001);
  nor csa_tree_add_51_79_groupi_g34978__1881(csa_tree_add_51_79_groupi_n_11077 ,csa_tree_add_51_79_groupi_n_11036 ,csa_tree_add_51_79_groupi_n_11024);
  and csa_tree_add_51_79_groupi_g34979__5115(csa_tree_add_51_79_groupi_n_11076 ,csa_tree_add_51_79_groupi_n_11005 ,csa_tree_add_51_79_groupi_n_11051);
  or csa_tree_add_51_79_groupi_g34980__7482(csa_tree_add_51_79_groupi_n_11075 ,csa_tree_add_51_79_groupi_n_11005 ,csa_tree_add_51_79_groupi_n_11051);
  or csa_tree_add_51_79_groupi_g34981__4733(csa_tree_add_51_79_groupi_n_11074 ,csa_tree_add_51_79_groupi_n_11037 ,csa_tree_add_51_79_groupi_n_11023);
  nor csa_tree_add_51_79_groupi_g34982__6161(csa_tree_add_51_79_groupi_n_11073 ,csa_tree_add_51_79_groupi_n_11049 ,csa_tree_add_51_79_groupi_n_11002);
  nor csa_tree_add_51_79_groupi_g34983__9315(csa_tree_add_51_79_groupi_n_11072 ,csa_tree_add_51_79_groupi_n_11015 ,csa_tree_add_51_79_groupi_n_39);
  or csa_tree_add_51_79_groupi_g34984__9945(csa_tree_add_51_79_groupi_n_11071 ,csa_tree_add_51_79_groupi_n_11045 ,csa_tree_add_51_79_groupi_n_11055);
  and csa_tree_add_51_79_groupi_g34985__2883(csa_tree_add_51_79_groupi_n_11084 ,csa_tree_add_51_79_groupi_n_10979 ,csa_tree_add_51_79_groupi_n_11044);
  and csa_tree_add_51_79_groupi_g34986__2346(csa_tree_add_51_79_groupi_n_11083 ,csa_tree_add_51_79_groupi_n_11043 ,csa_tree_add_51_79_groupi_n_11012);
  or csa_tree_add_51_79_groupi_g34987__1666(csa_tree_add_51_79_groupi_n_11082 ,csa_tree_add_51_79_groupi_n_11021 ,csa_tree_add_51_79_groupi_n_11047);
  and csa_tree_add_51_79_groupi_g34988__7410(csa_tree_add_51_79_groupi_n_11080 ,csa_tree_add_51_79_groupi_n_10947 ,csa_tree_add_51_79_groupi_n_11035);
  not csa_tree_add_51_79_groupi_g34989(csa_tree_add_51_79_groupi_n_11068 ,csa_tree_add_51_79_groupi_n_41);
  not csa_tree_add_51_79_groupi_g34990(csa_tree_add_51_79_groupi_n_11067 ,csa_tree_add_51_79_groupi_n_11066);
  not csa_tree_add_51_79_groupi_g34991(csa_tree_add_51_79_groupi_n_11065 ,csa_tree_add_51_79_groupi_n_11064);
  not csa_tree_add_51_79_groupi_g34992(csa_tree_add_51_79_groupi_n_11063 ,csa_tree_add_51_79_groupi_n_42);
  xnor csa_tree_add_51_79_groupi_g34993__6417(out1[6] ,csa_tree_add_51_79_groupi_n_11027 ,csa_tree_add_51_79_groupi_n_10995);
  nor csa_tree_add_51_79_groupi_g34994__5477(csa_tree_add_51_79_groupi_n_11061 ,csa_tree_add_51_79_groupi_n_10953 ,csa_tree_add_51_79_groupi_n_11039);
  or csa_tree_add_51_79_groupi_g34995__2398(csa_tree_add_51_79_groupi_n_11060 ,csa_tree_add_51_79_groupi_n_10952 ,csa_tree_add_51_79_groupi_n_11038);
  xnor csa_tree_add_51_79_groupi_g34996__5107(csa_tree_add_51_79_groupi_n_11059 ,csa_tree_add_51_79_groupi_n_10960 ,csa_tree_add_51_79_groupi_n_11004);
  xor csa_tree_add_51_79_groupi_g34997__6260(csa_tree_add_51_79_groupi_n_11058 ,csa_tree_add_51_79_groupi_n_11026 ,csa_tree_add_51_79_groupi_n_10954);
  xnor csa_tree_add_51_79_groupi_g34998__4319(csa_tree_add_51_79_groupi_n_11057 ,csa_tree_add_51_79_groupi_n_11000 ,csa_tree_add_51_79_groupi_n_10913);
  xnor csa_tree_add_51_79_groupi_g34999__8428(csa_tree_add_51_79_groupi_n_11070 ,csa_tree_add_51_79_groupi_n_10966 ,csa_tree_add_51_79_groupi_n_10993);
  xnor csa_tree_add_51_79_groupi_g35000__5526(csa_tree_add_51_79_groupi_n_11069 ,csa_tree_add_51_79_groupi_n_10905 ,csa_tree_add_51_79_groupi_n_10990);
  xnor csa_tree_add_51_79_groupi_g35002__6783(csa_tree_add_51_79_groupi_n_11066 ,csa_tree_add_51_79_groupi_n_11008 ,csa_tree_add_51_79_groupi_n_10992);
  xnor csa_tree_add_51_79_groupi_g35003__3680(csa_tree_add_51_79_groupi_n_11064 ,csa_tree_add_51_79_groupi_n_10938 ,csa_tree_add_51_79_groupi_n_10991);
  not csa_tree_add_51_79_groupi_g35005(csa_tree_add_51_79_groupi_n_11053 ,csa_tree_add_51_79_groupi_n_11052);
  not csa_tree_add_51_79_groupi_g35006(csa_tree_add_51_79_groupi_n_11049 ,csa_tree_add_51_79_groupi_n_11050);
  or csa_tree_add_51_79_groupi_g35007__1617(csa_tree_add_51_79_groupi_n_11048 ,csa_tree_add_51_79_groupi_n_40 ,csa_tree_add_51_79_groupi_n_10912);
  nor csa_tree_add_51_79_groupi_g35008__2802(csa_tree_add_51_79_groupi_n_11047 ,csa_tree_add_51_79_groupi_n_10988 ,csa_tree_add_51_79_groupi_n_11020);
  nor csa_tree_add_51_79_groupi_g35009__1705(csa_tree_add_51_79_groupi_n_11046 ,csa_tree_add_51_79_groupi_n_10959 ,csa_tree_add_51_79_groupi_n_11004);
  nor csa_tree_add_51_79_groupi_g35010__5122(csa_tree_add_51_79_groupi_n_11045 ,csa_tree_add_51_79_groupi_n_11000 ,csa_tree_add_51_79_groupi_n_10913);
  or csa_tree_add_51_79_groupi_g35011__8246(csa_tree_add_51_79_groupi_n_11044 ,csa_tree_add_51_79_groupi_n_10978 ,csa_tree_add_51_79_groupi_n_11027);
  or csa_tree_add_51_79_groupi_g35012__7098(csa_tree_add_51_79_groupi_n_11043 ,csa_tree_add_51_79_groupi_n_11014 ,csa_tree_add_51_79_groupi_n_11025);
  and csa_tree_add_51_79_groupi_g35013__6131(csa_tree_add_51_79_groupi_n_11056 ,csa_tree_add_51_79_groupi_n_10982 ,csa_tree_add_51_79_groupi_n_11022);
  and csa_tree_add_51_79_groupi_g35014__1881(csa_tree_add_51_79_groupi_n_11055 ,csa_tree_add_51_79_groupi_n_10923 ,csa_tree_add_51_79_groupi_n_11017);
  and csa_tree_add_51_79_groupi_g35015__5115(csa_tree_add_51_79_groupi_n_11054 ,csa_tree_add_51_79_groupi_n_11018 ,csa_tree_add_51_79_groupi_n_10973);
  or csa_tree_add_51_79_groupi_g35016__7482(csa_tree_add_51_79_groupi_n_11052 ,csa_tree_add_51_79_groupi_n_11016 ,csa_tree_add_51_79_groupi_n_10925);
  and csa_tree_add_51_79_groupi_g35017__4733(csa_tree_add_51_79_groupi_n_11051 ,csa_tree_add_51_79_groupi_n_10969 ,csa_tree_add_51_79_groupi_n_11019);
  and csa_tree_add_51_79_groupi_g35018__6161(csa_tree_add_51_79_groupi_n_11050 ,csa_tree_add_51_79_groupi_n_11013 ,csa_tree_add_51_79_groupi_n_10972);
  not csa_tree_add_51_79_groupi_g35020(csa_tree_add_51_79_groupi_n_11041 ,csa_tree_add_51_79_groupi_n_11040);
  not csa_tree_add_51_79_groupi_g35021(csa_tree_add_51_79_groupi_n_11039 ,csa_tree_add_51_79_groupi_n_11038);
  not csa_tree_add_51_79_groupi_g35022(csa_tree_add_51_79_groupi_n_11037 ,csa_tree_add_51_79_groupi_n_11036);
  or csa_tree_add_51_79_groupi_g35023__9315(csa_tree_add_51_79_groupi_n_11035 ,csa_tree_add_51_79_groupi_n_11009 ,csa_tree_add_51_79_groupi_n_10950);
  or csa_tree_add_51_79_groupi_g35024__9945(csa_tree_add_51_79_groupi_n_11034 ,csa_tree_add_51_79_groupi_n_10960 ,csa_tree_add_51_79_groupi_n_11003);
  xnor csa_tree_add_51_79_groupi_g35025__2883(out1[5] ,csa_tree_add_51_79_groupi_n_10887 ,csa_tree_add_51_79_groupi_n_10943);
  xnor csa_tree_add_51_79_groupi_g35026__2346(csa_tree_add_51_79_groupi_n_11032 ,csa_tree_add_51_79_groupi_n_10936 ,csa_tree_add_51_79_groupi_n_10958);
  xnor csa_tree_add_51_79_groupi_g35027__1666(csa_tree_add_51_79_groupi_n_11031 ,csa_tree_add_51_79_groupi_n_10956 ,csa_tree_add_51_79_groupi_n_10909);
  xnor csa_tree_add_51_79_groupi_g35028__7410(csa_tree_add_51_79_groupi_n_11030 ,csa_tree_add_51_79_groupi_n_10965 ,csa_tree_add_51_79_groupi_n_10983);
  xor csa_tree_add_51_79_groupi_g35029__6417(csa_tree_add_51_79_groupi_n_11029 ,csa_tree_add_51_79_groupi_n_10988 ,csa_tree_add_51_79_groupi_n_10883);
  xnor csa_tree_add_51_79_groupi_g35030__5477(csa_tree_add_51_79_groupi_n_11028 ,csa_tree_add_51_79_groupi_n_10962 ,csa_tree_add_51_79_groupi_n_10928);
  and csa_tree_add_51_79_groupi_g35031__2398(csa_tree_add_51_79_groupi_n_11042 ,csa_tree_add_51_79_groupi_n_10951 ,csa_tree_add_51_79_groupi_n_10999);
  xnor csa_tree_add_51_79_groupi_g35033__5107(csa_tree_add_51_79_groupi_n_11040 ,csa_tree_add_51_79_groupi_n_10791 ,csa_tree_add_51_79_groupi_n_10945);
  xnor csa_tree_add_51_79_groupi_g35034__6260(csa_tree_add_51_79_groupi_n_11038 ,csa_tree_add_51_79_groupi_n_10986 ,csa_tree_add_51_79_groupi_n_10946);
  xnor csa_tree_add_51_79_groupi_g35035__4319(csa_tree_add_51_79_groupi_n_11036 ,csa_tree_add_51_79_groupi_n_10967 ,csa_tree_add_51_79_groupi_n_10942);
  not csa_tree_add_51_79_groupi_g35036(csa_tree_add_51_79_groupi_n_11024 ,csa_tree_add_51_79_groupi_n_11023);
  or csa_tree_add_51_79_groupi_g35037__8428(csa_tree_add_51_79_groupi_n_11022 ,csa_tree_add_51_79_groupi_n_10981 ,csa_tree_add_51_79_groupi_n_10966);
  nor csa_tree_add_51_79_groupi_g35038__5526(csa_tree_add_51_79_groupi_n_11021 ,csa_tree_add_51_79_groupi_n_10883 ,csa_tree_add_51_79_groupi_n_10964);
  and csa_tree_add_51_79_groupi_g35039__6783(csa_tree_add_51_79_groupi_n_11020 ,csa_tree_add_51_79_groupi_n_10883 ,csa_tree_add_51_79_groupi_n_10964);
  or csa_tree_add_51_79_groupi_g35040__3680(csa_tree_add_51_79_groupi_n_11019 ,csa_tree_add_51_79_groupi_n_10938 ,csa_tree_add_51_79_groupi_n_10968);
  or csa_tree_add_51_79_groupi_g35041__1617(csa_tree_add_51_79_groupi_n_11018 ,csa_tree_add_51_79_groupi_n_10971 ,csa_tree_add_51_79_groupi_n_10941);
  or csa_tree_add_51_79_groupi_g35042__2802(csa_tree_add_51_79_groupi_n_11017 ,csa_tree_add_51_79_groupi_n_10893 ,csa_tree_add_51_79_groupi_n_10986);
  and csa_tree_add_51_79_groupi_g35043__1705(csa_tree_add_51_79_groupi_n_11016 ,csa_tree_add_51_79_groupi_n_10967 ,csa_tree_add_51_79_groupi_n_10924);
  nor csa_tree_add_51_79_groupi_g35044__5122(csa_tree_add_51_79_groupi_n_11015 ,csa_tree_add_51_79_groupi_n_10965 ,csa_tree_add_51_79_groupi_n_10983);
  nor csa_tree_add_51_79_groupi_g35045__8246(csa_tree_add_51_79_groupi_n_11014 ,csa_tree_add_51_79_groupi_n_10962 ,csa_tree_add_51_79_groupi_n_10928);
  or csa_tree_add_51_79_groupi_g35046__7098(csa_tree_add_51_79_groupi_n_11013 ,csa_tree_add_51_79_groupi_n_10976 ,csa_tree_add_51_79_groupi_n_10940);
  or csa_tree_add_51_79_groupi_g35047__6131(csa_tree_add_51_79_groupi_n_11012 ,csa_tree_add_51_79_groupi_n_10961 ,csa_tree_add_51_79_groupi_n_10927);
  and csa_tree_add_51_79_groupi_g35048__1881(csa_tree_add_51_79_groupi_n_11011 ,csa_tree_add_51_79_groupi_n_10965 ,csa_tree_add_51_79_groupi_n_10983);
  nor csa_tree_add_51_79_groupi_g35049__5115(csa_tree_add_51_79_groupi_n_11010 ,csa_tree_add_51_79_groupi_n_10955 ,csa_tree_add_51_79_groupi_n_10909);
  and csa_tree_add_51_79_groupi_g35050__7482(csa_tree_add_51_79_groupi_n_11027 ,csa_tree_add_51_79_groupi_n_10977 ,csa_tree_add_51_79_groupi_n_10896);
  and csa_tree_add_51_79_groupi_g35051__4733(csa_tree_add_51_79_groupi_n_11026 ,csa_tree_add_51_79_groupi_n_10974 ,csa_tree_add_51_79_groupi_n_10926);
  and csa_tree_add_51_79_groupi_g35052__6161(csa_tree_add_51_79_groupi_n_11025 ,csa_tree_add_51_79_groupi_n_10866 ,csa_tree_add_51_79_groupi_n_10975);
  and csa_tree_add_51_79_groupi_g35053__9315(csa_tree_add_51_79_groupi_n_11023 ,csa_tree_add_51_79_groupi_n_10875 ,csa_tree_add_51_79_groupi_n_10980);
  not csa_tree_add_51_79_groupi_g35054(csa_tree_add_51_79_groupi_n_11009 ,csa_tree_add_51_79_groupi_n_11008);
  not csa_tree_add_51_79_groupi_g35055(csa_tree_add_51_79_groupi_n_11007 ,csa_tree_add_51_79_groupi_n_11006);
  not csa_tree_add_51_79_groupi_g35056(csa_tree_add_51_79_groupi_n_11004 ,csa_tree_add_51_79_groupi_n_11003);
  not csa_tree_add_51_79_groupi_g35057(csa_tree_add_51_79_groupi_n_11002 ,csa_tree_add_51_79_groupi_n_11001);
  not csa_tree_add_51_79_groupi_g35058(csa_tree_add_51_79_groupi_n_11000 ,csa_tree_add_51_79_groupi_n_40);
  or csa_tree_add_51_79_groupi_g35059__9945(csa_tree_add_51_79_groupi_n_10999 ,csa_tree_add_51_79_groupi_n_10948 ,csa_tree_add_51_79_groupi_n_10987);
  or csa_tree_add_51_79_groupi_g35060__2883(csa_tree_add_51_79_groupi_n_10998 ,csa_tree_add_51_79_groupi_n_10956 ,csa_tree_add_51_79_groupi_n_10908);
  nor csa_tree_add_51_79_groupi_g35061__2346(csa_tree_add_51_79_groupi_n_10997 ,csa_tree_add_51_79_groupi_n_10935 ,csa_tree_add_51_79_groupi_n_10958);
  or csa_tree_add_51_79_groupi_g35062__1666(csa_tree_add_51_79_groupi_n_10996 ,csa_tree_add_51_79_groupi_n_10936 ,csa_tree_add_51_79_groupi_n_10957);
  xnor csa_tree_add_51_79_groupi_g35063__7410(csa_tree_add_51_79_groupi_n_10995 ,csa_tree_add_51_79_groupi_n_10830 ,csa_tree_add_51_79_groupi_n_10907);
  xnor csa_tree_add_51_79_groupi_g35065__6417(csa_tree_add_51_79_groupi_n_10994 ,csa_tree_add_51_79_groupi_n_10934 ,csa_tree_add_51_79_groupi_n_10901);
  xnor csa_tree_add_51_79_groupi_g35066__5477(csa_tree_add_51_79_groupi_n_10993 ,csa_tree_add_51_79_groupi_n_10930 ,csa_tree_add_51_79_groupi_n_10899);
  xnor csa_tree_add_51_79_groupi_g35067__2398(csa_tree_add_51_79_groupi_n_10992 ,csa_tree_add_51_79_groupi_n_10932 ,csa_tree_add_51_79_groupi_n_10911);
  xnor csa_tree_add_51_79_groupi_g35068__5107(csa_tree_add_51_79_groupi_n_10991 ,csa_tree_add_51_79_groupi_n_10903 ,csa_tree_add_51_79_groupi_n_10886);
  xnor csa_tree_add_51_79_groupi_g35069__6260(csa_tree_add_51_79_groupi_n_10990 ,csa_tree_add_51_79_groupi_n_10797 ,csa_tree_add_51_79_groupi_n_10941);
  xnor csa_tree_add_51_79_groupi_g35070__4319(csa_tree_add_51_79_groupi_n_10989 ,csa_tree_add_51_79_groupi_n_10855 ,csa_tree_add_51_79_groupi_n_10915);
  xnor csa_tree_add_51_79_groupi_g35071__8428(csa_tree_add_51_79_groupi_n_11008 ,csa_tree_add_51_79_groupi_n_10831 ,csa_tree_add_51_79_groupi_n_36);
  xnor csa_tree_add_51_79_groupi_g35072__5526(csa_tree_add_51_79_groupi_n_11006 ,csa_tree_add_51_79_groupi_n_10795 ,csa_tree_add_51_79_groupi_n_10892);
  xnor csa_tree_add_51_79_groupi_g35073__6783(csa_tree_add_51_79_groupi_n_11005 ,csa_tree_add_51_79_groupi_n_10786 ,csa_tree_add_51_79_groupi_n_10891);
  xnor csa_tree_add_51_79_groupi_g35074__3680(csa_tree_add_51_79_groupi_n_11003 ,csa_tree_add_51_79_groupi_n_10916 ,csa_tree_add_51_79_groupi_n_10890);
  xnor csa_tree_add_51_79_groupi_g35075__1617(csa_tree_add_51_79_groupi_n_11001 ,csa_tree_add_51_79_groupi_n_10888 ,csa_tree_add_51_79_groupi_n_10889);
  not csa_tree_add_51_79_groupi_g35078(csa_tree_add_51_79_groupi_n_10984 ,csa_tree_add_51_79_groupi_n_10985);
  or csa_tree_add_51_79_groupi_g35079__2802(csa_tree_add_51_79_groupi_n_10982 ,csa_tree_add_51_79_groupi_n_10899 ,csa_tree_add_51_79_groupi_n_10930);
  and csa_tree_add_51_79_groupi_g35080__1705(csa_tree_add_51_79_groupi_n_10981 ,csa_tree_add_51_79_groupi_n_10899 ,csa_tree_add_51_79_groupi_n_10930);
  or csa_tree_add_51_79_groupi_g35081__5122(csa_tree_add_51_79_groupi_n_10980 ,csa_tree_add_51_79_groupi_n_10874 ,csa_tree_add_51_79_groupi_n_10916);
  or csa_tree_add_51_79_groupi_g35082__8246(csa_tree_add_51_79_groupi_n_10979 ,csa_tree_add_51_79_groupi_n_10830 ,csa_tree_add_51_79_groupi_n_10906);
  nor csa_tree_add_51_79_groupi_g35083__7098(csa_tree_add_51_79_groupi_n_10978 ,csa_tree_add_51_79_groupi_n_10829 ,csa_tree_add_51_79_groupi_n_10907);
  or csa_tree_add_51_79_groupi_g35084__6131(csa_tree_add_51_79_groupi_n_10977 ,csa_tree_add_51_79_groupi_n_10898 ,csa_tree_add_51_79_groupi_n_10887);
  nor csa_tree_add_51_79_groupi_g35085__1881(csa_tree_add_51_79_groupi_n_10976 ,csa_tree_add_51_79_groupi_n_10855 ,csa_tree_add_51_79_groupi_n_10915);
  or csa_tree_add_51_79_groupi_g35086__5115(csa_tree_add_51_79_groupi_n_10975 ,csa_tree_add_51_79_groupi_n_10939 ,csa_tree_add_51_79_groupi_n_10849);
  or csa_tree_add_51_79_groupi_g35087__7482(csa_tree_add_51_79_groupi_n_10974 ,csa_tree_add_51_79_groupi_n_10920 ,csa_tree_add_51_79_groupi_n_10937);
  or csa_tree_add_51_79_groupi_g35088__4733(csa_tree_add_51_79_groupi_n_10973 ,csa_tree_add_51_79_groupi_n_10796 ,csa_tree_add_51_79_groupi_n_10904);
  or csa_tree_add_51_79_groupi_g35089__6161(csa_tree_add_51_79_groupi_n_10972 ,csa_tree_add_51_79_groupi_n_10854 ,csa_tree_add_51_79_groupi_n_10914);
  nor csa_tree_add_51_79_groupi_g35090__9315(csa_tree_add_51_79_groupi_n_10971 ,csa_tree_add_51_79_groupi_n_10797 ,csa_tree_add_51_79_groupi_n_10905);
  or csa_tree_add_51_79_groupi_g35091__9945(csa_tree_add_51_79_groupi_n_10970 ,csa_tree_add_51_79_groupi_n_10721 ,csa_tree_add_51_79_groupi_n_10929);
  or csa_tree_add_51_79_groupi_g35092__2883(csa_tree_add_51_79_groupi_n_10969 ,csa_tree_add_51_79_groupi_n_10902 ,csa_tree_add_51_79_groupi_n_10885);
  nor csa_tree_add_51_79_groupi_g35093__2346(csa_tree_add_51_79_groupi_n_10968 ,csa_tree_add_51_79_groupi_n_10903 ,csa_tree_add_51_79_groupi_n_10886);
  and csa_tree_add_51_79_groupi_g35094__1666(csa_tree_add_51_79_groupi_n_10988 ,csa_tree_add_51_79_groupi_n_10921 ,csa_tree_add_51_79_groupi_n_10870);
  and csa_tree_add_51_79_groupi_g35095__7410(csa_tree_add_51_79_groupi_n_10987 ,csa_tree_add_51_79_groupi_n_10922 ,csa_tree_add_51_79_groupi_n_10808);
  and csa_tree_add_51_79_groupi_g35096__6417(csa_tree_add_51_79_groupi_n_10986 ,csa_tree_add_51_79_groupi_n_10845 ,csa_tree_add_51_79_groupi_n_10897);
  and csa_tree_add_51_79_groupi_g35097__5477(csa_tree_add_51_79_groupi_n_10985 ,csa_tree_add_51_79_groupi_n_10917 ,csa_tree_add_51_79_groupi_n_10865);
  or csa_tree_add_51_79_groupi_g35098__2398(csa_tree_add_51_79_groupi_n_10983 ,csa_tree_add_51_79_groupi_n_10869 ,csa_tree_add_51_79_groupi_n_10918);
  not csa_tree_add_51_79_groupi_g35099(csa_tree_add_51_79_groupi_n_10964 ,csa_tree_add_51_79_groupi_n_10963);
  not csa_tree_add_51_79_groupi_g35100(csa_tree_add_51_79_groupi_n_10962 ,csa_tree_add_51_79_groupi_n_10961);
  not csa_tree_add_51_79_groupi_g35101(csa_tree_add_51_79_groupi_n_10960 ,csa_tree_add_51_79_groupi_n_10959);
  not csa_tree_add_51_79_groupi_g35102(csa_tree_add_51_79_groupi_n_10958 ,csa_tree_add_51_79_groupi_n_10957);
  not csa_tree_add_51_79_groupi_g35103(csa_tree_add_51_79_groupi_n_10956 ,csa_tree_add_51_79_groupi_n_10955);
  not csa_tree_add_51_79_groupi_g35104(csa_tree_add_51_79_groupi_n_10953 ,csa_tree_add_51_79_groupi_n_10952);
  or csa_tree_add_51_79_groupi_g35105__5107(csa_tree_add_51_79_groupi_n_10951 ,csa_tree_add_51_79_groupi_n_10934 ,csa_tree_add_51_79_groupi_n_10900);
  nor csa_tree_add_51_79_groupi_g35106__6260(csa_tree_add_51_79_groupi_n_10950 ,csa_tree_add_51_79_groupi_n_10931 ,csa_tree_add_51_79_groupi_n_10911);
  and csa_tree_add_51_79_groupi_g35107__4319(csa_tree_add_51_79_groupi_n_10949 ,csa_tree_add_51_79_groupi_n_10721 ,csa_tree_add_51_79_groupi_n_10929);
  nor csa_tree_add_51_79_groupi_g35108__8428(csa_tree_add_51_79_groupi_n_10948 ,csa_tree_add_51_79_groupi_n_10933 ,csa_tree_add_51_79_groupi_n_10901);
  or csa_tree_add_51_79_groupi_g35109__5526(csa_tree_add_51_79_groupi_n_10947 ,csa_tree_add_51_79_groupi_n_10932 ,csa_tree_add_51_79_groupi_n_10910);
  xnor csa_tree_add_51_79_groupi_g35110__6783(csa_tree_add_51_79_groupi_n_10946 ,csa_tree_add_51_79_groupi_n_10799 ,csa_tree_add_51_79_groupi_n_10853);
  xnor csa_tree_add_51_79_groupi_g35111__3680(csa_tree_add_51_79_groupi_n_10945 ,csa_tree_add_51_79_groupi_n_10861 ,csa_tree_add_51_79_groupi_n_10647);
  xnor csa_tree_add_51_79_groupi_g35112__1617(csa_tree_add_51_79_groupi_n_10944 ,csa_tree_add_51_79_groupi_n_10784 ,csa_tree_add_51_79_groupi_n_10859);
  xnor csa_tree_add_51_79_groupi_g35113__2802(csa_tree_add_51_79_groupi_n_10943 ,csa_tree_add_51_79_groupi_n_10857 ,csa_tree_add_51_79_groupi_n_10686);
  xnor csa_tree_add_51_79_groupi_g35114__1705(csa_tree_add_51_79_groupi_n_10942 ,csa_tree_add_51_79_groupi_n_10884 ,csa_tree_add_51_79_groupi_n_10860);
  xnor csa_tree_add_51_79_groupi_g35115__5122(csa_tree_add_51_79_groupi_n_10967 ,csa_tree_add_51_79_groupi_n_10726 ,csa_tree_add_51_79_groupi_n_35);
  xnor csa_tree_add_51_79_groupi_g35116__8246(csa_tree_add_51_79_groupi_n_10966 ,csa_tree_add_51_79_groupi_n_10862 ,csa_tree_add_51_79_groupi_n_10843);
  xnor csa_tree_add_51_79_groupi_g35117__7098(csa_tree_add_51_79_groupi_n_10965 ,csa_tree_add_51_79_groupi_n_10764 ,csa_tree_add_51_79_groupi_n_10840);
  xnor csa_tree_add_51_79_groupi_g35118__6131(csa_tree_add_51_79_groupi_n_10963 ,csa_tree_add_51_79_groupi_n_10719 ,csa_tree_add_51_79_groupi_n_10839);
  xnor csa_tree_add_51_79_groupi_g35119__1881(csa_tree_add_51_79_groupi_n_10961 ,csa_tree_add_51_79_groupi_n_10802 ,csa_tree_add_51_79_groupi_n_10842);
  or csa_tree_add_51_79_groupi_g35120__5115(csa_tree_add_51_79_groupi_n_10959 ,csa_tree_add_51_79_groupi_n_10777 ,csa_tree_add_51_79_groupi_n_10895);
  xnor csa_tree_add_51_79_groupi_g35121__7482(csa_tree_add_51_79_groupi_n_10957 ,csa_tree_add_51_79_groupi_n_10864 ,csa_tree_add_51_79_groupi_n_10844);
  or csa_tree_add_51_79_groupi_g35122__4733(csa_tree_add_51_79_groupi_n_10955 ,csa_tree_add_51_79_groupi_n_10848 ,csa_tree_add_51_79_groupi_n_10919);
  xnor csa_tree_add_51_79_groupi_g35123__6161(csa_tree_add_51_79_groupi_n_10954 ,csa_tree_add_51_79_groupi_n_10834 ,csa_tree_add_51_79_groupi_n_10841);
  xnor csa_tree_add_51_79_groupi_g35124__9315(csa_tree_add_51_79_groupi_n_10952 ,csa_tree_add_51_79_groupi_n_10727 ,csa_tree_add_51_79_groupi_n_10838);
  not csa_tree_add_51_79_groupi_g35128(csa_tree_add_51_79_groupi_n_10935 ,csa_tree_add_51_79_groupi_n_10936);
  not csa_tree_add_51_79_groupi_g35129(csa_tree_add_51_79_groupi_n_10933 ,csa_tree_add_51_79_groupi_n_10934);
  not csa_tree_add_51_79_groupi_g35130(csa_tree_add_51_79_groupi_n_10931 ,csa_tree_add_51_79_groupi_n_10932);
  not csa_tree_add_51_79_groupi_g35132(csa_tree_add_51_79_groupi_n_10928 ,csa_tree_add_51_79_groupi_n_10927);
  or csa_tree_add_51_79_groupi_g35133__9945(csa_tree_add_51_79_groupi_n_10926 ,csa_tree_add_51_79_groupi_n_10783 ,csa_tree_add_51_79_groupi_n_10859);
  and csa_tree_add_51_79_groupi_g35134__2883(csa_tree_add_51_79_groupi_n_10925 ,csa_tree_add_51_79_groupi_n_10884 ,csa_tree_add_51_79_groupi_n_10860);
  or csa_tree_add_51_79_groupi_g35135__2346(csa_tree_add_51_79_groupi_n_10924 ,csa_tree_add_51_79_groupi_n_10884 ,csa_tree_add_51_79_groupi_n_10860);
  or csa_tree_add_51_79_groupi_g35136__1666(csa_tree_add_51_79_groupi_n_10923 ,csa_tree_add_51_79_groupi_n_10798 ,csa_tree_add_51_79_groupi_n_10852);
  or csa_tree_add_51_79_groupi_g35137__7410(csa_tree_add_51_79_groupi_n_10922 ,csa_tree_add_51_79_groupi_n_10863 ,csa_tree_add_51_79_groupi_n_10809);
  or csa_tree_add_51_79_groupi_g35138__6417(csa_tree_add_51_79_groupi_n_10921 ,csa_tree_add_51_79_groupi_n_10861 ,csa_tree_add_51_79_groupi_n_10871);
  nor csa_tree_add_51_79_groupi_g35139__5477(csa_tree_add_51_79_groupi_n_10920 ,csa_tree_add_51_79_groupi_n_10784 ,csa_tree_add_51_79_groupi_n_10858);
  and csa_tree_add_51_79_groupi_g35140__2398(csa_tree_add_51_79_groupi_n_10919 ,csa_tree_add_51_79_groupi_n_10851 ,csa_tree_add_51_79_groupi_n_10888);
  nor csa_tree_add_51_79_groupi_g35141__5107(csa_tree_add_51_79_groupi_n_10918 ,csa_tree_add_51_79_groupi_n_10868 ,csa_tree_add_51_79_groupi_n_10801);
  or csa_tree_add_51_79_groupi_g35142__6260(csa_tree_add_51_79_groupi_n_10917 ,csa_tree_add_51_79_groupi_n_10867 ,csa_tree_add_51_79_groupi_n_10836);
  and csa_tree_add_51_79_groupi_g35143__4319(csa_tree_add_51_79_groupi_n_10941 ,csa_tree_add_51_79_groupi_n_10807 ,csa_tree_add_51_79_groupi_n_10877);
  and csa_tree_add_51_79_groupi_g35144__8428(csa_tree_add_51_79_groupi_n_10940 ,csa_tree_add_51_79_groupi_n_10880 ,csa_tree_add_51_79_groupi_n_10824);
  and csa_tree_add_51_79_groupi_g35145__5526(csa_tree_add_51_79_groupi_n_10939 ,csa_tree_add_51_79_groupi_n_10850 ,csa_tree_add_51_79_groupi_n_10821);
  and csa_tree_add_51_79_groupi_g35146__6783(csa_tree_add_51_79_groupi_n_10938 ,csa_tree_add_51_79_groupi_n_10878 ,csa_tree_add_51_79_groupi_n_10817);
  and csa_tree_add_51_79_groupi_g35147__3680(csa_tree_add_51_79_groupi_n_10937 ,csa_tree_add_51_79_groupi_n_10879 ,csa_tree_add_51_79_groupi_n_10741);
  and csa_tree_add_51_79_groupi_g35148__1617(csa_tree_add_51_79_groupi_n_10936 ,csa_tree_add_51_79_groupi_n_10740 ,csa_tree_add_51_79_groupi_n_10882);
  and csa_tree_add_51_79_groupi_g35149__2802(csa_tree_add_51_79_groupi_n_10934 ,csa_tree_add_51_79_groupi_n_10872 ,csa_tree_add_51_79_groupi_n_10810);
  and csa_tree_add_51_79_groupi_g35150__1705(csa_tree_add_51_79_groupi_n_10932 ,csa_tree_add_51_79_groupi_n_10846 ,csa_tree_add_51_79_groupi_n_10779);
  and csa_tree_add_51_79_groupi_g35151__5122(csa_tree_add_51_79_groupi_n_10930 ,csa_tree_add_51_79_groupi_n_10881 ,csa_tree_add_51_79_groupi_n_10818);
  and csa_tree_add_51_79_groupi_g35152__8246(csa_tree_add_51_79_groupi_n_10929 ,csa_tree_add_51_79_groupi_n_10876 ,csa_tree_add_51_79_groupi_n_10630);
  and csa_tree_add_51_79_groupi_g35153__7098(csa_tree_add_51_79_groupi_n_10927 ,csa_tree_add_51_79_groupi_n_10826 ,csa_tree_add_51_79_groupi_n_10873);
  not csa_tree_add_51_79_groupi_g35154(csa_tree_add_51_79_groupi_n_10915 ,csa_tree_add_51_79_groupi_n_10914);
  not csa_tree_add_51_79_groupi_g35155(csa_tree_add_51_79_groupi_n_10913 ,csa_tree_add_51_79_groupi_n_10912);
  not csa_tree_add_51_79_groupi_g35156(csa_tree_add_51_79_groupi_n_10911 ,csa_tree_add_51_79_groupi_n_10910);
  not csa_tree_add_51_79_groupi_g35157(csa_tree_add_51_79_groupi_n_10909 ,csa_tree_add_51_79_groupi_n_10908);
  not csa_tree_add_51_79_groupi_g35158(csa_tree_add_51_79_groupi_n_10907 ,csa_tree_add_51_79_groupi_n_10906);
  not csa_tree_add_51_79_groupi_g35159(csa_tree_add_51_79_groupi_n_10905 ,csa_tree_add_51_79_groupi_n_10904);
  not csa_tree_add_51_79_groupi_g35160(csa_tree_add_51_79_groupi_n_10903 ,csa_tree_add_51_79_groupi_n_10902);
  not csa_tree_add_51_79_groupi_g35161(csa_tree_add_51_79_groupi_n_10901 ,csa_tree_add_51_79_groupi_n_10900);
  nor csa_tree_add_51_79_groupi_g35162__6131(csa_tree_add_51_79_groupi_n_10898 ,csa_tree_add_51_79_groupi_n_10856 ,csa_tree_add_51_79_groupi_n_10686);
  or csa_tree_add_51_79_groupi_g35163__1881(csa_tree_add_51_79_groupi_n_10897 ,csa_tree_add_51_79_groupi_n_10805 ,csa_tree_add_51_79_groupi_n_10847);
  or csa_tree_add_51_79_groupi_g35164__5115(csa_tree_add_51_79_groupi_n_10896 ,csa_tree_add_51_79_groupi_n_10857 ,csa_tree_add_51_79_groupi_n_10685);
  nor csa_tree_add_51_79_groupi_g35165__7482(csa_tree_add_51_79_groupi_n_10895 ,csa_tree_add_51_79_groupi_n_10776 ,csa_tree_add_51_79_groupi_n_10864);
  xnor csa_tree_add_51_79_groupi_g35166__4733(out1[4] ,csa_tree_add_51_79_groupi_n_10694 ,csa_tree_add_51_79_groupi_n_10772);
  nor csa_tree_add_51_79_groupi_g35167__6161(csa_tree_add_51_79_groupi_n_10893 ,csa_tree_add_51_79_groupi_n_10799 ,csa_tree_add_51_79_groupi_n_10853);
  xnor csa_tree_add_51_79_groupi_g35168__9315(csa_tree_add_51_79_groupi_n_10892 ,csa_tree_add_51_79_groupi_n_10805 ,csa_tree_add_51_79_groupi_n_10650);
  xnor csa_tree_add_51_79_groupi_g35170__9945(csa_tree_add_51_79_groupi_n_10891 ,csa_tree_add_51_79_groupi_n_10788 ,csa_tree_add_51_79_groupi_n_10836);
  xnor csa_tree_add_51_79_groupi_g35171__2883(csa_tree_add_51_79_groupi_n_10890 ,csa_tree_add_51_79_groupi_n_10800 ,csa_tree_add_51_79_groupi_n_10828);
  xnor csa_tree_add_51_79_groupi_g35173__2346(csa_tree_add_51_79_groupi_n_10889 ,csa_tree_add_51_79_groupi_n_10640 ,csa_tree_add_51_79_groupi_n_10793);
  xnor csa_tree_add_51_79_groupi_g35174__1666(csa_tree_add_51_79_groupi_n_10916 ,csa_tree_add_51_79_groupi_n_10695 ,csa_tree_add_51_79_groupi_n_10769);
  xnor csa_tree_add_51_79_groupi_g35175__7410(csa_tree_add_51_79_groupi_n_10914 ,csa_tree_add_51_79_groupi_n_10730 ,csa_tree_add_51_79_groupi_n_10767);
  xnor csa_tree_add_51_79_groupi_g35176__6417(csa_tree_add_51_79_groupi_n_10912 ,csa_tree_add_51_79_groupi_n_10751 ,csa_tree_add_51_79_groupi_n_10766);
  xnor csa_tree_add_51_79_groupi_g35177__5477(csa_tree_add_51_79_groupi_n_10910 ,csa_tree_add_51_79_groupi_n_10833 ,csa_tree_add_51_79_groupi_n_10774);
  xnor csa_tree_add_51_79_groupi_g35178__2398(csa_tree_add_51_79_groupi_n_10908 ,csa_tree_add_51_79_groupi_n_10835 ,csa_tree_add_51_79_groupi_n_10696);
  xnor csa_tree_add_51_79_groupi_g35179__5107(csa_tree_add_51_79_groupi_n_10906 ,csa_tree_add_51_79_groupi_n_10803 ,csa_tree_add_51_79_groupi_n_10770);
  xnor csa_tree_add_51_79_groupi_g35180__6260(csa_tree_add_51_79_groupi_n_10904 ,csa_tree_add_51_79_groupi_n_10693 ,csa_tree_add_51_79_groupi_n_10768);
  xnor csa_tree_add_51_79_groupi_g35181__4319(csa_tree_add_51_79_groupi_n_10902 ,csa_tree_add_51_79_groupi_n_10765 ,csa_tree_add_51_79_groupi_n_10771);
  xnor csa_tree_add_51_79_groupi_g35182__8428(csa_tree_add_51_79_groupi_n_10900 ,csa_tree_add_51_79_groupi_n_10728 ,csa_tree_add_51_79_groupi_n_10773);
  xnor csa_tree_add_51_79_groupi_g35183__5526(csa_tree_add_51_79_groupi_n_10899 ,csa_tree_add_51_79_groupi_n_10717 ,csa_tree_add_51_79_groupi_n_10775);
  not csa_tree_add_51_79_groupi_g35184(csa_tree_add_51_79_groupi_n_10886 ,csa_tree_add_51_79_groupi_n_10885);
  or csa_tree_add_51_79_groupi_g35185__6783(csa_tree_add_51_79_groupi_n_10882 ,csa_tree_add_51_79_groupi_n_10804 ,csa_tree_add_51_79_groupi_n_10743);
  or csa_tree_add_51_79_groupi_g35186__3680(csa_tree_add_51_79_groupi_n_10881 ,csa_tree_add_51_79_groupi_n_10762 ,csa_tree_add_51_79_groupi_n_10819);
  or csa_tree_add_51_79_groupi_g35187__1617(csa_tree_add_51_79_groupi_n_10880 ,csa_tree_add_51_79_groupi_n_10802 ,csa_tree_add_51_79_groupi_n_10822);
  or csa_tree_add_51_79_groupi_g35188__2802(csa_tree_add_51_79_groupi_n_10879 ,csa_tree_add_51_79_groupi_n_10742 ,csa_tree_add_51_79_groupi_n_10833);
  or csa_tree_add_51_79_groupi_g35189__1705(csa_tree_add_51_79_groupi_n_10878 ,csa_tree_add_51_79_groupi_n_10816 ,csa_tree_add_51_79_groupi_n_10834);
  or csa_tree_add_51_79_groupi_g35190__5122(csa_tree_add_51_79_groupi_n_10877 ,csa_tree_add_51_79_groupi_n_10764 ,csa_tree_add_51_79_groupi_n_10806);
  or csa_tree_add_51_79_groupi_g35191__8246(csa_tree_add_51_79_groupi_n_10876 ,csa_tree_add_51_79_groupi_n_10637 ,csa_tree_add_51_79_groupi_n_10835);
  or csa_tree_add_51_79_groupi_g35192__7098(csa_tree_add_51_79_groupi_n_10875 ,csa_tree_add_51_79_groupi_n_10828 ,csa_tree_add_51_79_groupi_n_10800);
  and csa_tree_add_51_79_groupi_g35193__6131(csa_tree_add_51_79_groupi_n_10874 ,csa_tree_add_51_79_groupi_n_10828 ,csa_tree_add_51_79_groupi_n_10800);
  or csa_tree_add_51_79_groupi_g35194__1881(csa_tree_add_51_79_groupi_n_10873 ,csa_tree_add_51_79_groupi_n_10612 ,csa_tree_add_51_79_groupi_n_10825);
  or csa_tree_add_51_79_groupi_g35195__5115(csa_tree_add_51_79_groupi_n_10872 ,csa_tree_add_51_79_groupi_n_10811 ,csa_tree_add_51_79_groupi_n_10658);
  nor csa_tree_add_51_79_groupi_g35196__7482(csa_tree_add_51_79_groupi_n_10871 ,csa_tree_add_51_79_groupi_n_10646 ,csa_tree_add_51_79_groupi_n_10791);
  or csa_tree_add_51_79_groupi_g35197__4733(csa_tree_add_51_79_groupi_n_10870 ,csa_tree_add_51_79_groupi_n_10647 ,csa_tree_add_51_79_groupi_n_10790);
  nor csa_tree_add_51_79_groupi_g35198__6161(csa_tree_add_51_79_groupi_n_10869 ,csa_tree_add_51_79_groupi_n_10789 ,csa_tree_add_51_79_groupi_n_10831);
  and csa_tree_add_51_79_groupi_g35199__9315(csa_tree_add_51_79_groupi_n_10868 ,csa_tree_add_51_79_groupi_n_10789 ,csa_tree_add_51_79_groupi_n_10831);
  nor csa_tree_add_51_79_groupi_g35200__9945(csa_tree_add_51_79_groupi_n_10867 ,csa_tree_add_51_79_groupi_n_10786 ,csa_tree_add_51_79_groupi_n_10788);
  or csa_tree_add_51_79_groupi_g35201__2883(csa_tree_add_51_79_groupi_n_10866 ,csa_tree_add_51_79_groupi_n_10720 ,csa_tree_add_51_79_groupi_n_10832);
  or csa_tree_add_51_79_groupi_g35202__2346(csa_tree_add_51_79_groupi_n_10865 ,csa_tree_add_51_79_groupi_n_10785 ,csa_tree_add_51_79_groupi_n_10787);
  or csa_tree_add_51_79_groupi_g35203__1666(csa_tree_add_51_79_groupi_n_10888 ,csa_tree_add_51_79_groupi_n_10712 ,csa_tree_add_51_79_groupi_n_10782);
  and csa_tree_add_51_79_groupi_g35204__7410(csa_tree_add_51_79_groupi_n_10887 ,csa_tree_add_51_79_groupi_n_10812 ,csa_tree_add_51_79_groupi_n_10747);
  and csa_tree_add_51_79_groupi_g35205__6417(csa_tree_add_51_79_groupi_n_10885 ,csa_tree_add_51_79_groupi_n_10814 ,csa_tree_add_51_79_groupi_n_10711);
  or csa_tree_add_51_79_groupi_g35206__5477(csa_tree_add_51_79_groupi_n_10884 ,csa_tree_add_51_79_groupi_n_10815 ,csa_tree_add_51_79_groupi_n_10733);
  and csa_tree_add_51_79_groupi_g35207__2398(csa_tree_add_51_79_groupi_n_10883 ,csa_tree_add_51_79_groupi_n_10823 ,csa_tree_add_51_79_groupi_n_10734);
  not csa_tree_add_51_79_groupi_g35208(csa_tree_add_51_79_groupi_n_10863 ,csa_tree_add_51_79_groupi_n_10862);
  not csa_tree_add_51_79_groupi_g35209(csa_tree_add_51_79_groupi_n_10858 ,csa_tree_add_51_79_groupi_n_10859);
  not csa_tree_add_51_79_groupi_g35210(csa_tree_add_51_79_groupi_n_10857 ,csa_tree_add_51_79_groupi_n_10856);
  not csa_tree_add_51_79_groupi_g35211(csa_tree_add_51_79_groupi_n_10854 ,csa_tree_add_51_79_groupi_n_10855);
  not csa_tree_add_51_79_groupi_g35212(csa_tree_add_51_79_groupi_n_10853 ,csa_tree_add_51_79_groupi_n_10852);
  or csa_tree_add_51_79_groupi_g35213__5107(csa_tree_add_51_79_groupi_n_10851 ,csa_tree_add_51_79_groupi_n_10639 ,csa_tree_add_51_79_groupi_n_10793);
  or csa_tree_add_51_79_groupi_g35214__6260(csa_tree_add_51_79_groupi_n_10850 ,csa_tree_add_51_79_groupi_n_10820 ,csa_tree_add_51_79_groupi_n_10727);
  and csa_tree_add_51_79_groupi_g35215__4319(csa_tree_add_51_79_groupi_n_10849 ,csa_tree_add_51_79_groupi_n_10720 ,csa_tree_add_51_79_groupi_n_10832);
  nor csa_tree_add_51_79_groupi_g35216__8428(csa_tree_add_51_79_groupi_n_10848 ,csa_tree_add_51_79_groupi_n_10640 ,csa_tree_add_51_79_groupi_n_10792);
  nor csa_tree_add_51_79_groupi_g35217__5526(csa_tree_add_51_79_groupi_n_10847 ,csa_tree_add_51_79_groupi_n_10794 ,csa_tree_add_51_79_groupi_n_10650);
  or csa_tree_add_51_79_groupi_g35218__6783(csa_tree_add_51_79_groupi_n_10846 ,csa_tree_add_51_79_groupi_n_10780 ,csa_tree_add_51_79_groupi_n_10763);
  or csa_tree_add_51_79_groupi_g35219__3680(csa_tree_add_51_79_groupi_n_10845 ,csa_tree_add_51_79_groupi_n_10795 ,csa_tree_add_51_79_groupi_n_10649);
  xnor csa_tree_add_51_79_groupi_g35220__1617(csa_tree_add_51_79_groupi_n_10844 ,csa_tree_add_51_79_groupi_n_10722 ,csa_tree_add_51_79_groupi_n_10761);
  xnor csa_tree_add_51_79_groupi_g35221__2802(csa_tree_add_51_79_groupi_n_10843 ,csa_tree_add_51_79_groupi_n_10756 ,csa_tree_add_51_79_groupi_n_10753);
  xnor csa_tree_add_51_79_groupi_g35222__1705(csa_tree_add_51_79_groupi_n_10842 ,csa_tree_add_51_79_groupi_n_10610 ,csa_tree_add_51_79_groupi_n_10749);
  xnor csa_tree_add_51_79_groupi_g35223__5122(csa_tree_add_51_79_groupi_n_10841 ,csa_tree_add_51_79_groupi_n_10724 ,csa_tree_add_51_79_groupi_n_10758);
  xnor csa_tree_add_51_79_groupi_g35224__8246(csa_tree_add_51_79_groupi_n_10840 ,csa_tree_add_51_79_groupi_n_10714 ,csa_tree_add_51_79_groupi_n_10760);
  xnor csa_tree_add_51_79_groupi_g35226__7098(csa_tree_add_51_79_groupi_n_10839 ,csa_tree_add_51_79_groupi_n_10609 ,csa_tree_add_51_79_groupi_n_10762);
  xnor csa_tree_add_51_79_groupi_g35227__6131(csa_tree_add_51_79_groupi_n_10838 ,csa_tree_add_51_79_groupi_n_10716 ,csa_tree_add_51_79_groupi_n_10561);
  xnor csa_tree_add_51_79_groupi_g35228__1881(csa_tree_add_51_79_groupi_n_10837 ,csa_tree_add_51_79_groupi_n_10754 ,csa_tree_add_51_79_groupi_n_10268);
  xnor csa_tree_add_51_79_groupi_g35229__5115(csa_tree_add_51_79_groupi_n_10864 ,csa_tree_add_51_79_groupi_n_10575 ,csa_tree_add_51_79_groupi_n_10699);
  xnor csa_tree_add_51_79_groupi_g35230__7482(csa_tree_add_51_79_groupi_n_10862 ,csa_tree_add_51_79_groupi_n_10487 ,csa_tree_add_51_79_groupi_n_10700);
  xnor csa_tree_add_51_79_groupi_g35231__4733(csa_tree_add_51_79_groupi_n_10861 ,csa_tree_add_51_79_groupi_n_10616 ,csa_tree_add_51_79_groupi_n_10697);
  xnor csa_tree_add_51_79_groupi_g35232__6161(csa_tree_add_51_79_groupi_n_10860 ,csa_tree_add_51_79_groupi_n_10614 ,csa_tree_add_51_79_groupi_n_10698);
  xnor csa_tree_add_51_79_groupi_g35233__9315(csa_tree_add_51_79_groupi_n_10859 ,csa_tree_add_51_79_groupi_n_10566 ,csa_tree_add_51_79_groupi_n_10702);
  xnor csa_tree_add_51_79_groupi_g35234__9945(csa_tree_add_51_79_groupi_n_10856 ,csa_tree_add_51_79_groupi_n_10576 ,csa_tree_add_51_79_groupi_n_10701);
  or csa_tree_add_51_79_groupi_g35235__2883(csa_tree_add_51_79_groupi_n_10855 ,csa_tree_add_51_79_groupi_n_10708 ,csa_tree_add_51_79_groupi_n_10781);
  and csa_tree_add_51_79_groupi_g35236__2346(csa_tree_add_51_79_groupi_n_10852 ,csa_tree_add_51_79_groupi_n_10827 ,csa_tree_add_51_79_groupi_n_10705);
  not csa_tree_add_51_79_groupi_g35238(csa_tree_add_51_79_groupi_n_10829 ,csa_tree_add_51_79_groupi_n_10830);
  or csa_tree_add_51_79_groupi_g35239__1666(csa_tree_add_51_79_groupi_n_10827 ,csa_tree_add_51_79_groupi_n_10729 ,csa_tree_add_51_79_groupi_n_10706);
  or csa_tree_add_51_79_groupi_g35240__7410(csa_tree_add_51_79_groupi_n_10826 ,csa_tree_add_51_79_groupi_n_10750 ,csa_tree_add_51_79_groupi_n_10641);
  nor csa_tree_add_51_79_groupi_g35241__6417(csa_tree_add_51_79_groupi_n_10825 ,csa_tree_add_51_79_groupi_n_10751 ,csa_tree_add_51_79_groupi_n_10642);
  or csa_tree_add_51_79_groupi_g35242__5477(csa_tree_add_51_79_groupi_n_10824 ,csa_tree_add_51_79_groupi_n_10749 ,csa_tree_add_51_79_groupi_n_10610);
  or csa_tree_add_51_79_groupi_g35243__2398(csa_tree_add_51_79_groupi_n_10823 ,csa_tree_add_51_79_groupi_n_10735 ,csa_tree_add_51_79_groupi_n_10765);
  and csa_tree_add_51_79_groupi_g35244__5107(csa_tree_add_51_79_groupi_n_10822 ,csa_tree_add_51_79_groupi_n_10749 ,csa_tree_add_51_79_groupi_n_10610);
  or csa_tree_add_51_79_groupi_g35245__6260(csa_tree_add_51_79_groupi_n_10821 ,csa_tree_add_51_79_groupi_n_10715 ,csa_tree_add_51_79_groupi_n_10560);
  nor csa_tree_add_51_79_groupi_g35246__4319(csa_tree_add_51_79_groupi_n_10820 ,csa_tree_add_51_79_groupi_n_10716 ,csa_tree_add_51_79_groupi_n_10561);
  nor csa_tree_add_51_79_groupi_g35247__8428(csa_tree_add_51_79_groupi_n_10819 ,csa_tree_add_51_79_groupi_n_10719 ,csa_tree_add_51_79_groupi_n_10608);
  or csa_tree_add_51_79_groupi_g35248__5526(csa_tree_add_51_79_groupi_n_10818 ,csa_tree_add_51_79_groupi_n_10718 ,csa_tree_add_51_79_groupi_n_10609);
  or csa_tree_add_51_79_groupi_g35249__6783(csa_tree_add_51_79_groupi_n_10817 ,csa_tree_add_51_79_groupi_n_10723 ,csa_tree_add_51_79_groupi_n_10757);
  nor csa_tree_add_51_79_groupi_g35250__3680(csa_tree_add_51_79_groupi_n_10816 ,csa_tree_add_51_79_groupi_n_10724 ,csa_tree_add_51_79_groupi_n_10758);
  nor csa_tree_add_51_79_groupi_g35251__1617(csa_tree_add_51_79_groupi_n_10815 ,csa_tree_add_51_79_groupi_n_10732 ,csa_tree_add_51_79_groupi_n_10695);
  or csa_tree_add_51_79_groupi_g35252__2802(csa_tree_add_51_79_groupi_n_10814 ,csa_tree_add_51_79_groupi_n_10693 ,csa_tree_add_51_79_groupi_n_10748);
  and csa_tree_add_51_79_groupi_g35253__1705(csa_tree_add_51_79_groupi_n_10813 ,csa_tree_add_51_79_groupi_n_10754 ,csa_tree_add_51_79_groupi_n_10269);
  or csa_tree_add_51_79_groupi_g35254__5122(csa_tree_add_51_79_groupi_n_10812 ,csa_tree_add_51_79_groupi_n_10694 ,csa_tree_add_51_79_groupi_n_10745);
  and csa_tree_add_51_79_groupi_g35255__8246(csa_tree_add_51_79_groupi_n_10811 ,csa_tree_add_51_79_groupi_n_10690 ,csa_tree_add_51_79_groupi_n_10717);
  or csa_tree_add_51_79_groupi_g35256__7098(csa_tree_add_51_79_groupi_n_10810 ,csa_tree_add_51_79_groupi_n_10690 ,csa_tree_add_51_79_groupi_n_10717);
  nor csa_tree_add_51_79_groupi_g35257__6131(csa_tree_add_51_79_groupi_n_10809 ,csa_tree_add_51_79_groupi_n_10756 ,csa_tree_add_51_79_groupi_n_10752);
  or csa_tree_add_51_79_groupi_g35258__1881(csa_tree_add_51_79_groupi_n_10808 ,csa_tree_add_51_79_groupi_n_10755 ,csa_tree_add_51_79_groupi_n_10753);
  or csa_tree_add_51_79_groupi_g35259__5115(csa_tree_add_51_79_groupi_n_10807 ,csa_tree_add_51_79_groupi_n_10713 ,csa_tree_add_51_79_groupi_n_10760);
  nor csa_tree_add_51_79_groupi_g35260__7482(csa_tree_add_51_79_groupi_n_10806 ,csa_tree_add_51_79_groupi_n_10714 ,csa_tree_add_51_79_groupi_n_10759);
  and csa_tree_add_51_79_groupi_g35261__4733(csa_tree_add_51_79_groupi_n_10836 ,csa_tree_add_51_79_groupi_n_10736 ,csa_tree_add_51_79_groupi_n_10666);
  and csa_tree_add_51_79_groupi_g35262__6161(csa_tree_add_51_79_groupi_n_10835 ,csa_tree_add_51_79_groupi_n_10636 ,csa_tree_add_51_79_groupi_n_10703);
  and csa_tree_add_51_79_groupi_g35263__9315(csa_tree_add_51_79_groupi_n_10834 ,csa_tree_add_51_79_groupi_n_10671 ,csa_tree_add_51_79_groupi_n_10738);
  and csa_tree_add_51_79_groupi_g35264__9945(csa_tree_add_51_79_groupi_n_10833 ,csa_tree_add_51_79_groupi_n_10737 ,csa_tree_add_51_79_groupi_n_10668);
  and csa_tree_add_51_79_groupi_g35265__2883(csa_tree_add_51_79_groupi_n_10832 ,csa_tree_add_51_79_groupi_n_10746 ,csa_tree_add_51_79_groupi_n_10605);
  and csa_tree_add_51_79_groupi_g35266__2346(csa_tree_add_51_79_groupi_n_10831 ,csa_tree_add_51_79_groupi_n_10661 ,csa_tree_add_51_79_groupi_n_10731);
  and csa_tree_add_51_79_groupi_g35267__1666(csa_tree_add_51_79_groupi_n_10830 ,csa_tree_add_51_79_groupi_n_10672 ,csa_tree_add_51_79_groupi_n_10744);
  and csa_tree_add_51_79_groupi_g35268__7410(csa_tree_add_51_79_groupi_n_10828 ,csa_tree_add_51_79_groupi_n_10739 ,csa_tree_add_51_79_groupi_n_10662);
  not csa_tree_add_51_79_groupi_g35269(csa_tree_add_51_79_groupi_n_10804 ,csa_tree_add_51_79_groupi_n_10803);
  not csa_tree_add_51_79_groupi_g35270(csa_tree_add_51_79_groupi_n_10799 ,csa_tree_add_51_79_groupi_n_10798);
  not csa_tree_add_51_79_groupi_g35271(csa_tree_add_51_79_groupi_n_10797 ,csa_tree_add_51_79_groupi_n_10796);
  not csa_tree_add_51_79_groupi_g35272(csa_tree_add_51_79_groupi_n_10795 ,csa_tree_add_51_79_groupi_n_10794);
  not csa_tree_add_51_79_groupi_g35273(csa_tree_add_51_79_groupi_n_10793 ,csa_tree_add_51_79_groupi_n_10792);
  not csa_tree_add_51_79_groupi_g35274(csa_tree_add_51_79_groupi_n_10791 ,csa_tree_add_51_79_groupi_n_10790);
  not csa_tree_add_51_79_groupi_g35276(csa_tree_add_51_79_groupi_n_10788 ,csa_tree_add_51_79_groupi_n_10787);
  not csa_tree_add_51_79_groupi_g35277(csa_tree_add_51_79_groupi_n_10786 ,csa_tree_add_51_79_groupi_n_10785);
  not csa_tree_add_51_79_groupi_g35278(csa_tree_add_51_79_groupi_n_10784 ,csa_tree_add_51_79_groupi_n_10783);
  nor csa_tree_add_51_79_groupi_g35279__6417(csa_tree_add_51_79_groupi_n_10782 ,csa_tree_add_51_79_groupi_n_10709 ,csa_tree_add_51_79_groupi_n_10730);
  nor csa_tree_add_51_79_groupi_g35280__5477(csa_tree_add_51_79_groupi_n_10781 ,csa_tree_add_51_79_groupi_n_10707 ,csa_tree_add_51_79_groupi_n_10525);
  and csa_tree_add_51_79_groupi_g35281__2398(csa_tree_add_51_79_groupi_n_10780 ,csa_tree_add_51_79_groupi_n_10726 ,csa_tree_add_51_79_groupi_n_10725);
  or csa_tree_add_51_79_groupi_g35282__5107(csa_tree_add_51_79_groupi_n_10779 ,csa_tree_add_51_79_groupi_n_10726 ,csa_tree_add_51_79_groupi_n_10725);
  nor csa_tree_add_51_79_groupi_g35283__6260(csa_tree_add_51_79_groupi_n_10778 ,csa_tree_add_51_79_groupi_n_10754 ,csa_tree_add_51_79_groupi_n_10269);
  and csa_tree_add_51_79_groupi_g35284__4319(csa_tree_add_51_79_groupi_n_10777 ,csa_tree_add_51_79_groupi_n_10722 ,csa_tree_add_51_79_groupi_n_10761);
  nor csa_tree_add_51_79_groupi_g35285__8428(csa_tree_add_51_79_groupi_n_10776 ,csa_tree_add_51_79_groupi_n_10722 ,csa_tree_add_51_79_groupi_n_10761);
  xnor csa_tree_add_51_79_groupi_g35286__5526(csa_tree_add_51_79_groupi_n_10775 ,csa_tree_add_51_79_groupi_n_10658 ,csa_tree_add_51_79_groupi_n_10690);
  xnor csa_tree_add_51_79_groupi_g35287__6783(csa_tree_add_51_79_groupi_n_10774 ,csa_tree_add_51_79_groupi_n_10687 ,csa_tree_add_51_79_groupi_n_10645);
  xnor csa_tree_add_51_79_groupi_g35288__3680(csa_tree_add_51_79_groupi_n_10773 ,csa_tree_add_51_79_groupi_n_10556 ,csa_tree_add_51_79_groupi_n_10684);
  xnor csa_tree_add_51_79_groupi_g35289__1617(csa_tree_add_51_79_groupi_n_10772 ,csa_tree_add_51_79_groupi_n_10331 ,csa_tree_add_51_79_groupi_n_10652);
  xnor csa_tree_add_51_79_groupi_g35290__2802(csa_tree_add_51_79_groupi_n_10771 ,csa_tree_add_51_79_groupi_n_10691 ,csa_tree_add_51_79_groupi_n_10565);
  xnor csa_tree_add_51_79_groupi_g35291__1705(csa_tree_add_51_79_groupi_n_10770 ,csa_tree_add_51_79_groupi_n_10657 ,csa_tree_add_51_79_groupi_n_10689);
  xnor csa_tree_add_51_79_groupi_g35292__5122(csa_tree_add_51_79_groupi_n_10769 ,csa_tree_add_51_79_groupi_n_10464 ,csa_tree_add_51_79_groupi_n_10655);
  xnor csa_tree_add_51_79_groupi_g35293__8246(csa_tree_add_51_79_groupi_n_10768 ,csa_tree_add_51_79_groupi_n_10654 ,csa_tree_add_51_79_groupi_n_10644);
  xnor csa_tree_add_51_79_groupi_g35294__7098(csa_tree_add_51_79_groupi_n_10767 ,csa_tree_add_51_79_groupi_n_10473 ,csa_tree_add_51_79_groupi_n_10638);
  xnor csa_tree_add_51_79_groupi_g35295__6131(csa_tree_add_51_79_groupi_n_10766 ,csa_tree_add_51_79_groupi_n_10612 ,csa_tree_add_51_79_groupi_n_10642);
  and csa_tree_add_51_79_groupi_g35296__1881(csa_tree_add_51_79_groupi_n_10805 ,csa_tree_add_51_79_groupi_n_10632 ,csa_tree_add_51_79_groupi_n_10704);
  xnor csa_tree_add_51_79_groupi_g35297__5115(csa_tree_add_51_79_groupi_n_10803 ,csa_tree_add_51_79_groupi_n_10481 ,csa_tree_add_51_79_groupi_n_34);
  xnor csa_tree_add_51_79_groupi_g35298__7482(csa_tree_add_51_79_groupi_n_10802 ,csa_tree_add_51_79_groupi_n_10648 ,csa_tree_add_51_79_groupi_n_10622);
  xnor csa_tree_add_51_79_groupi_g35299__4733(csa_tree_add_51_79_groupi_n_10801 ,csa_tree_add_51_79_groupi_n_10477 ,csa_tree_add_51_79_groupi_n_10623);
  xnor csa_tree_add_51_79_groupi_g35300__6161(csa_tree_add_51_79_groupi_n_10800 ,csa_tree_add_51_79_groupi_n_10485 ,csa_tree_add_51_79_groupi_n_10619);
  xnor csa_tree_add_51_79_groupi_g35301__9315(csa_tree_add_51_79_groupi_n_10798 ,csa_tree_add_51_79_groupi_n_10692 ,csa_tree_add_51_79_groupi_n_10629);
  xnor csa_tree_add_51_79_groupi_g35302__9945(csa_tree_add_51_79_groupi_n_10796 ,csa_tree_add_51_79_groupi_n_10468 ,csa_tree_add_51_79_groupi_n_10625);
  xnor csa_tree_add_51_79_groupi_g35303__2883(csa_tree_add_51_79_groupi_n_10794 ,csa_tree_add_51_79_groupi_n_10479 ,csa_tree_add_51_79_groupi_n_10621);
  xnor csa_tree_add_51_79_groupi_g35304__2346(csa_tree_add_51_79_groupi_n_10792 ,csa_tree_add_51_79_groupi_n_10574 ,csa_tree_add_51_79_groupi_n_10626);
  xnor csa_tree_add_51_79_groupi_g35305__1666(csa_tree_add_51_79_groupi_n_10790 ,csa_tree_add_51_79_groupi_n_10459 ,csa_tree_add_51_79_groupi_n_10627);
  xnor csa_tree_add_51_79_groupi_g35306__7410(csa_tree_add_51_79_groupi_n_10789 ,csa_tree_add_51_79_groupi_n_10484 ,csa_tree_add_51_79_groupi_n_10618);
  xnor csa_tree_add_51_79_groupi_g35307__6417(csa_tree_add_51_79_groupi_n_10787 ,csa_tree_add_51_79_groupi_n_10457 ,csa_tree_add_51_79_groupi_n_10628);
  xnor csa_tree_add_51_79_groupi_g35308__5477(csa_tree_add_51_79_groupi_n_10785 ,csa_tree_add_51_79_groupi_n_10577 ,csa_tree_add_51_79_groupi_n_10620);
  xnor csa_tree_add_51_79_groupi_g35309__2398(csa_tree_add_51_79_groupi_n_10783 ,csa_tree_add_51_79_groupi_n_10483 ,csa_tree_add_51_79_groupi_n_10624);
  not csa_tree_add_51_79_groupi_g35311(csa_tree_add_51_79_groupi_n_10759 ,csa_tree_add_51_79_groupi_n_10760);
  not csa_tree_add_51_79_groupi_g35312(csa_tree_add_51_79_groupi_n_10758 ,csa_tree_add_51_79_groupi_n_10757);
  not csa_tree_add_51_79_groupi_g35313(csa_tree_add_51_79_groupi_n_10756 ,csa_tree_add_51_79_groupi_n_10755);
  not csa_tree_add_51_79_groupi_g35314(csa_tree_add_51_79_groupi_n_10752 ,csa_tree_add_51_79_groupi_n_10753);
  not csa_tree_add_51_79_groupi_g35315(csa_tree_add_51_79_groupi_n_10750 ,csa_tree_add_51_79_groupi_n_10751);
  nor csa_tree_add_51_79_groupi_g35316__5107(csa_tree_add_51_79_groupi_n_10748 ,csa_tree_add_51_79_groupi_n_10654 ,csa_tree_add_51_79_groupi_n_10644);
  or csa_tree_add_51_79_groupi_g35317__6260(csa_tree_add_51_79_groupi_n_10747 ,csa_tree_add_51_79_groupi_n_10331 ,csa_tree_add_51_79_groupi_n_10651);
  or csa_tree_add_51_79_groupi_g35318__4319(csa_tree_add_51_79_groupi_n_10746 ,csa_tree_add_51_79_groupi_n_10606 ,csa_tree_add_51_79_groupi_n_10692);
  nor csa_tree_add_51_79_groupi_g35319__8428(csa_tree_add_51_79_groupi_n_10745 ,csa_tree_add_51_79_groupi_n_10330 ,csa_tree_add_51_79_groupi_n_10652);
  or csa_tree_add_51_79_groupi_g35320__5526(csa_tree_add_51_79_groupi_n_10744 ,csa_tree_add_51_79_groupi_n_10576 ,csa_tree_add_51_79_groupi_n_10674);
  nor csa_tree_add_51_79_groupi_g35321__6783(csa_tree_add_51_79_groupi_n_10743 ,csa_tree_add_51_79_groupi_n_10657 ,csa_tree_add_51_79_groupi_n_10688);
  and csa_tree_add_51_79_groupi_g35322__3680(csa_tree_add_51_79_groupi_n_10742 ,csa_tree_add_51_79_groupi_n_10645 ,csa_tree_add_51_79_groupi_n_10687);
  or csa_tree_add_51_79_groupi_g35323__1617(csa_tree_add_51_79_groupi_n_10741 ,csa_tree_add_51_79_groupi_n_10645 ,csa_tree_add_51_79_groupi_n_10687);
  or csa_tree_add_51_79_groupi_g35324__2802(csa_tree_add_51_79_groupi_n_10740 ,csa_tree_add_51_79_groupi_n_10656 ,csa_tree_add_51_79_groupi_n_10689);
  or csa_tree_add_51_79_groupi_g35325__1705(csa_tree_add_51_79_groupi_n_10739 ,csa_tree_add_51_79_groupi_n_10575 ,csa_tree_add_51_79_groupi_n_10659);
  or csa_tree_add_51_79_groupi_g35326__5122(csa_tree_add_51_79_groupi_n_10738 ,csa_tree_add_51_79_groupi_n_10613 ,csa_tree_add_51_79_groupi_n_10670);
  or csa_tree_add_51_79_groupi_g35327__8246(csa_tree_add_51_79_groupi_n_10737 ,csa_tree_add_51_79_groupi_n_10433 ,csa_tree_add_51_79_groupi_n_10669);
  or csa_tree_add_51_79_groupi_g35328__7098(csa_tree_add_51_79_groupi_n_10736 ,csa_tree_add_51_79_groupi_n_10616 ,csa_tree_add_51_79_groupi_n_10667);
  and csa_tree_add_51_79_groupi_g35329__6131(csa_tree_add_51_79_groupi_n_10735 ,csa_tree_add_51_79_groupi_n_10565 ,csa_tree_add_51_79_groupi_n_10691);
  or csa_tree_add_51_79_groupi_g35330__1881(csa_tree_add_51_79_groupi_n_10734 ,csa_tree_add_51_79_groupi_n_10565 ,csa_tree_add_51_79_groupi_n_10691);
  nor csa_tree_add_51_79_groupi_g35331__5115(csa_tree_add_51_79_groupi_n_10733 ,csa_tree_add_51_79_groupi_n_10655 ,csa_tree_add_51_79_groupi_n_10464);
  and csa_tree_add_51_79_groupi_g35332__7482(csa_tree_add_51_79_groupi_n_10732 ,csa_tree_add_51_79_groupi_n_10655 ,csa_tree_add_51_79_groupi_n_10464);
  or csa_tree_add_51_79_groupi_g35333__4733(csa_tree_add_51_79_groupi_n_10731 ,csa_tree_add_51_79_groupi_n_10660 ,csa_tree_add_51_79_groupi_n_10615);
  and csa_tree_add_51_79_groupi_g35334__6161(csa_tree_add_51_79_groupi_n_10765 ,csa_tree_add_51_79_groupi_n_10680 ,csa_tree_add_51_79_groupi_n_10554);
  and csa_tree_add_51_79_groupi_g35335__9315(csa_tree_add_51_79_groupi_n_10764 ,csa_tree_add_51_79_groupi_n_10550 ,csa_tree_add_51_79_groupi_n_10663);
  and csa_tree_add_51_79_groupi_g35336__9945(csa_tree_add_51_79_groupi_n_10763 ,csa_tree_add_51_79_groupi_n_10597 ,csa_tree_add_51_79_groupi_n_10676);
  and csa_tree_add_51_79_groupi_g35337__2883(csa_tree_add_51_79_groupi_n_10762 ,csa_tree_add_51_79_groupi_n_10681 ,csa_tree_add_51_79_groupi_n_10599);
  or csa_tree_add_51_79_groupi_g35338__2346(csa_tree_add_51_79_groupi_n_10761 ,csa_tree_add_51_79_groupi_n_10583 ,csa_tree_add_51_79_groupi_n_10665);
  and csa_tree_add_51_79_groupi_g35339__1666(csa_tree_add_51_79_groupi_n_10760 ,csa_tree_add_51_79_groupi_n_10677 ,csa_tree_add_51_79_groupi_n_10600);
  and csa_tree_add_51_79_groupi_g35340__7410(csa_tree_add_51_79_groupi_n_10757 ,csa_tree_add_51_79_groupi_n_10587 ,csa_tree_add_51_79_groupi_n_10664);
  and csa_tree_add_51_79_groupi_g35341__6417(csa_tree_add_51_79_groupi_n_10755 ,csa_tree_add_51_79_groupi_n_10673 ,csa_tree_add_51_79_groupi_n_10592);
  and csa_tree_add_51_79_groupi_g35342__5477(csa_tree_add_51_79_groupi_n_10754 ,csa_tree_add_51_79_groupi_n_10675 ,csa_tree_add_51_79_groupi_n_10362);
  and csa_tree_add_51_79_groupi_g35343__2398(csa_tree_add_51_79_groupi_n_10753 ,csa_tree_add_51_79_groupi_n_10584 ,csa_tree_add_51_79_groupi_n_10679);
  or csa_tree_add_51_79_groupi_g35344__5107(csa_tree_add_51_79_groupi_n_10751 ,csa_tree_add_51_79_groupi_n_10682 ,csa_tree_add_51_79_groupi_n_10604);
  and csa_tree_add_51_79_groupi_g35345__6260(csa_tree_add_51_79_groupi_n_10749 ,csa_tree_add_51_79_groupi_n_10544 ,csa_tree_add_51_79_groupi_n_10678);
  not csa_tree_add_51_79_groupi_g35346(csa_tree_add_51_79_groupi_n_10729 ,csa_tree_add_51_79_groupi_n_10728);
  not csa_tree_add_51_79_groupi_g35347(csa_tree_add_51_79_groupi_n_10724 ,csa_tree_add_51_79_groupi_n_10723);
  not csa_tree_add_51_79_groupi_g35348(csa_tree_add_51_79_groupi_n_10718 ,csa_tree_add_51_79_groupi_n_10719);
  not csa_tree_add_51_79_groupi_g35349(csa_tree_add_51_79_groupi_n_10716 ,csa_tree_add_51_79_groupi_n_10715);
  not csa_tree_add_51_79_groupi_g35350(csa_tree_add_51_79_groupi_n_10714 ,csa_tree_add_51_79_groupi_n_10713);
  and csa_tree_add_51_79_groupi_g35351__4319(csa_tree_add_51_79_groupi_n_10712 ,csa_tree_add_51_79_groupi_n_10473 ,csa_tree_add_51_79_groupi_n_10638);
  or csa_tree_add_51_79_groupi_g35352__8428(csa_tree_add_51_79_groupi_n_10711 ,csa_tree_add_51_79_groupi_n_10653 ,csa_tree_add_51_79_groupi_n_10643);
  xnor csa_tree_add_51_79_groupi_g35353__5526(out1[3] ,csa_tree_add_51_79_groupi_n_10340 ,csa_tree_add_51_79_groupi_n_10541);
  nor csa_tree_add_51_79_groupi_g35354__6783(csa_tree_add_51_79_groupi_n_10709 ,csa_tree_add_51_79_groupi_n_10473 ,csa_tree_add_51_79_groupi_n_10638);
  and csa_tree_add_51_79_groupi_g35355__3680(csa_tree_add_51_79_groupi_n_10708 ,csa_tree_add_51_79_groupi_n_10482 ,csa_tree_add_51_79_groupi_n_10648);
  nor csa_tree_add_51_79_groupi_g35356__1617(csa_tree_add_51_79_groupi_n_10707 ,csa_tree_add_51_79_groupi_n_10482 ,csa_tree_add_51_79_groupi_n_10648);
  nor csa_tree_add_51_79_groupi_g35357__2802(csa_tree_add_51_79_groupi_n_10706 ,csa_tree_add_51_79_groupi_n_10555 ,csa_tree_add_51_79_groupi_n_10684);
  or csa_tree_add_51_79_groupi_g35358__1705(csa_tree_add_51_79_groupi_n_10705 ,csa_tree_add_51_79_groupi_n_10556 ,csa_tree_add_51_79_groupi_n_10683);
  or csa_tree_add_51_79_groupi_g35359__5122(csa_tree_add_51_79_groupi_n_10704 ,csa_tree_add_51_79_groupi_n_10631 ,csa_tree_add_51_79_groupi_n_10488);
  or csa_tree_add_51_79_groupi_g35360__8246(csa_tree_add_51_79_groupi_n_10703 ,csa_tree_add_51_79_groupi_n_10635 ,csa_tree_add_51_79_groupi_n_10489);
  xnor csa_tree_add_51_79_groupi_g35361__7098(csa_tree_add_51_79_groupi_n_10702 ,csa_tree_add_51_79_groupi_n_10469 ,csa_tree_add_51_79_groupi_n_10613);
  xnor csa_tree_add_51_79_groupi_g35362__6131(csa_tree_add_51_79_groupi_n_10701 ,csa_tree_add_51_79_groupi_n_10572 ,csa_tree_add_51_79_groupi_n_10429);
  xnor csa_tree_add_51_79_groupi_g35363__1881(csa_tree_add_51_79_groupi_n_10700 ,csa_tree_add_51_79_groupi_n_10570 ,csa_tree_add_51_79_groupi_n_10420);
  xnor csa_tree_add_51_79_groupi_g35364__5115(csa_tree_add_51_79_groupi_n_10699 ,csa_tree_add_51_79_groupi_n_10562 ,csa_tree_add_51_79_groupi_n_10611);
  xnor csa_tree_add_51_79_groupi_g35365__7482(csa_tree_add_51_79_groupi_n_10698 ,csa_tree_add_51_79_groupi_n_10517 ,csa_tree_add_51_79_groupi_n_10557);
  xnor csa_tree_add_51_79_groupi_g35366__4733(csa_tree_add_51_79_groupi_n_10697 ,csa_tree_add_51_79_groupi_n_10563 ,csa_tree_add_51_79_groupi_n_10521);
  xnor csa_tree_add_51_79_groupi_g35367__6161(csa_tree_add_51_79_groupi_n_10696 ,csa_tree_add_51_79_groupi_n_10559 ,csa_tree_add_51_79_groupi_n_10568);
  xnor csa_tree_add_51_79_groupi_g35368__9315(csa_tree_add_51_79_groupi_n_10730 ,csa_tree_add_51_79_groupi_n_10387 ,csa_tree_add_51_79_groupi_n_10533);
  or csa_tree_add_51_79_groupi_g35369__9945(csa_tree_add_51_79_groupi_n_10728 ,csa_tree_add_51_79_groupi_n_10546 ,csa_tree_add_51_79_groupi_n_10633);
  and csa_tree_add_51_79_groupi_g35370__2883(csa_tree_add_51_79_groupi_n_10727 ,csa_tree_add_51_79_groupi_n_10634 ,csa_tree_add_51_79_groupi_n_10547);
  xnor csa_tree_add_51_79_groupi_g35371__2346(csa_tree_add_51_79_groupi_n_10726 ,csa_tree_add_51_79_groupi_n_10564 ,csa_tree_add_51_79_groupi_n_10535);
  xnor csa_tree_add_51_79_groupi_g35372__1666(csa_tree_add_51_79_groupi_n_10725 ,csa_tree_add_51_79_groupi_n_10385 ,csa_tree_add_51_79_groupi_n_10542);
  xnor csa_tree_add_51_79_groupi_g35373__7410(csa_tree_add_51_79_groupi_n_10723 ,csa_tree_add_51_79_groupi_n_10436 ,csa_tree_add_51_79_groupi_n_10537);
  xnor csa_tree_add_51_79_groupi_g35374__6417(csa_tree_add_51_79_groupi_n_10722 ,csa_tree_add_51_79_groupi_n_10426 ,csa_tree_add_51_79_groupi_n_10536);
  xnor csa_tree_add_51_79_groupi_g35375__5477(csa_tree_add_51_79_groupi_n_10721 ,csa_tree_add_51_79_groupi_n_10617 ,csa_tree_add_51_79_groupi_n_10448);
  xnor csa_tree_add_51_79_groupi_g35376__2398(csa_tree_add_51_79_groupi_n_10720 ,csa_tree_add_51_79_groupi_n_10470 ,csa_tree_add_51_79_groupi_n_10540);
  xnor csa_tree_add_51_79_groupi_g35377__5107(csa_tree_add_51_79_groupi_n_10719 ,csa_tree_add_51_79_groupi_n_10366 ,csa_tree_add_51_79_groupi_n_10543);
  xnor csa_tree_add_51_79_groupi_g35378__6260(csa_tree_add_51_79_groupi_n_10717 ,csa_tree_add_51_79_groupi_n_10480 ,csa_tree_add_51_79_groupi_n_10538);
  xnor csa_tree_add_51_79_groupi_g35379__4319(csa_tree_add_51_79_groupi_n_10715 ,csa_tree_add_51_79_groupi_n_10466 ,csa_tree_add_51_79_groupi_n_10534);
  xnor csa_tree_add_51_79_groupi_g35380__8428(csa_tree_add_51_79_groupi_n_10713 ,csa_tree_add_51_79_groupi_n_10432 ,csa_tree_add_51_79_groupi_n_10539);
  not csa_tree_add_51_79_groupi_g35381(csa_tree_add_51_79_groupi_n_10688 ,csa_tree_add_51_79_groupi_n_10689);
  not csa_tree_add_51_79_groupi_g35382(csa_tree_add_51_79_groupi_n_10686 ,csa_tree_add_51_79_groupi_n_10685);
  not csa_tree_add_51_79_groupi_g35383(csa_tree_add_51_79_groupi_n_10684 ,csa_tree_add_51_79_groupi_n_10683);
  and csa_tree_add_51_79_groupi_g35384__5526(csa_tree_add_51_79_groupi_n_10682 ,csa_tree_add_51_79_groupi_n_10342 ,csa_tree_add_51_79_groupi_n_10602);
  or csa_tree_add_51_79_groupi_g35385__6783(csa_tree_add_51_79_groupi_n_10681 ,csa_tree_add_51_79_groupi_n_10598 ,csa_tree_add_51_79_groupi_n_10531);
  or csa_tree_add_51_79_groupi_g35386__3680(csa_tree_add_51_79_groupi_n_10680 ,csa_tree_add_51_79_groupi_n_10530 ,csa_tree_add_51_79_groupi_n_10607);
  or csa_tree_add_51_79_groupi_g35387__1617(csa_tree_add_51_79_groupi_n_10679 ,csa_tree_add_51_79_groupi_n_10526 ,csa_tree_add_51_79_groupi_n_10591);
  or csa_tree_add_51_79_groupi_g35388__2802(csa_tree_add_51_79_groupi_n_10678 ,csa_tree_add_51_79_groupi_n_10553 ,csa_tree_add_51_79_groupi_n_10435);
  or csa_tree_add_51_79_groupi_g35389__1705(csa_tree_add_51_79_groupi_n_10677 ,csa_tree_add_51_79_groupi_n_10601 ,csa_tree_add_51_79_groupi_n_10484);
  or csa_tree_add_51_79_groupi_g35390__5122(csa_tree_add_51_79_groupi_n_10676 ,csa_tree_add_51_79_groupi_n_10596 ,csa_tree_add_51_79_groupi_n_10485);
  or csa_tree_add_51_79_groupi_g35391__8246(csa_tree_add_51_79_groupi_n_10675 ,csa_tree_add_51_79_groupi_n_10617 ,csa_tree_add_51_79_groupi_n_10363);
  nor csa_tree_add_51_79_groupi_g35392__7098(csa_tree_add_51_79_groupi_n_10674 ,csa_tree_add_51_79_groupi_n_10572 ,csa_tree_add_51_79_groupi_n_10428);
  or csa_tree_add_51_79_groupi_g35393__6131(csa_tree_add_51_79_groupi_n_10673 ,csa_tree_add_51_79_groupi_n_10578 ,csa_tree_add_51_79_groupi_n_10593);
  or csa_tree_add_51_79_groupi_g35394__1881(csa_tree_add_51_79_groupi_n_10672 ,csa_tree_add_51_79_groupi_n_10571 ,csa_tree_add_51_79_groupi_n_10429);
  or csa_tree_add_51_79_groupi_g35395__5115(csa_tree_add_51_79_groupi_n_10671 ,csa_tree_add_51_79_groupi_n_10566 ,csa_tree_add_51_79_groupi_n_10469);
  and csa_tree_add_51_79_groupi_g35396__7482(csa_tree_add_51_79_groupi_n_10670 ,csa_tree_add_51_79_groupi_n_10566 ,csa_tree_add_51_79_groupi_n_10469);
  and csa_tree_add_51_79_groupi_g35397__4733(csa_tree_add_51_79_groupi_n_10669 ,csa_tree_add_51_79_groupi_n_10564 ,csa_tree_add_51_79_groupi_n_10374);
  or csa_tree_add_51_79_groupi_g35398__6161(csa_tree_add_51_79_groupi_n_10668 ,csa_tree_add_51_79_groupi_n_10564 ,csa_tree_add_51_79_groupi_n_10374);
  and csa_tree_add_51_79_groupi_g35399__9315(csa_tree_add_51_79_groupi_n_10667 ,csa_tree_add_51_79_groupi_n_10521 ,csa_tree_add_51_79_groupi_n_10563);
  or csa_tree_add_51_79_groupi_g35400__9945(csa_tree_add_51_79_groupi_n_10666 ,csa_tree_add_51_79_groupi_n_10521 ,csa_tree_add_51_79_groupi_n_10563);
  nor csa_tree_add_51_79_groupi_g35401__2883(csa_tree_add_51_79_groupi_n_10665 ,csa_tree_add_51_79_groupi_n_10589 ,csa_tree_add_51_79_groupi_n_10281);
  or csa_tree_add_51_79_groupi_g35402__2346(csa_tree_add_51_79_groupi_n_10664 ,csa_tree_add_51_79_groupi_n_10586 ,csa_tree_add_51_79_groupi_n_10532);
  or csa_tree_add_51_79_groupi_g35403__1666(csa_tree_add_51_79_groupi_n_10663 ,csa_tree_add_51_79_groupi_n_10529 ,csa_tree_add_51_79_groupi_n_10549);
  or csa_tree_add_51_79_groupi_g35404__7410(csa_tree_add_51_79_groupi_n_10662 ,csa_tree_add_51_79_groupi_n_10611 ,csa_tree_add_51_79_groupi_n_10562);
  or csa_tree_add_51_79_groupi_g35405__6417(csa_tree_add_51_79_groupi_n_10661 ,csa_tree_add_51_79_groupi_n_10557 ,csa_tree_add_51_79_groupi_n_10517);
  and csa_tree_add_51_79_groupi_g35406__5477(csa_tree_add_51_79_groupi_n_10660 ,csa_tree_add_51_79_groupi_n_10557 ,csa_tree_add_51_79_groupi_n_10517);
  and csa_tree_add_51_79_groupi_g35407__2398(csa_tree_add_51_79_groupi_n_10659 ,csa_tree_add_51_79_groupi_n_10611 ,csa_tree_add_51_79_groupi_n_10562);
  and csa_tree_add_51_79_groupi_g35408__5107(csa_tree_add_51_79_groupi_n_10695 ,csa_tree_add_51_79_groupi_n_10595 ,csa_tree_add_51_79_groupi_n_10503);
  and csa_tree_add_51_79_groupi_g35409__6260(csa_tree_add_51_79_groupi_n_10694 ,csa_tree_add_51_79_groupi_n_10581 ,csa_tree_add_51_79_groupi_n_10499);
  and csa_tree_add_51_79_groupi_g35410__4319(csa_tree_add_51_79_groupi_n_10693 ,csa_tree_add_51_79_groupi_n_10497 ,csa_tree_add_51_79_groupi_n_10590);
  and csa_tree_add_51_79_groupi_g35411__8428(csa_tree_add_51_79_groupi_n_10692 ,csa_tree_add_51_79_groupi_n_10455 ,csa_tree_add_51_79_groupi_n_10551);
  and csa_tree_add_51_79_groupi_g35412__5526(csa_tree_add_51_79_groupi_n_10691 ,csa_tree_add_51_79_groupi_n_10494 ,csa_tree_add_51_79_groupi_n_10588);
  and csa_tree_add_51_79_groupi_g35413__6783(csa_tree_add_51_79_groupi_n_10690 ,csa_tree_add_51_79_groupi_n_10580 ,csa_tree_add_51_79_groupi_n_10505);
  and csa_tree_add_51_79_groupi_g35414__3680(csa_tree_add_51_79_groupi_n_10689 ,csa_tree_add_51_79_groupi_n_10594 ,csa_tree_add_51_79_groupi_n_10501);
  and csa_tree_add_51_79_groupi_g35415__1617(csa_tree_add_51_79_groupi_n_10687 ,csa_tree_add_51_79_groupi_n_10492 ,csa_tree_add_51_79_groupi_n_10585);
  and csa_tree_add_51_79_groupi_g35416__2802(csa_tree_add_51_79_groupi_n_10685 ,csa_tree_add_51_79_groupi_n_10283 ,csa_tree_add_51_79_groupi_n_10582);
  and csa_tree_add_51_79_groupi_g35417__1705(csa_tree_add_51_79_groupi_n_10683 ,csa_tree_add_51_79_groupi_n_10511 ,csa_tree_add_51_79_groupi_n_10603);
  not csa_tree_add_51_79_groupi_g35418(csa_tree_add_51_79_groupi_n_10657 ,csa_tree_add_51_79_groupi_n_10656);
  not csa_tree_add_51_79_groupi_g35419(csa_tree_add_51_79_groupi_n_10654 ,csa_tree_add_51_79_groupi_n_10653);
  not csa_tree_add_51_79_groupi_g35420(csa_tree_add_51_79_groupi_n_10652 ,csa_tree_add_51_79_groupi_n_10651);
  not csa_tree_add_51_79_groupi_g35421(csa_tree_add_51_79_groupi_n_10650 ,csa_tree_add_51_79_groupi_n_10649);
  not csa_tree_add_51_79_groupi_g35422(csa_tree_add_51_79_groupi_n_10646 ,csa_tree_add_51_79_groupi_n_10647);
  not csa_tree_add_51_79_groupi_g35423(csa_tree_add_51_79_groupi_n_10644 ,csa_tree_add_51_79_groupi_n_10643);
  not csa_tree_add_51_79_groupi_g35424(csa_tree_add_51_79_groupi_n_10642 ,csa_tree_add_51_79_groupi_n_10641);
  not csa_tree_add_51_79_groupi_g35425(csa_tree_add_51_79_groupi_n_10639 ,csa_tree_add_51_79_groupi_n_10640);
  nor csa_tree_add_51_79_groupi_g35426__5122(csa_tree_add_51_79_groupi_n_10637 ,csa_tree_add_51_79_groupi_n_10559 ,csa_tree_add_51_79_groupi_n_10568);
  or csa_tree_add_51_79_groupi_g35427__8246(csa_tree_add_51_79_groupi_n_10636 ,csa_tree_add_51_79_groupi_n_10573 ,csa_tree_add_51_79_groupi_n_10325);
  nor csa_tree_add_51_79_groupi_g35428__7098(csa_tree_add_51_79_groupi_n_10635 ,csa_tree_add_51_79_groupi_n_10574 ,csa_tree_add_51_79_groupi_n_10326);
  or csa_tree_add_51_79_groupi_g35429__6131(csa_tree_add_51_79_groupi_n_10634 ,csa_tree_add_51_79_groupi_n_10528 ,csa_tree_add_51_79_groupi_n_10548);
  nor csa_tree_add_51_79_groupi_g35430__1881(csa_tree_add_51_79_groupi_n_10633 ,csa_tree_add_51_79_groupi_n_10389 ,csa_tree_add_51_79_groupi_n_10545);
  or csa_tree_add_51_79_groupi_g35431__5115(csa_tree_add_51_79_groupi_n_10632 ,csa_tree_add_51_79_groupi_n_10569 ,csa_tree_add_51_79_groupi_n_10419);
  nor csa_tree_add_51_79_groupi_g35432__7482(csa_tree_add_51_79_groupi_n_10631 ,csa_tree_add_51_79_groupi_n_10570 ,csa_tree_add_51_79_groupi_n_10420);
  or csa_tree_add_51_79_groupi_g35433__4733(csa_tree_add_51_79_groupi_n_10630 ,csa_tree_add_51_79_groupi_n_10558 ,csa_tree_add_51_79_groupi_n_10567);
  xnor csa_tree_add_51_79_groupi_g35434__6161(csa_tree_add_51_79_groupi_n_10629 ,csa_tree_add_51_79_groupi_n_10422 ,csa_tree_add_51_79_groupi_n_10516);
  xnor csa_tree_add_51_79_groupi_g35435__9315(csa_tree_add_51_79_groupi_n_10628 ,csa_tree_add_51_79_groupi_n_10526 ,csa_tree_add_51_79_groupi_n_10373);
  xnor csa_tree_add_51_79_groupi_g35436__9945(csa_tree_add_51_79_groupi_n_10627 ,csa_tree_add_51_79_groupi_n_10463 ,csa_tree_add_51_79_groupi_n_10531);
  xnor csa_tree_add_51_79_groupi_g35437__2883(csa_tree_add_51_79_groupi_n_10626 ,csa_tree_add_51_79_groupi_n_10489 ,csa_tree_add_51_79_groupi_n_10326);
  xnor csa_tree_add_51_79_groupi_g35438__2346(csa_tree_add_51_79_groupi_n_10625 ,csa_tree_add_51_79_groupi_n_10530 ,csa_tree_add_51_79_groupi_n_10472);
  xnor csa_tree_add_51_79_groupi_g35439__1666(csa_tree_add_51_79_groupi_n_10624 ,csa_tree_add_51_79_groupi_n_10532 ,csa_tree_add_51_79_groupi_n_10371);
  xnor csa_tree_add_51_79_groupi_g35440__7410(csa_tree_add_51_79_groupi_n_10623 ,csa_tree_add_51_79_groupi_n_10529 ,csa_tree_add_51_79_groupi_n_10475);
  xnor csa_tree_add_51_79_groupi_g35441__6417(csa_tree_add_51_79_groupi_n_10622 ,csa_tree_add_51_79_groupi_n_10482 ,csa_tree_add_51_79_groupi_n_10525);
  xnor csa_tree_add_51_79_groupi_g35443__5477(csa_tree_add_51_79_groupi_n_10621 ,csa_tree_add_51_79_groupi_n_10527 ,csa_tree_add_51_79_groupi_n_10369);
  xnor csa_tree_add_51_79_groupi_g35444__2398(csa_tree_add_51_79_groupi_n_10620 ,csa_tree_add_51_79_groupi_n_10524 ,csa_tree_add_51_79_groupi_n_10461);
  xnor csa_tree_add_51_79_groupi_g35445__5107(csa_tree_add_51_79_groupi_n_10619 ,csa_tree_add_51_79_groupi_n_10518 ,csa_tree_add_51_79_groupi_n_10522);
  xnor csa_tree_add_51_79_groupi_g35446__6260(csa_tree_add_51_79_groupi_n_10618 ,csa_tree_add_51_79_groupi_n_10337 ,csa_tree_add_51_79_groupi_n_10520);
  xnor csa_tree_add_51_79_groupi_g35447__4319(csa_tree_add_51_79_groupi_n_10658 ,csa_tree_add_51_79_groupi_n_10424 ,csa_tree_add_51_79_groupi_n_10440);
  xnor csa_tree_add_51_79_groupi_g35448__8428(csa_tree_add_51_79_groupi_n_10656 ,csa_tree_add_51_79_groupi_n_10264 ,csa_tree_add_51_79_groupi_n_10443);
  xnor csa_tree_add_51_79_groupi_g35449__5526(csa_tree_add_51_79_groupi_n_10655 ,csa_tree_add_51_79_groupi_n_10280 ,csa_tree_add_51_79_groupi_n_10447);
  xnor csa_tree_add_51_79_groupi_g35450__6783(csa_tree_add_51_79_groupi_n_10653 ,csa_tree_add_51_79_groupi_n_10154 ,csa_tree_add_51_79_groupi_n_10442);
  xnor csa_tree_add_51_79_groupi_g35451__3680(csa_tree_add_51_79_groupi_n_10651 ,csa_tree_add_51_79_groupi_n_10486 ,csa_tree_add_51_79_groupi_n_10349);
  xnor csa_tree_add_51_79_groupi_g35452__1617(csa_tree_add_51_79_groupi_n_10649 ,csa_tree_add_51_79_groupi_n_10381 ,csa_tree_add_51_79_groupi_n_10439);
  xnor csa_tree_add_51_79_groupi_g35453__2802(csa_tree_add_51_79_groupi_n_10648 ,csa_tree_add_51_79_groupi_n_10379 ,csa_tree_add_51_79_groupi_n_10438);
  xnor csa_tree_add_51_79_groupi_g35454__1705(csa_tree_add_51_79_groupi_n_10647 ,csa_tree_add_51_79_groupi_n_10431 ,csa_tree_add_51_79_groupi_n_10444);
  xnor csa_tree_add_51_79_groupi_g35455__5122(csa_tree_add_51_79_groupi_n_10645 ,csa_tree_add_51_79_groupi_n_10276 ,csa_tree_add_51_79_groupi_n_10445);
  xnor csa_tree_add_51_79_groupi_g35456__8246(csa_tree_add_51_79_groupi_n_10643 ,csa_tree_add_51_79_groupi_n_10277 ,csa_tree_add_51_79_groupi_n_10441);
  xnor csa_tree_add_51_79_groupi_g35457__7098(csa_tree_add_51_79_groupi_n_10641 ,csa_tree_add_51_79_groupi_n_10437 ,csa_tree_add_51_79_groupi_n_10446);
  and csa_tree_add_51_79_groupi_g35458__6131(csa_tree_add_51_79_groupi_n_10640 ,csa_tree_add_51_79_groupi_n_10449 ,csa_tree_add_51_79_groupi_n_10579);
  or csa_tree_add_51_79_groupi_g35459__1881(csa_tree_add_51_79_groupi_n_10638 ,csa_tree_add_51_79_groupi_n_10552 ,csa_tree_add_51_79_groupi_n_10451);
  not csa_tree_add_51_79_groupi_g35460(csa_tree_add_51_79_groupi_n_10615 ,csa_tree_add_51_79_groupi_n_10614);
  not csa_tree_add_51_79_groupi_g35461(csa_tree_add_51_79_groupi_n_10608 ,csa_tree_add_51_79_groupi_n_10609);
  nor csa_tree_add_51_79_groupi_g35462__5115(csa_tree_add_51_79_groupi_n_10607 ,csa_tree_add_51_79_groupi_n_10468 ,csa_tree_add_51_79_groupi_n_10472);
  nor csa_tree_add_51_79_groupi_g35463__7482(csa_tree_add_51_79_groupi_n_10606 ,csa_tree_add_51_79_groupi_n_10422 ,csa_tree_add_51_79_groupi_n_10516);
  or csa_tree_add_51_79_groupi_g35464__4733(csa_tree_add_51_79_groupi_n_10605 ,csa_tree_add_51_79_groupi_n_10421 ,csa_tree_add_51_79_groupi_n_10515);
  nor csa_tree_add_51_79_groupi_g35465__6161(csa_tree_add_51_79_groupi_n_10604 ,csa_tree_add_51_79_groupi_n_10375 ,csa_tree_add_51_79_groupi_n_10466);
  or csa_tree_add_51_79_groupi_g35466__9315(csa_tree_add_51_79_groupi_n_10603 ,csa_tree_add_51_79_groupi_n_10278 ,csa_tree_add_51_79_groupi_n_10509);
  or csa_tree_add_51_79_groupi_g35467__9945(csa_tree_add_51_79_groupi_n_10602 ,csa_tree_add_51_79_groupi_n_10376 ,csa_tree_add_51_79_groupi_n_10465);
  and csa_tree_add_51_79_groupi_g35468__2883(csa_tree_add_51_79_groupi_n_10601 ,csa_tree_add_51_79_groupi_n_10520 ,csa_tree_add_51_79_groupi_n_10337);
  or csa_tree_add_51_79_groupi_g35469__2346(csa_tree_add_51_79_groupi_n_10600 ,csa_tree_add_51_79_groupi_n_10520 ,csa_tree_add_51_79_groupi_n_10337);
  or csa_tree_add_51_79_groupi_g35470__1666(csa_tree_add_51_79_groupi_n_10599 ,csa_tree_add_51_79_groupi_n_10458 ,csa_tree_add_51_79_groupi_n_10462);
  nor csa_tree_add_51_79_groupi_g35471__7410(csa_tree_add_51_79_groupi_n_10598 ,csa_tree_add_51_79_groupi_n_10459 ,csa_tree_add_51_79_groupi_n_10463);
  or csa_tree_add_51_79_groupi_g35472__6417(csa_tree_add_51_79_groupi_n_10597 ,csa_tree_add_51_79_groupi_n_10522 ,csa_tree_add_51_79_groupi_n_10518);
  and csa_tree_add_51_79_groupi_g35473__5477(csa_tree_add_51_79_groupi_n_10596 ,csa_tree_add_51_79_groupi_n_10522 ,csa_tree_add_51_79_groupi_n_10518);
  or csa_tree_add_51_79_groupi_g35474__2398(csa_tree_add_51_79_groupi_n_10595 ,csa_tree_add_51_79_groupi_n_10504 ,csa_tree_add_51_79_groupi_n_10390);
  or csa_tree_add_51_79_groupi_g35475__5107(csa_tree_add_51_79_groupi_n_10594 ,csa_tree_add_51_79_groupi_n_10514 ,csa_tree_add_51_79_groupi_n_10082);
  nor csa_tree_add_51_79_groupi_g35476__6260(csa_tree_add_51_79_groupi_n_10593 ,csa_tree_add_51_79_groupi_n_10524 ,csa_tree_add_51_79_groupi_n_10460);
  or csa_tree_add_51_79_groupi_g35477__4319(csa_tree_add_51_79_groupi_n_10592 ,csa_tree_add_51_79_groupi_n_10523 ,csa_tree_add_51_79_groupi_n_10461);
  nor csa_tree_add_51_79_groupi_g35478__8428(csa_tree_add_51_79_groupi_n_10591 ,csa_tree_add_51_79_groupi_n_10457 ,csa_tree_add_51_79_groupi_n_10373);
  or csa_tree_add_51_79_groupi_g35479__5526(csa_tree_add_51_79_groupi_n_10590 ,csa_tree_add_51_79_groupi_n_10432 ,csa_tree_add_51_79_groupi_n_10496);
  and csa_tree_add_51_79_groupi_g35480__6783(csa_tree_add_51_79_groupi_n_10589 ,csa_tree_add_51_79_groupi_n_10481 ,csa_tree_add_51_79_groupi_n_10519);
  or csa_tree_add_51_79_groupi_g35481__3680(csa_tree_add_51_79_groupi_n_10588 ,csa_tree_add_51_79_groupi_n_10493 ,csa_tree_add_51_79_groupi_n_10436);
  or csa_tree_add_51_79_groupi_g35482__1617(csa_tree_add_51_79_groupi_n_10587 ,csa_tree_add_51_79_groupi_n_10371 ,csa_tree_add_51_79_groupi_n_10483);
  and csa_tree_add_51_79_groupi_g35483__2802(csa_tree_add_51_79_groupi_n_10586 ,csa_tree_add_51_79_groupi_n_10371 ,csa_tree_add_51_79_groupi_n_10483);
  or csa_tree_add_51_79_groupi_g35484__1705(csa_tree_add_51_79_groupi_n_10585 ,csa_tree_add_51_79_groupi_n_10491 ,csa_tree_add_51_79_groupi_n_10434);
  or csa_tree_add_51_79_groupi_g35485__5122(csa_tree_add_51_79_groupi_n_10584 ,csa_tree_add_51_79_groupi_n_10456 ,csa_tree_add_51_79_groupi_n_10372);
  nor csa_tree_add_51_79_groupi_g35486__8246(csa_tree_add_51_79_groupi_n_10583 ,csa_tree_add_51_79_groupi_n_10481 ,csa_tree_add_51_79_groupi_n_10519);
  or csa_tree_add_51_79_groupi_g35487__7098(csa_tree_add_51_79_groupi_n_10582 ,csa_tree_add_51_79_groupi_n_10316 ,csa_tree_add_51_79_groupi_n_10486);
  or csa_tree_add_51_79_groupi_g35488__6131(csa_tree_add_51_79_groupi_n_10581 ,csa_tree_add_51_79_groupi_n_10495 ,csa_tree_add_51_79_groupi_n_10340);
  or csa_tree_add_51_79_groupi_g35489__1881(csa_tree_add_51_79_groupi_n_10580 ,csa_tree_add_51_79_groupi_n_10500 ,csa_tree_add_51_79_groupi_n_10430);
  or csa_tree_add_51_79_groupi_g35490__5115(csa_tree_add_51_79_groupi_n_10579 ,csa_tree_add_51_79_groupi_n_10513 ,csa_tree_add_51_79_groupi_n_10388);
  and csa_tree_add_51_79_groupi_g35491__7482(csa_tree_add_51_79_groupi_n_10617 ,csa_tree_add_51_79_groupi_n_10508 ,csa_tree_add_51_79_groupi_n_10315);
  and csa_tree_add_51_79_groupi_g35492__4733(csa_tree_add_51_79_groupi_n_10616 ,csa_tree_add_51_79_groupi_n_10502 ,csa_tree_add_51_79_groupi_n_10414);
  or csa_tree_add_51_79_groupi_g35493__6161(csa_tree_add_51_79_groupi_n_10614 ,csa_tree_add_51_79_groupi_n_10395 ,csa_tree_add_51_79_groupi_n_10506);
  and csa_tree_add_51_79_groupi_g35494__9315(csa_tree_add_51_79_groupi_n_10613 ,csa_tree_add_51_79_groupi_n_10401 ,csa_tree_add_51_79_groupi_n_10507);
  and csa_tree_add_51_79_groupi_g35495__9945(csa_tree_add_51_79_groupi_n_10612 ,csa_tree_add_51_79_groupi_n_10361 ,csa_tree_add_51_79_groupi_n_10512);
  and csa_tree_add_51_79_groupi_g35496__2883(csa_tree_add_51_79_groupi_n_10611 ,csa_tree_add_51_79_groupi_n_10410 ,csa_tree_add_51_79_groupi_n_10490);
  and csa_tree_add_51_79_groupi_g35497__2346(csa_tree_add_51_79_groupi_n_10610 ,csa_tree_add_51_79_groupi_n_10510 ,csa_tree_add_51_79_groupi_n_10417);
  and csa_tree_add_51_79_groupi_g35498__1666(csa_tree_add_51_79_groupi_n_10609 ,csa_tree_add_51_79_groupi_n_10498 ,csa_tree_add_51_79_groupi_n_10402);
  not csa_tree_add_51_79_groupi_g35499(csa_tree_add_51_79_groupi_n_10578 ,csa_tree_add_51_79_groupi_n_10577);
  not csa_tree_add_51_79_groupi_g35500(csa_tree_add_51_79_groupi_n_10574 ,csa_tree_add_51_79_groupi_n_10573);
  not csa_tree_add_51_79_groupi_g35501(csa_tree_add_51_79_groupi_n_10572 ,csa_tree_add_51_79_groupi_n_10571);
  not csa_tree_add_51_79_groupi_g35502(csa_tree_add_51_79_groupi_n_10570 ,csa_tree_add_51_79_groupi_n_10569);
  not csa_tree_add_51_79_groupi_g35503(csa_tree_add_51_79_groupi_n_10568 ,csa_tree_add_51_79_groupi_n_10567);
  not csa_tree_add_51_79_groupi_g35504(csa_tree_add_51_79_groupi_n_10561 ,csa_tree_add_51_79_groupi_n_10560);
  not csa_tree_add_51_79_groupi_g35505(csa_tree_add_51_79_groupi_n_10558 ,csa_tree_add_51_79_groupi_n_10559);
  not csa_tree_add_51_79_groupi_g35506(csa_tree_add_51_79_groupi_n_10556 ,csa_tree_add_51_79_groupi_n_10555);
  or csa_tree_add_51_79_groupi_g35507__7410(csa_tree_add_51_79_groupi_n_10554 ,csa_tree_add_51_79_groupi_n_10467 ,csa_tree_add_51_79_groupi_n_10471);
  and csa_tree_add_51_79_groupi_g35508__6417(csa_tree_add_51_79_groupi_n_10553 ,csa_tree_add_51_79_groupi_n_10470 ,csa_tree_add_51_79_groupi_n_10367);
  nor csa_tree_add_51_79_groupi_g35509__5477(csa_tree_add_51_79_groupi_n_10552 ,csa_tree_add_51_79_groupi_n_10273 ,csa_tree_add_51_79_groupi_n_10452);
  or csa_tree_add_51_79_groupi_g35510__2398(csa_tree_add_51_79_groupi_n_10551 ,csa_tree_add_51_79_groupi_n_10218 ,csa_tree_add_51_79_groupi_n_10453);
  or csa_tree_add_51_79_groupi_g35511__5107(csa_tree_add_51_79_groupi_n_10550 ,csa_tree_add_51_79_groupi_n_10474 ,csa_tree_add_51_79_groupi_n_10476);
  nor csa_tree_add_51_79_groupi_g35512__6260(csa_tree_add_51_79_groupi_n_10549 ,csa_tree_add_51_79_groupi_n_10475 ,csa_tree_add_51_79_groupi_n_10477);
  nor csa_tree_add_51_79_groupi_g35513__4319(csa_tree_add_51_79_groupi_n_10548 ,csa_tree_add_51_79_groupi_n_10479 ,csa_tree_add_51_79_groupi_n_10369);
  or csa_tree_add_51_79_groupi_g35514__8428(csa_tree_add_51_79_groupi_n_10547 ,csa_tree_add_51_79_groupi_n_10478 ,csa_tree_add_51_79_groupi_n_10368);
  nor csa_tree_add_51_79_groupi_g35515__5526(csa_tree_add_51_79_groupi_n_10546 ,csa_tree_add_51_79_groupi_n_10480 ,csa_tree_add_51_79_groupi_n_10386);
  and csa_tree_add_51_79_groupi_g35516__6783(csa_tree_add_51_79_groupi_n_10545 ,csa_tree_add_51_79_groupi_n_10480 ,csa_tree_add_51_79_groupi_n_10386);
  or csa_tree_add_51_79_groupi_g35517__3680(csa_tree_add_51_79_groupi_n_10544 ,csa_tree_add_51_79_groupi_n_10470 ,csa_tree_add_51_79_groupi_n_10367);
  xnor csa_tree_add_51_79_groupi_g35518__1617(csa_tree_add_51_79_groupi_n_10543 ,csa_tree_add_51_79_groupi_n_10263 ,csa_tree_add_51_79_groupi_n_10430);
  xnor csa_tree_add_51_79_groupi_g35519__2802(csa_tree_add_51_79_groupi_n_10542 ,csa_tree_add_51_79_groupi_n_10135 ,csa_tree_add_51_79_groupi_n_10434);
  xnor csa_tree_add_51_79_groupi_g35520__1705(csa_tree_add_51_79_groupi_n_10541 ,csa_tree_add_51_79_groupi_n_10129 ,csa_tree_add_51_79_groupi_n_10383);
  xnor csa_tree_add_51_79_groupi_g35521__5122(csa_tree_add_51_79_groupi_n_10540 ,csa_tree_add_51_79_groupi_n_10367 ,csa_tree_add_51_79_groupi_n_10435);
  xnor csa_tree_add_51_79_groupi_g35522__8246(csa_tree_add_51_79_groupi_n_10539 ,csa_tree_add_51_79_groupi_n_10423 ,csa_tree_add_51_79_groupi_n_10266);
  xnor csa_tree_add_51_79_groupi_g35523__7098(csa_tree_add_51_79_groupi_n_10538 ,csa_tree_add_51_79_groupi_n_10386 ,csa_tree_add_51_79_groupi_n_10389);
  xnor csa_tree_add_51_79_groupi_g35524__6131(csa_tree_add_51_79_groupi_n_10537 ,csa_tree_add_51_79_groupi_n_10384 ,csa_tree_add_51_79_groupi_n_10427);
  xnor csa_tree_add_51_79_groupi_g35525__1881(csa_tree_add_51_79_groupi_n_10536 ,csa_tree_add_51_79_groupi_n_10139 ,csa_tree_add_51_79_groupi_n_10390);
  xnor csa_tree_add_51_79_groupi_g35526__5115(csa_tree_add_51_79_groupi_n_10535 ,csa_tree_add_51_79_groupi_n_10374 ,csa_tree_add_51_79_groupi_n_10433);
  xnor csa_tree_add_51_79_groupi_g35527__7482(csa_tree_add_51_79_groupi_n_10534 ,csa_tree_add_51_79_groupi_n_10376 ,csa_tree_add_51_79_groupi_n_10342);
  xnor csa_tree_add_51_79_groupi_g35528__4733(csa_tree_add_51_79_groupi_n_10533 ,csa_tree_add_51_79_groupi_n_10329 ,csa_tree_add_51_79_groupi_n_10378);
  xnor csa_tree_add_51_79_groupi_g35529__6161(csa_tree_add_51_79_groupi_n_10577 ,csa_tree_add_51_79_groupi_n_10282 ,csa_tree_add_51_79_groupi_n_10352);
  xnor csa_tree_add_51_79_groupi_g35530__9315(csa_tree_add_51_79_groupi_n_10576 ,csa_tree_add_51_79_groupi_n_10370 ,csa_tree_add_51_79_groupi_n_10354);
  xnor csa_tree_add_51_79_groupi_g35531__9945(csa_tree_add_51_79_groupi_n_10575 ,csa_tree_add_51_79_groupi_n_10220 ,csa_tree_add_51_79_groupi_n_10356);
  xnor csa_tree_add_51_79_groupi_g35532__2883(csa_tree_add_51_79_groupi_n_10573 ,csa_tree_add_51_79_groupi_n_10391 ,csa_tree_add_51_79_groupi_n_10235);
  xnor csa_tree_add_51_79_groupi_g35533__2346(csa_tree_add_51_79_groupi_n_10571 ,csa_tree_add_51_79_groupi_n_9869 ,csa_tree_add_51_79_groupi_n_10347);
  xnor csa_tree_add_51_79_groupi_g35534__1666(csa_tree_add_51_79_groupi_n_10569 ,csa_tree_add_51_79_groupi_n_10152 ,csa_tree_add_51_79_groupi_n_10346);
  xnor csa_tree_add_51_79_groupi_g35535__7410(csa_tree_add_51_79_groupi_n_10567 ,csa_tree_add_51_79_groupi_n_10392 ,csa_tree_add_51_79_groupi_n_10355);
  xnor csa_tree_add_51_79_groupi_g35536__6417(csa_tree_add_51_79_groupi_n_10566 ,csa_tree_add_51_79_groupi_n_10145 ,csa_tree_add_51_79_groupi_n_10351);
  xnor csa_tree_add_51_79_groupi_g35537__5477(csa_tree_add_51_79_groupi_n_10565 ,csa_tree_add_51_79_groupi_n_10339 ,csa_tree_add_51_79_groupi_n_10348);
  xnor csa_tree_add_51_79_groupi_g35538__2398(csa_tree_add_51_79_groupi_n_10564 ,csa_tree_add_51_79_groupi_n_10077 ,csa_tree_add_51_79_groupi_n_10350);
  xnor csa_tree_add_51_79_groupi_g35539__5107(csa_tree_add_51_79_groupi_n_10563 ,csa_tree_add_51_79_groupi_n_10010 ,csa_tree_add_51_79_groupi_n_10353);
  xnor csa_tree_add_51_79_groupi_g35540__6260(csa_tree_add_51_79_groupi_n_10562 ,csa_tree_add_51_79_groupi_n_10155 ,csa_tree_add_51_79_groupi_n_10357);
  xnor csa_tree_add_51_79_groupi_g35541__4319(csa_tree_add_51_79_groupi_n_10560 ,csa_tree_add_51_79_groupi_n_10270 ,csa_tree_add_51_79_groupi_n_10343);
  or csa_tree_add_51_79_groupi_g35542__8428(csa_tree_add_51_79_groupi_n_10559 ,csa_tree_add_51_79_groupi_n_10454 ,csa_tree_add_51_79_groupi_n_10122);
  xnor csa_tree_add_51_79_groupi_g35543__5526(csa_tree_add_51_79_groupi_n_10557 ,csa_tree_add_51_79_groupi_n_10223 ,csa_tree_add_51_79_groupi_n_10344);
  xnor csa_tree_add_51_79_groupi_g35544__6783(csa_tree_add_51_79_groupi_n_10555 ,csa_tree_add_51_79_groupi_n_10274 ,csa_tree_add_51_79_groupi_n_10345);
  not csa_tree_add_51_79_groupi_g35545(csa_tree_add_51_79_groupi_n_10528 ,csa_tree_add_51_79_groupi_n_10527);
  not csa_tree_add_51_79_groupi_g35546(csa_tree_add_51_79_groupi_n_10524 ,csa_tree_add_51_79_groupi_n_10523);
  not csa_tree_add_51_79_groupi_g35548(csa_tree_add_51_79_groupi_n_10515 ,csa_tree_add_51_79_groupi_n_10516);
  and csa_tree_add_51_79_groupi_g35549__3680(csa_tree_add_51_79_groupi_n_10514 ,csa_tree_add_51_79_groupi_n_10370 ,csa_tree_add_51_79_groupi_n_10131);
  nor csa_tree_add_51_79_groupi_g35550__1617(csa_tree_add_51_79_groupi_n_10513 ,csa_tree_add_51_79_groupi_n_10328 ,csa_tree_add_51_79_groupi_n_10378);
  or csa_tree_add_51_79_groupi_g35551__2802(csa_tree_add_51_79_groupi_n_10512 ,csa_tree_add_51_79_groupi_n_10360 ,csa_tree_add_51_79_groupi_n_10222);
  or csa_tree_add_51_79_groupi_g35552__1705(csa_tree_add_51_79_groupi_n_10511 ,csa_tree_add_51_79_groupi_n_10424 ,csa_tree_add_51_79_groupi_n_10335);
  or csa_tree_add_51_79_groupi_g35553__5122(csa_tree_add_51_79_groupi_n_10510 ,csa_tree_add_51_79_groupi_n_10404 ,csa_tree_add_51_79_groupi_n_10437);
  and csa_tree_add_51_79_groupi_g35554__8246(csa_tree_add_51_79_groupi_n_10509 ,csa_tree_add_51_79_groupi_n_10424 ,csa_tree_add_51_79_groupi_n_10335);
  or csa_tree_add_51_79_groupi_g35555__7098(csa_tree_add_51_79_groupi_n_10508 ,csa_tree_add_51_79_groupi_n_10392 ,csa_tree_add_51_79_groupi_n_10314);
  or csa_tree_add_51_79_groupi_g35556__6131(csa_tree_add_51_79_groupi_n_10507 ,csa_tree_add_51_79_groupi_n_10276 ,csa_tree_add_51_79_groupi_n_10400);
  nor csa_tree_add_51_79_groupi_g35557__1881(csa_tree_add_51_79_groupi_n_10506 ,csa_tree_add_51_79_groupi_n_10394 ,csa_tree_add_51_79_groupi_n_10280);
  or csa_tree_add_51_79_groupi_g35558__5115(csa_tree_add_51_79_groupi_n_10505 ,csa_tree_add_51_79_groupi_n_10262 ,csa_tree_add_51_79_groupi_n_10366);
  nor csa_tree_add_51_79_groupi_g35559__7482(csa_tree_add_51_79_groupi_n_10504 ,csa_tree_add_51_79_groupi_n_10425 ,csa_tree_add_51_79_groupi_n_10139);
  or csa_tree_add_51_79_groupi_g35560__4733(csa_tree_add_51_79_groupi_n_10503 ,csa_tree_add_51_79_groupi_n_10426 ,csa_tree_add_51_79_groupi_n_10138);
  or csa_tree_add_51_79_groupi_g35561__6161(csa_tree_add_51_79_groupi_n_10502 ,csa_tree_add_51_79_groupi_n_10415 ,csa_tree_add_51_79_groupi_n_10277);
  or csa_tree_add_51_79_groupi_g35562__9315(csa_tree_add_51_79_groupi_n_10501 ,csa_tree_add_51_79_groupi_n_10370 ,csa_tree_add_51_79_groupi_n_10131);
  nor csa_tree_add_51_79_groupi_g35563__9945(csa_tree_add_51_79_groupi_n_10500 ,csa_tree_add_51_79_groupi_n_10263 ,csa_tree_add_51_79_groupi_n_10365);
  or csa_tree_add_51_79_groupi_g35564__2883(csa_tree_add_51_79_groupi_n_10499 ,csa_tree_add_51_79_groupi_n_10129 ,csa_tree_add_51_79_groupi_n_10382);
  or csa_tree_add_51_79_groupi_g35565__2346(csa_tree_add_51_79_groupi_n_10498 ,csa_tree_add_51_79_groupi_n_10431 ,csa_tree_add_51_79_groupi_n_10399);
  or csa_tree_add_51_79_groupi_g35566__1666(csa_tree_add_51_79_groupi_n_10497 ,csa_tree_add_51_79_groupi_n_10266 ,csa_tree_add_51_79_groupi_n_10423);
  and csa_tree_add_51_79_groupi_g35567__7410(csa_tree_add_51_79_groupi_n_10496 ,csa_tree_add_51_79_groupi_n_10266 ,csa_tree_add_51_79_groupi_n_10423);
  nor csa_tree_add_51_79_groupi_g35568__6417(csa_tree_add_51_79_groupi_n_10495 ,csa_tree_add_51_79_groupi_n_10128 ,csa_tree_add_51_79_groupi_n_10383);
  or csa_tree_add_51_79_groupi_g35569__5477(csa_tree_add_51_79_groupi_n_10494 ,csa_tree_add_51_79_groupi_n_10427 ,csa_tree_add_51_79_groupi_n_10384);
  and csa_tree_add_51_79_groupi_g35570__2398(csa_tree_add_51_79_groupi_n_10493 ,csa_tree_add_51_79_groupi_n_10427 ,csa_tree_add_51_79_groupi_n_10384);
  or csa_tree_add_51_79_groupi_g35571__5107(csa_tree_add_51_79_groupi_n_10492 ,csa_tree_add_51_79_groupi_n_10385 ,csa_tree_add_51_79_groupi_n_10135);
  and csa_tree_add_51_79_groupi_g35572__6260(csa_tree_add_51_79_groupi_n_10491 ,csa_tree_add_51_79_groupi_n_10385 ,csa_tree_add_51_79_groupi_n_10135);
  or csa_tree_add_51_79_groupi_g35573__4319(csa_tree_add_51_79_groupi_n_10490 ,csa_tree_add_51_79_groupi_n_10413 ,csa_tree_add_51_79_groupi_n_10341);
  and csa_tree_add_51_79_groupi_g35574__8428(csa_tree_add_51_79_groupi_n_10532 ,csa_tree_add_51_79_groupi_n_10213 ,csa_tree_add_51_79_groupi_n_10396);
  and csa_tree_add_51_79_groupi_g35575__5526(csa_tree_add_51_79_groupi_n_10531 ,csa_tree_add_51_79_groupi_n_10416 ,csa_tree_add_51_79_groupi_n_10292);
  and csa_tree_add_51_79_groupi_g35576__6783(csa_tree_add_51_79_groupi_n_10530 ,csa_tree_add_51_79_groupi_n_10290 ,csa_tree_add_51_79_groupi_n_10411);
  and csa_tree_add_51_79_groupi_g35577__3680(csa_tree_add_51_79_groupi_n_10529 ,csa_tree_add_51_79_groupi_n_10260 ,csa_tree_add_51_79_groupi_n_10405);
  or csa_tree_add_51_79_groupi_g35578__1617(csa_tree_add_51_79_groupi_n_10527 ,csa_tree_add_51_79_groupi_n_10409 ,csa_tree_add_51_79_groupi_n_10310);
  and csa_tree_add_51_79_groupi_g35579__2802(csa_tree_add_51_79_groupi_n_10526 ,csa_tree_add_51_79_groupi_n_10397 ,csa_tree_add_51_79_groupi_n_10284);
  and csa_tree_add_51_79_groupi_g35580__1705(csa_tree_add_51_79_groupi_n_10525 ,csa_tree_add_51_79_groupi_n_10407 ,csa_tree_add_51_79_groupi_n_10307);
  and csa_tree_add_51_79_groupi_g35581__5122(csa_tree_add_51_79_groupi_n_10523 ,csa_tree_add_51_79_groupi_n_10418 ,csa_tree_add_51_79_groupi_n_10302);
  and csa_tree_add_51_79_groupi_g35582__8246(csa_tree_add_51_79_groupi_n_10522 ,csa_tree_add_51_79_groupi_n_10406 ,csa_tree_add_51_79_groupi_n_10305);
  and csa_tree_add_51_79_groupi_g35583__7098(csa_tree_add_51_79_groupi_n_10521 ,csa_tree_add_51_79_groupi_n_10258 ,csa_tree_add_51_79_groupi_n_10403);
  and csa_tree_add_51_79_groupi_g35584__6131(csa_tree_add_51_79_groupi_n_10520 ,csa_tree_add_51_79_groupi_n_10287 ,csa_tree_add_51_79_groupi_n_10398);
  and csa_tree_add_51_79_groupi_g35585__1881(csa_tree_add_51_79_groupi_n_10519 ,csa_tree_add_51_79_groupi_n_10358 ,csa_tree_add_51_79_groupi_n_10252);
  and csa_tree_add_51_79_groupi_g35586__5115(csa_tree_add_51_79_groupi_n_10518 ,csa_tree_add_51_79_groupi_n_10297 ,csa_tree_add_51_79_groupi_n_10393);
  and csa_tree_add_51_79_groupi_g35587__7482(csa_tree_add_51_79_groupi_n_10517 ,csa_tree_add_51_79_groupi_n_10201 ,csa_tree_add_51_79_groupi_n_10408);
  or csa_tree_add_51_79_groupi_g35588__4733(csa_tree_add_51_79_groupi_n_10516 ,csa_tree_add_51_79_groupi_n_10318 ,csa_tree_add_51_79_groupi_n_10412);
  not csa_tree_add_51_79_groupi_g35589(csa_tree_add_51_79_groupi_n_10488 ,csa_tree_add_51_79_groupi_n_10487);
  not csa_tree_add_51_79_groupi_g35590(csa_tree_add_51_79_groupi_n_10479 ,csa_tree_add_51_79_groupi_n_10478);
  not csa_tree_add_51_79_groupi_g35591(csa_tree_add_51_79_groupi_n_10477 ,csa_tree_add_51_79_groupi_n_10476);
  not csa_tree_add_51_79_groupi_g35592(csa_tree_add_51_79_groupi_n_10475 ,csa_tree_add_51_79_groupi_n_10474);
  not csa_tree_add_51_79_groupi_g35593(csa_tree_add_51_79_groupi_n_10472 ,csa_tree_add_51_79_groupi_n_10471);
  not csa_tree_add_51_79_groupi_g35594(csa_tree_add_51_79_groupi_n_10468 ,csa_tree_add_51_79_groupi_n_10467);
  not csa_tree_add_51_79_groupi_g35595(csa_tree_add_51_79_groupi_n_10466 ,csa_tree_add_51_79_groupi_n_10465);
  not csa_tree_add_51_79_groupi_g35596(csa_tree_add_51_79_groupi_n_10463 ,csa_tree_add_51_79_groupi_n_10462);
  not csa_tree_add_51_79_groupi_g35597(csa_tree_add_51_79_groupi_n_10460 ,csa_tree_add_51_79_groupi_n_10461);
  not csa_tree_add_51_79_groupi_g35598(csa_tree_add_51_79_groupi_n_10459 ,csa_tree_add_51_79_groupi_n_10458);
  not csa_tree_add_51_79_groupi_g35599(csa_tree_add_51_79_groupi_n_10457 ,csa_tree_add_51_79_groupi_n_10456);
  or csa_tree_add_51_79_groupi_g35600__6161(csa_tree_add_51_79_groupi_n_10455 ,csa_tree_add_51_79_groupi_n_10380 ,csa_tree_add_51_79_groupi_n_10323);
  and csa_tree_add_51_79_groupi_g35601__9315(csa_tree_add_51_79_groupi_n_10454 ,csa_tree_add_51_79_groupi_n_10391 ,csa_tree_add_51_79_groupi_n_10124);
  nor csa_tree_add_51_79_groupi_g35602__9945(csa_tree_add_51_79_groupi_n_10453 ,csa_tree_add_51_79_groupi_n_10381 ,csa_tree_add_51_79_groupi_n_10324);
  and csa_tree_add_51_79_groupi_g35603__2883(csa_tree_add_51_79_groupi_n_10452 ,csa_tree_add_51_79_groupi_n_10160 ,csa_tree_add_51_79_groupi_n_10379);
  nor csa_tree_add_51_79_groupi_g35604__2346(csa_tree_add_51_79_groupi_n_10451 ,csa_tree_add_51_79_groupi_n_10160 ,csa_tree_add_51_79_groupi_n_10379);
  xnor csa_tree_add_51_79_groupi_g35605__1666(out1[2] ,csa_tree_add_51_79_groupi_n_9793 ,csa_tree_add_51_79_groupi_n_10244);
  or csa_tree_add_51_79_groupi_g35606__7410(csa_tree_add_51_79_groupi_n_10449 ,csa_tree_add_51_79_groupi_n_10329 ,csa_tree_add_51_79_groupi_n_10377);
  xnor csa_tree_add_51_79_groupi_g35607__6417(csa_tree_add_51_79_groupi_n_10448 ,csa_tree_add_51_79_groupi_n_10336 ,csa_tree_add_51_79_groupi_n_9999);
  xnor csa_tree_add_51_79_groupi_g35608__5477(csa_tree_add_51_79_groupi_n_10447 ,csa_tree_add_51_79_groupi_n_10267 ,csa_tree_add_51_79_groupi_n_10332);
  xnor csa_tree_add_51_79_groupi_g35609__2398(csa_tree_add_51_79_groupi_n_10446 ,csa_tree_add_51_79_groupi_n_10271 ,csa_tree_add_51_79_groupi_n_10327);
  xnor csa_tree_add_51_79_groupi_g35610__5107(csa_tree_add_51_79_groupi_n_10445 ,csa_tree_add_51_79_groupi_n_10140 ,csa_tree_add_51_79_groupi_n_10333);
  xnor csa_tree_add_51_79_groupi_g35611__6260(csa_tree_add_51_79_groupi_n_10444 ,csa_tree_add_51_79_groupi_n_10272 ,csa_tree_add_51_79_groupi_n_10334);
  xnor csa_tree_add_51_79_groupi_g35612__4319(csa_tree_add_51_79_groupi_n_10443 ,csa_tree_add_51_79_groupi_n_10265 ,csa_tree_add_51_79_groupi_n_10341);
  xnor csa_tree_add_51_79_groupi_g35613__8428(csa_tree_add_51_79_groupi_n_10442 ,csa_tree_add_51_79_groupi_n_10158 ,csa_tree_add_51_79_groupi_n_10338);
  xnor csa_tree_add_51_79_groupi_g35614__5526(csa_tree_add_51_79_groupi_n_10441 ,csa_tree_add_51_79_groupi_n_10214 ,csa_tree_add_51_79_groupi_n_10322);
  xnor csa_tree_add_51_79_groupi_g35615__6783(csa_tree_add_51_79_groupi_n_10440 ,csa_tree_add_51_79_groupi_n_10335 ,csa_tree_add_51_79_groupi_n_10278);
  xnor csa_tree_add_51_79_groupi_g35616__3680(csa_tree_add_51_79_groupi_n_10439 ,csa_tree_add_51_79_groupi_n_10218 ,csa_tree_add_51_79_groupi_n_10324);
  xnor csa_tree_add_51_79_groupi_g35617__1617(csa_tree_add_51_79_groupi_n_10438 ,csa_tree_add_51_79_groupi_n_10159 ,csa_tree_add_51_79_groupi_n_10273);
  and csa_tree_add_51_79_groupi_g35618__2802(csa_tree_add_51_79_groupi_n_10489 ,csa_tree_add_51_79_groupi_n_10251 ,csa_tree_add_51_79_groupi_n_10359);
  or csa_tree_add_51_79_groupi_g35619__1705(csa_tree_add_51_79_groupi_n_10487 ,csa_tree_add_51_79_groupi_n_10364 ,csa_tree_add_51_79_groupi_n_10261);
  xnor csa_tree_add_51_79_groupi_g35620__5122(csa_tree_add_51_79_groupi_n_10486 ,csa_tree_add_51_79_groupi_n_10081 ,csa_tree_add_51_79_groupi_n_10225);
  xnor csa_tree_add_51_79_groupi_g35621__8246(csa_tree_add_51_79_groupi_n_10485 ,csa_tree_add_51_79_groupi_n_10074 ,csa_tree_add_51_79_groupi_n_10228);
  xnor csa_tree_add_51_79_groupi_g35622__7098(csa_tree_add_51_79_groupi_n_10484 ,csa_tree_add_51_79_groupi_n_10072 ,csa_tree_add_51_79_groupi_n_10227);
  xnor csa_tree_add_51_79_groupi_g35623__6131(csa_tree_add_51_79_groupi_n_10483 ,csa_tree_add_51_79_groupi_n_10024 ,csa_tree_add_51_79_groupi_n_10239);
  xnor csa_tree_add_51_79_groupi_g35624__1881(csa_tree_add_51_79_groupi_n_10482 ,csa_tree_add_51_79_groupi_n_10219 ,csa_tree_add_51_79_groupi_n_10231);
  xnor csa_tree_add_51_79_groupi_g35625__5115(csa_tree_add_51_79_groupi_n_10481 ,csa_tree_add_51_79_groupi_n_10083 ,csa_tree_add_51_79_groupi_n_10226);
  xnor csa_tree_add_51_79_groupi_g35626__7482(csa_tree_add_51_79_groupi_n_10480 ,csa_tree_add_51_79_groupi_n_9987 ,csa_tree_add_51_79_groupi_n_10232);
  xnor csa_tree_add_51_79_groupi_g35627__4733(csa_tree_add_51_79_groupi_n_10478 ,csa_tree_add_51_79_groupi_n_10089 ,csa_tree_add_51_79_groupi_n_10233);
  xnor csa_tree_add_51_79_groupi_g35628__6161(csa_tree_add_51_79_groupi_n_10476 ,csa_tree_add_51_79_groupi_n_10279 ,csa_tree_add_51_79_groupi_n_10245);
  xnor csa_tree_add_51_79_groupi_g35629__9315(csa_tree_add_51_79_groupi_n_10474 ,csa_tree_add_51_79_groupi_n_10091 ,csa_tree_add_51_79_groupi_n_10230);
  xnor csa_tree_add_51_79_groupi_g35630__9945(csa_tree_add_51_79_groupi_n_10473 ,csa_tree_add_51_79_groupi_n_10148 ,csa_tree_add_51_79_groupi_n_10236);
  xnor csa_tree_add_51_79_groupi_g35631__2883(csa_tree_add_51_79_groupi_n_10471 ,csa_tree_add_51_79_groupi_n_10134 ,csa_tree_add_51_79_groupi_n_10238);
  xnor csa_tree_add_51_79_groupi_g35632__2346(csa_tree_add_51_79_groupi_n_10470 ,csa_tree_add_51_79_groupi_n_10156 ,csa_tree_add_51_79_groupi_n_10229);
  xnor csa_tree_add_51_79_groupi_g35633__1666(csa_tree_add_51_79_groupi_n_10469 ,csa_tree_add_51_79_groupi_n_10163 ,csa_tree_add_51_79_groupi_n_10240);
  xnor csa_tree_add_51_79_groupi_g35634__7410(csa_tree_add_51_79_groupi_n_10467 ,csa_tree_add_51_79_groupi_n_10014 ,csa_tree_add_51_79_groupi_n_10237);
  xnor csa_tree_add_51_79_groupi_g35635__6417(csa_tree_add_51_79_groupi_n_10465 ,csa_tree_add_51_79_groupi_n_10088 ,csa_tree_add_51_79_groupi_n_10241);
  xnor csa_tree_add_51_79_groupi_g35636__5477(csa_tree_add_51_79_groupi_n_10464 ,csa_tree_add_51_79_groupi_n_10275 ,csa_tree_add_51_79_groupi_n_10246);
  xnor csa_tree_add_51_79_groupi_g35637__2398(csa_tree_add_51_79_groupi_n_10462 ,csa_tree_add_51_79_groupi_n_10137 ,csa_tree_add_51_79_groupi_n_10243);
  xnor csa_tree_add_51_79_groupi_g35638__5107(csa_tree_add_51_79_groupi_n_10461 ,csa_tree_add_51_79_groupi_n_9983 ,csa_tree_add_51_79_groupi_n_10247);
  xnor csa_tree_add_51_79_groupi_g35639__6260(csa_tree_add_51_79_groupi_n_10458 ,csa_tree_add_51_79_groupi_n_10011 ,csa_tree_add_51_79_groupi_n_10234);
  xnor csa_tree_add_51_79_groupi_g35640__4319(csa_tree_add_51_79_groupi_n_10456 ,csa_tree_add_51_79_groupi_n_10085 ,csa_tree_add_51_79_groupi_n_10242);
  not csa_tree_add_51_79_groupi_g35641(csa_tree_add_51_79_groupi_n_10428 ,csa_tree_add_51_79_groupi_n_10429);
  not csa_tree_add_51_79_groupi_g35642(csa_tree_add_51_79_groupi_n_10425 ,csa_tree_add_51_79_groupi_n_10426);
  not csa_tree_add_51_79_groupi_g35643(csa_tree_add_51_79_groupi_n_10421 ,csa_tree_add_51_79_groupi_n_10422);
  not csa_tree_add_51_79_groupi_g35644(csa_tree_add_51_79_groupi_n_10420 ,csa_tree_add_51_79_groupi_n_10419);
  or csa_tree_add_51_79_groupi_g35645__8428(csa_tree_add_51_79_groupi_n_10418 ,csa_tree_add_51_79_groupi_n_10339 ,csa_tree_add_51_79_groupi_n_10320);
  or csa_tree_add_51_79_groupi_g35646__5526(csa_tree_add_51_79_groupi_n_10417 ,csa_tree_add_51_79_groupi_n_10327 ,csa_tree_add_51_79_groupi_n_10271);
  or csa_tree_add_51_79_groupi_g35647__6783(csa_tree_add_51_79_groupi_n_10416 ,csa_tree_add_51_79_groupi_n_10090 ,csa_tree_add_51_79_groupi_n_10291);
  and csa_tree_add_51_79_groupi_g35648__3680(csa_tree_add_51_79_groupi_n_10415 ,csa_tree_add_51_79_groupi_n_10322 ,csa_tree_add_51_79_groupi_n_10214);
  or csa_tree_add_51_79_groupi_g35649__1617(csa_tree_add_51_79_groupi_n_10414 ,csa_tree_add_51_79_groupi_n_10322 ,csa_tree_add_51_79_groupi_n_10214);
  and csa_tree_add_51_79_groupi_g35650__2802(csa_tree_add_51_79_groupi_n_10413 ,csa_tree_add_51_79_groupi_n_10264 ,csa_tree_add_51_79_groupi_n_10265);
  and csa_tree_add_51_79_groupi_g35651__1705(csa_tree_add_51_79_groupi_n_10412 ,csa_tree_add_51_79_groupi_n_10274 ,csa_tree_add_51_79_groupi_n_10317);
  or csa_tree_add_51_79_groupi_g35652__5122(csa_tree_add_51_79_groupi_n_10411 ,csa_tree_add_51_79_groupi_n_10217 ,csa_tree_add_51_79_groupi_n_10289);
  or csa_tree_add_51_79_groupi_g35653__8246(csa_tree_add_51_79_groupi_n_10410 ,csa_tree_add_51_79_groupi_n_10264 ,csa_tree_add_51_79_groupi_n_10265);
  nor csa_tree_add_51_79_groupi_g35654__7098(csa_tree_add_51_79_groupi_n_10409 ,csa_tree_add_51_79_groupi_n_10311 ,csa_tree_add_51_79_groupi_n_10084);
  or csa_tree_add_51_79_groupi_g35655__6131(csa_tree_add_51_79_groupi_n_10408 ,csa_tree_add_51_79_groupi_n_10275 ,csa_tree_add_51_79_groupi_n_10200);
  or csa_tree_add_51_79_groupi_g35656__1881(csa_tree_add_51_79_groupi_n_10407 ,csa_tree_add_51_79_groupi_n_10309 ,csa_tree_add_51_79_groupi_n_10094);
  or csa_tree_add_51_79_groupi_g35657__5115(csa_tree_add_51_79_groupi_n_10406 ,csa_tree_add_51_79_groupi_n_10224 ,csa_tree_add_51_79_groupi_n_10303);
  or csa_tree_add_51_79_groupi_g35658__7482(csa_tree_add_51_79_groupi_n_10405 ,csa_tree_add_51_79_groupi_n_10259 ,csa_tree_add_51_79_groupi_n_10223);
  and csa_tree_add_51_79_groupi_g35659__4733(csa_tree_add_51_79_groupi_n_10404 ,csa_tree_add_51_79_groupi_n_10327 ,csa_tree_add_51_79_groupi_n_10271);
  or csa_tree_add_51_79_groupi_g35660__6161(csa_tree_add_51_79_groupi_n_10403 ,csa_tree_add_51_79_groupi_n_10338 ,csa_tree_add_51_79_groupi_n_10256);
  or csa_tree_add_51_79_groupi_g35661__9315(csa_tree_add_51_79_groupi_n_10402 ,csa_tree_add_51_79_groupi_n_10334 ,csa_tree_add_51_79_groupi_n_10272);
  or csa_tree_add_51_79_groupi_g35662__9945(csa_tree_add_51_79_groupi_n_10401 ,csa_tree_add_51_79_groupi_n_10333 ,csa_tree_add_51_79_groupi_n_10140);
  and csa_tree_add_51_79_groupi_g35663__2883(csa_tree_add_51_79_groupi_n_10400 ,csa_tree_add_51_79_groupi_n_10333 ,csa_tree_add_51_79_groupi_n_10140);
  and csa_tree_add_51_79_groupi_g35664__2346(csa_tree_add_51_79_groupi_n_10399 ,csa_tree_add_51_79_groupi_n_10334 ,csa_tree_add_51_79_groupi_n_10272);
  or csa_tree_add_51_79_groupi_g35665__1666(csa_tree_add_51_79_groupi_n_10398 ,csa_tree_add_51_79_groupi_n_10286 ,csa_tree_add_51_79_groupi_n_10077);
  or csa_tree_add_51_79_groupi_g35666__7410(csa_tree_add_51_79_groupi_n_10397 ,csa_tree_add_51_79_groupi_n_10096 ,csa_tree_add_51_79_groupi_n_10285);
  or csa_tree_add_51_79_groupi_g35667__6417(csa_tree_add_51_79_groupi_n_10396 ,csa_tree_add_51_79_groupi_n_10182 ,csa_tree_add_51_79_groupi_n_10279);
  nor csa_tree_add_51_79_groupi_g35668__5477(csa_tree_add_51_79_groupi_n_10395 ,csa_tree_add_51_79_groupi_n_10332 ,csa_tree_add_51_79_groupi_n_10267);
  and csa_tree_add_51_79_groupi_g35669__2398(csa_tree_add_51_79_groupi_n_10394 ,csa_tree_add_51_79_groupi_n_10332 ,csa_tree_add_51_79_groupi_n_10267);
  or csa_tree_add_51_79_groupi_g35670__5107(csa_tree_add_51_79_groupi_n_10393 ,csa_tree_add_51_79_groupi_n_10220 ,csa_tree_add_51_79_groupi_n_10296);
  and csa_tree_add_51_79_groupi_g35671__6260(csa_tree_add_51_79_groupi_n_10437 ,csa_tree_add_51_79_groupi_n_10321 ,csa_tree_add_51_79_groupi_n_10209);
  and csa_tree_add_51_79_groupi_g35672__4319(csa_tree_add_51_79_groupi_n_10436 ,csa_tree_add_51_79_groupi_n_10185 ,csa_tree_add_51_79_groupi_n_10299);
  and csa_tree_add_51_79_groupi_g35673__8428(csa_tree_add_51_79_groupi_n_10435 ,csa_tree_add_51_79_groupi_n_10115 ,csa_tree_add_51_79_groupi_n_10306);
  and csa_tree_add_51_79_groupi_g35674__5526(csa_tree_add_51_79_groupi_n_10434 ,csa_tree_add_51_79_groupi_n_10171 ,csa_tree_add_51_79_groupi_n_10298);
  and csa_tree_add_51_79_groupi_g35675__6783(csa_tree_add_51_79_groupi_n_10433 ,csa_tree_add_51_79_groupi_n_10301 ,csa_tree_add_51_79_groupi_n_10190);
  and csa_tree_add_51_79_groupi_g35676__3680(csa_tree_add_51_79_groupi_n_10432 ,csa_tree_add_51_79_groupi_n_10174 ,csa_tree_add_51_79_groupi_n_10288);
  and csa_tree_add_51_79_groupi_g35677__1617(csa_tree_add_51_79_groupi_n_10431 ,csa_tree_add_51_79_groupi_n_10294 ,csa_tree_add_51_79_groupi_n_10113);
  and csa_tree_add_51_79_groupi_g35678__2802(csa_tree_add_51_79_groupi_n_10430 ,csa_tree_add_51_79_groupi_n_10194 ,csa_tree_add_51_79_groupi_n_10295);
  and csa_tree_add_51_79_groupi_g35679__1705(csa_tree_add_51_79_groupi_n_10429 ,csa_tree_add_51_79_groupi_n_10177 ,csa_tree_add_51_79_groupi_n_10293);
  and csa_tree_add_51_79_groupi_g35680__5122(csa_tree_add_51_79_groupi_n_10427 ,csa_tree_add_51_79_groupi_n_10187 ,csa_tree_add_51_79_groupi_n_10300);
  and csa_tree_add_51_79_groupi_g35681__8246(csa_tree_add_51_79_groupi_n_10426 ,csa_tree_add_51_79_groupi_n_10312 ,csa_tree_add_51_79_groupi_n_10165);
  and csa_tree_add_51_79_groupi_g35682__7098(csa_tree_add_51_79_groupi_n_10424 ,csa_tree_add_51_79_groupi_n_10308 ,csa_tree_add_51_79_groupi_n_10198);
  and csa_tree_add_51_79_groupi_g35683__6131(csa_tree_add_51_79_groupi_n_10423 ,csa_tree_add_51_79_groupi_n_10313 ,csa_tree_add_51_79_groupi_n_10205);
  or csa_tree_add_51_79_groupi_g35684__1881(csa_tree_add_51_79_groupi_n_10422 ,csa_tree_add_51_79_groupi_n_10126 ,csa_tree_add_51_79_groupi_n_10319);
  and csa_tree_add_51_79_groupi_g35685__5115(csa_tree_add_51_79_groupi_n_10419 ,csa_tree_add_51_79_groupi_n_10304 ,csa_tree_add_51_79_groupi_n_10196);
  not csa_tree_add_51_79_groupi_g35686(csa_tree_add_51_79_groupi_n_10388 ,csa_tree_add_51_79_groupi_n_10387);
  not csa_tree_add_51_79_groupi_g35687(csa_tree_add_51_79_groupi_n_10383 ,csa_tree_add_51_79_groupi_n_10382);
  not csa_tree_add_51_79_groupi_g35688(csa_tree_add_51_79_groupi_n_10381 ,csa_tree_add_51_79_groupi_n_10380);
  not csa_tree_add_51_79_groupi_g35689(csa_tree_add_51_79_groupi_n_10378 ,csa_tree_add_51_79_groupi_n_10377);
  not csa_tree_add_51_79_groupi_g35690(csa_tree_add_51_79_groupi_n_10376 ,csa_tree_add_51_79_groupi_n_10375);
  not csa_tree_add_51_79_groupi_g35691(csa_tree_add_51_79_groupi_n_10373 ,csa_tree_add_51_79_groupi_n_10372);
  not csa_tree_add_51_79_groupi_g35692(csa_tree_add_51_79_groupi_n_10369 ,csa_tree_add_51_79_groupi_n_10368);
  not csa_tree_add_51_79_groupi_g35693(csa_tree_add_51_79_groupi_n_10365 ,csa_tree_add_51_79_groupi_n_10366);
  and csa_tree_add_51_79_groupi_g35694__7482(csa_tree_add_51_79_groupi_n_10364 ,csa_tree_add_51_79_groupi_n_10282 ,csa_tree_add_51_79_groupi_n_10249);
  and csa_tree_add_51_79_groupi_g35695__4733(csa_tree_add_51_79_groupi_n_10363 ,csa_tree_add_51_79_groupi_n_9999 ,csa_tree_add_51_79_groupi_n_10336);
  or csa_tree_add_51_79_groupi_g35696__6161(csa_tree_add_51_79_groupi_n_10362 ,csa_tree_add_51_79_groupi_n_9999 ,csa_tree_add_51_79_groupi_n_10336);
  or csa_tree_add_51_79_groupi_g35697__9315(csa_tree_add_51_79_groupi_n_10361 ,csa_tree_add_51_79_groupi_n_10161 ,csa_tree_add_51_79_groupi_n_10270);
  and csa_tree_add_51_79_groupi_g35698__9945(csa_tree_add_51_79_groupi_n_10360 ,csa_tree_add_51_79_groupi_n_10161 ,csa_tree_add_51_79_groupi_n_10270);
  or csa_tree_add_51_79_groupi_g35699__2883(csa_tree_add_51_79_groupi_n_10359 ,csa_tree_add_51_79_groupi_n_10250 ,csa_tree_add_51_79_groupi_n_10095);
  or csa_tree_add_51_79_groupi_g35700__2346(csa_tree_add_51_79_groupi_n_10358 ,csa_tree_add_51_79_groupi_n_9869 ,csa_tree_add_51_79_groupi_n_10253);
  xnor csa_tree_add_51_79_groupi_g35701__1666(csa_tree_add_51_79_groupi_n_10357 ,csa_tree_add_51_79_groupi_n_10224 ,csa_tree_add_51_79_groupi_n_9862);
  xnor csa_tree_add_51_79_groupi_g35702__7410(csa_tree_add_51_79_groupi_n_10356 ,csa_tree_add_51_79_groupi_n_10133 ,csa_tree_add_51_79_groupi_n_10075);
  xnor csa_tree_add_51_79_groupi_g35703__6417(csa_tree_add_51_79_groupi_n_10355 ,csa_tree_add_51_79_groupi_n_9795 ,csa_tree_add_51_79_groupi_n_10216);
  xnor csa_tree_add_51_79_groupi_g35704__5477(csa_tree_add_51_79_groupi_n_10354 ,csa_tree_add_51_79_groupi_n_10131 ,csa_tree_add_51_79_groupi_n_10082);
  xnor csa_tree_add_51_79_groupi_g35705__2398(csa_tree_add_51_79_groupi_n_10353 ,csa_tree_add_51_79_groupi_n_9989 ,csa_tree_add_51_79_groupi_n_10221);
  xnor csa_tree_add_51_79_groupi_g35706__5107(csa_tree_add_51_79_groupi_n_10352 ,csa_tree_add_51_79_groupi_n_10147 ,csa_tree_add_51_79_groupi_n_10146);
  xnor csa_tree_add_51_79_groupi_g35707__6260(csa_tree_add_51_79_groupi_n_10351 ,csa_tree_add_51_79_groupi_n_10141 ,csa_tree_add_51_79_groupi_n_10217);
  xnor csa_tree_add_51_79_groupi_g35708__4319(csa_tree_add_51_79_groupi_n_10350 ,csa_tree_add_51_79_groupi_n_10144 ,csa_tree_add_51_79_groupi_n_10073);
  xnor csa_tree_add_51_79_groupi_g35709__8428(csa_tree_add_51_79_groupi_n_10349 ,csa_tree_add_51_79_groupi_n_9982 ,csa_tree_add_51_79_groupi_n_10130);
  xnor csa_tree_add_51_79_groupi_g35710__5526(csa_tree_add_51_79_groupi_n_10348 ,csa_tree_add_51_79_groupi_n_10143 ,csa_tree_add_51_79_groupi_n_10127);
  xnor csa_tree_add_51_79_groupi_g35711__6783(csa_tree_add_51_79_groupi_n_10347 ,csa_tree_add_51_79_groupi_n_9866 ,csa_tree_add_51_79_groupi_n_10151);
  xnor csa_tree_add_51_79_groupi_g35712__3680(csa_tree_add_51_79_groupi_n_10346 ,csa_tree_add_51_79_groupi_n_10162 ,csa_tree_add_51_79_groupi_n_10084);
  xnor csa_tree_add_51_79_groupi_g35713__1617(csa_tree_add_51_79_groupi_n_10345 ,csa_tree_add_51_79_groupi_n_10149 ,csa_tree_add_51_79_groupi_n_10132);
  xnor csa_tree_add_51_79_groupi_g35714__2802(csa_tree_add_51_79_groupi_n_10344 ,csa_tree_add_51_79_groupi_n_10005 ,csa_tree_add_51_79_groupi_n_10142);
  xnor csa_tree_add_51_79_groupi_g35715__1705(csa_tree_add_51_79_groupi_n_10343 ,csa_tree_add_51_79_groupi_n_10161 ,csa_tree_add_51_79_groupi_n_10222);
  xnor csa_tree_add_51_79_groupi_g35716__5122(csa_tree_add_51_79_groupi_n_10392 ,csa_tree_add_51_79_groupi_n_31 ,csa_tree_add_51_79_groupi_n_10101);
  xnor csa_tree_add_51_79_groupi_g35717__8246(csa_tree_add_51_79_groupi_n_10391 ,csa_tree_add_51_79_groupi_n_9676 ,csa_tree_add_51_79_groupi_n_10109);
  xnor csa_tree_add_51_79_groupi_g35718__7098(csa_tree_add_51_79_groupi_n_10390 ,csa_tree_add_51_79_groupi_n_9873 ,csa_tree_add_51_79_groupi_n_10103);
  and csa_tree_add_51_79_groupi_g35719__6131(csa_tree_add_51_79_groupi_n_10389 ,csa_tree_add_51_79_groupi_n_10254 ,csa_tree_add_51_79_groupi_n_10116);
  or csa_tree_add_51_79_groupi_g35720__1881(csa_tree_add_51_79_groupi_n_10387 ,csa_tree_add_51_79_groupi_n_10257 ,csa_tree_add_51_79_groupi_n_10121);
  xnor csa_tree_add_51_79_groupi_g35721__5115(csa_tree_add_51_79_groupi_n_10386 ,csa_tree_add_51_79_groupi_n_10021 ,csa_tree_add_51_79_groupi_n_10106);
  xnor csa_tree_add_51_79_groupi_g35722__7482(csa_tree_add_51_79_groupi_n_10385 ,csa_tree_add_51_79_groupi_n_9864 ,csa_tree_add_51_79_groupi_n_10099);
  xnor csa_tree_add_51_79_groupi_g35723__4733(csa_tree_add_51_79_groupi_n_10384 ,csa_tree_add_51_79_groupi_n_9936 ,csa_tree_add_51_79_groupi_n_10110);
  xnor csa_tree_add_51_79_groupi_g35724__6161(csa_tree_add_51_79_groupi_n_10382 ,csa_tree_add_51_79_groupi_n_10080 ,csa_tree_add_51_79_groupi_n_10102);
  xnor csa_tree_add_51_79_groupi_g35725__9315(csa_tree_add_51_79_groupi_n_10380 ,csa_tree_add_51_79_groupi_n_10087 ,csa_tree_add_51_79_groupi_n_10111);
  xnor csa_tree_add_51_79_groupi_g35726__9945(csa_tree_add_51_79_groupi_n_10379 ,csa_tree_add_51_79_groupi_n_10025 ,csa_tree_add_51_79_groupi_n_10105);
  xnor csa_tree_add_51_79_groupi_g35727__2883(csa_tree_add_51_79_groupi_n_10377 ,csa_tree_add_51_79_groupi_n_9941 ,csa_tree_add_51_79_groupi_n_10112);
  xnor csa_tree_add_51_79_groupi_g35728__2346(csa_tree_add_51_79_groupi_n_10375 ,csa_tree_add_51_79_groupi_n_9985 ,csa_tree_add_51_79_groupi_n_10107);
  xnor csa_tree_add_51_79_groupi_g35729__1666(csa_tree_add_51_79_groupi_n_10374 ,csa_tree_add_51_79_groupi_n_9930 ,csa_tree_add_51_79_groupi_n_10098);
  xnor csa_tree_add_51_79_groupi_g35730__7410(csa_tree_add_51_79_groupi_n_10372 ,csa_tree_add_51_79_groupi_n_9984 ,csa_tree_add_51_79_groupi_n_10100);
  xnor csa_tree_add_51_79_groupi_g35731__6417(csa_tree_add_51_79_groupi_n_10371 ,csa_tree_add_51_79_groupi_n_9937 ,csa_tree_add_51_79_groupi_n_10108);
  xnor csa_tree_add_51_79_groupi_g35732__5477(csa_tree_add_51_79_groupi_n_10370 ,csa_tree_add_51_79_groupi_n_9870 ,csa_tree_add_51_79_groupi_n_10097);
  and csa_tree_add_51_79_groupi_g35733__2398(csa_tree_add_51_79_groupi_n_10368 ,csa_tree_add_51_79_groupi_n_10119 ,csa_tree_add_51_79_groupi_n_10255);
  xnor csa_tree_add_51_79_groupi_g35734__5107(csa_tree_add_51_79_groupi_n_10367 ,csa_tree_add_51_79_groupi_n_9939 ,csa_tree_add_51_79_groupi_n_10104);
  and csa_tree_add_51_79_groupi_g35735__6260(csa_tree_add_51_79_groupi_n_10366 ,csa_tree_add_51_79_groupi_n_10248 ,csa_tree_add_51_79_groupi_n_10188);
  not csa_tree_add_51_79_groupi_g35736(csa_tree_add_51_79_groupi_n_10330 ,csa_tree_add_51_79_groupi_n_10331);
  not csa_tree_add_51_79_groupi_g35737(csa_tree_add_51_79_groupi_n_10329 ,csa_tree_add_51_79_groupi_n_10328);
  not csa_tree_add_51_79_groupi_g35738(csa_tree_add_51_79_groupi_n_10326 ,csa_tree_add_51_79_groupi_n_10325);
  not csa_tree_add_51_79_groupi_g35739(csa_tree_add_51_79_groupi_n_10324 ,csa_tree_add_51_79_groupi_n_10323);
  or csa_tree_add_51_79_groupi_g35740__4319(csa_tree_add_51_79_groupi_n_10321 ,csa_tree_add_51_79_groupi_n_9947 ,csa_tree_add_51_79_groupi_n_10207);
  and csa_tree_add_51_79_groupi_g35741__8428(csa_tree_add_51_79_groupi_n_10320 ,csa_tree_add_51_79_groupi_n_10127 ,csa_tree_add_51_79_groupi_n_10143);
  and csa_tree_add_51_79_groupi_g35742__5526(csa_tree_add_51_79_groupi_n_10319 ,csa_tree_add_51_79_groupi_n_10125 ,csa_tree_add_51_79_groupi_n_10089);
  and csa_tree_add_51_79_groupi_g35743__6783(csa_tree_add_51_79_groupi_n_10318 ,csa_tree_add_51_79_groupi_n_10149 ,csa_tree_add_51_79_groupi_n_10132);
  or csa_tree_add_51_79_groupi_g35744__3680(csa_tree_add_51_79_groupi_n_10317 ,csa_tree_add_51_79_groupi_n_10149 ,csa_tree_add_51_79_groupi_n_10132);
  and csa_tree_add_51_79_groupi_g35745__1617(csa_tree_add_51_79_groupi_n_10316 ,csa_tree_add_51_79_groupi_n_10130 ,csa_tree_add_51_79_groupi_n_9982);
  or csa_tree_add_51_79_groupi_g35746__2802(csa_tree_add_51_79_groupi_n_10315 ,csa_tree_add_51_79_groupi_n_9794 ,csa_tree_add_51_79_groupi_n_10215);
  nor csa_tree_add_51_79_groupi_g35747__1705(csa_tree_add_51_79_groupi_n_10314 ,csa_tree_add_51_79_groupi_n_9795 ,csa_tree_add_51_79_groupi_n_10216);
  or csa_tree_add_51_79_groupi_g35748__5122(csa_tree_add_51_79_groupi_n_10313 ,csa_tree_add_51_79_groupi_n_10018 ,csa_tree_add_51_79_groupi_n_10206);
  or csa_tree_add_51_79_groupi_g35749__8246(csa_tree_add_51_79_groupi_n_10312 ,csa_tree_add_51_79_groupi_n_10083 ,csa_tree_add_51_79_groupi_n_10166);
  nor csa_tree_add_51_79_groupi_g35750__7098(csa_tree_add_51_79_groupi_n_10311 ,csa_tree_add_51_79_groupi_n_10152 ,csa_tree_add_51_79_groupi_n_10162);
  and csa_tree_add_51_79_groupi_g35751__6131(csa_tree_add_51_79_groupi_n_10310 ,csa_tree_add_51_79_groupi_n_10152 ,csa_tree_add_51_79_groupi_n_10162);
  and csa_tree_add_51_79_groupi_g35752__1881(csa_tree_add_51_79_groupi_n_10309 ,csa_tree_add_51_79_groupi_n_9978 ,csa_tree_add_51_79_groupi_n_10156);
  or csa_tree_add_51_79_groupi_g35753__5115(csa_tree_add_51_79_groupi_n_10308 ,csa_tree_add_51_79_groupi_n_10092 ,csa_tree_add_51_79_groupi_n_10199);
  or csa_tree_add_51_79_groupi_g35754__7482(csa_tree_add_51_79_groupi_n_10307 ,csa_tree_add_51_79_groupi_n_9978 ,csa_tree_add_51_79_groupi_n_10156);
  or csa_tree_add_51_79_groupi_g35755__4733(csa_tree_add_51_79_groupi_n_10306 ,csa_tree_add_51_79_groupi_n_10114 ,csa_tree_add_51_79_groupi_n_10088);
  or csa_tree_add_51_79_groupi_g35756__6161(csa_tree_add_51_79_groupi_n_10305 ,csa_tree_add_51_79_groupi_n_9862 ,csa_tree_add_51_79_groupi_n_10155);
  or csa_tree_add_51_79_groupi_g35757__9315(csa_tree_add_51_79_groupi_n_10304 ,csa_tree_add_51_79_groupi_n_10197 ,csa_tree_add_51_79_groupi_n_10086);
  and csa_tree_add_51_79_groupi_g35758__9945(csa_tree_add_51_79_groupi_n_10303 ,csa_tree_add_51_79_groupi_n_9862 ,csa_tree_add_51_79_groupi_n_10155);
  or csa_tree_add_51_79_groupi_g35759__2883(csa_tree_add_51_79_groupi_n_10302 ,csa_tree_add_51_79_groupi_n_10127 ,csa_tree_add_51_79_groupi_n_10143);
  or csa_tree_add_51_79_groupi_g35760__2346(csa_tree_add_51_79_groupi_n_10301 ,csa_tree_add_51_79_groupi_n_10022 ,csa_tree_add_51_79_groupi_n_10191);
  or csa_tree_add_51_79_groupi_g35761__1666(csa_tree_add_51_79_groupi_n_10300 ,csa_tree_add_51_79_groupi_n_10186 ,csa_tree_add_51_79_groupi_n_10024);
  or csa_tree_add_51_79_groupi_g35762__7410(csa_tree_add_51_79_groupi_n_10299 ,csa_tree_add_51_79_groupi_n_10184 ,csa_tree_add_51_79_groupi_n_10163);
  or csa_tree_add_51_79_groupi_g35763__6417(csa_tree_add_51_79_groupi_n_10298 ,csa_tree_add_51_79_groupi_n_9802 ,csa_tree_add_51_79_groupi_n_10170);
  or csa_tree_add_51_79_groupi_g35764__5477(csa_tree_add_51_79_groupi_n_10297 ,csa_tree_add_51_79_groupi_n_10075 ,csa_tree_add_51_79_groupi_n_10133);
  and csa_tree_add_51_79_groupi_g35765__2398(csa_tree_add_51_79_groupi_n_10296 ,csa_tree_add_51_79_groupi_n_10075 ,csa_tree_add_51_79_groupi_n_10133);
  or csa_tree_add_51_79_groupi_g35766__5107(csa_tree_add_51_79_groupi_n_10295 ,csa_tree_add_51_79_groupi_n_10203 ,csa_tree_add_51_79_groupi_n_10221);
  or csa_tree_add_51_79_groupi_g35767__6260(csa_tree_add_51_79_groupi_n_10294 ,csa_tree_add_51_79_groupi_n_10093 ,csa_tree_add_51_79_groupi_n_10212);
  or csa_tree_add_51_79_groupi_g35768__4319(csa_tree_add_51_79_groupi_n_10293 ,csa_tree_add_51_79_groupi_n_10081 ,csa_tree_add_51_79_groupi_n_10178);
  or csa_tree_add_51_79_groupi_g35769__8428(csa_tree_add_51_79_groupi_n_10292 ,csa_tree_add_51_79_groupi_n_10134 ,csa_tree_add_51_79_groupi_n_10002);
  and csa_tree_add_51_79_groupi_g35770__5526(csa_tree_add_51_79_groupi_n_10291 ,csa_tree_add_51_79_groupi_n_10134 ,csa_tree_add_51_79_groupi_n_10002);
  or csa_tree_add_51_79_groupi_g35771__6783(csa_tree_add_51_79_groupi_n_10290 ,csa_tree_add_51_79_groupi_n_10145 ,csa_tree_add_51_79_groupi_n_10141);
  and csa_tree_add_51_79_groupi_g35772__3680(csa_tree_add_51_79_groupi_n_10289 ,csa_tree_add_51_79_groupi_n_10145 ,csa_tree_add_51_79_groupi_n_10141);
  or csa_tree_add_51_79_groupi_g35773__1617(csa_tree_add_51_79_groupi_n_10288 ,csa_tree_add_51_79_groupi_n_10173 ,csa_tree_add_51_79_groupi_n_10091);
  or csa_tree_add_51_79_groupi_g35774__2802(csa_tree_add_51_79_groupi_n_10287 ,csa_tree_add_51_79_groupi_n_10073 ,csa_tree_add_51_79_groupi_n_10144);
  and csa_tree_add_51_79_groupi_g35775__1705(csa_tree_add_51_79_groupi_n_10286 ,csa_tree_add_51_79_groupi_n_10073 ,csa_tree_add_51_79_groupi_n_10144);
  nor csa_tree_add_51_79_groupi_g35776__5122(csa_tree_add_51_79_groupi_n_10285 ,csa_tree_add_51_79_groupi_n_10137 ,csa_tree_add_51_79_groupi_n_10068);
  or csa_tree_add_51_79_groupi_g35777__8246(csa_tree_add_51_79_groupi_n_10284 ,csa_tree_add_51_79_groupi_n_10136 ,csa_tree_add_51_79_groupi_n_10067);
  or csa_tree_add_51_79_groupi_g35778__7098(csa_tree_add_51_79_groupi_n_10283 ,csa_tree_add_51_79_groupi_n_10130 ,csa_tree_add_51_79_groupi_n_9982);
  or csa_tree_add_51_79_groupi_g35779__6131(csa_tree_add_51_79_groupi_n_10342 ,csa_tree_add_51_79_groupi_n_10183 ,csa_tree_add_51_79_groupi_n_9968);
  and csa_tree_add_51_79_groupi_g35780__1881(csa_tree_add_51_79_groupi_n_10341 ,csa_tree_add_51_79_groupi_n_10034 ,csa_tree_add_51_79_groupi_n_10189);
  and csa_tree_add_51_79_groupi_g35781__5115(csa_tree_add_51_79_groupi_n_10340 ,csa_tree_add_51_79_groupi_n_9843 ,csa_tree_add_51_79_groupi_n_10167);
  and csa_tree_add_51_79_groupi_g35782__7482(csa_tree_add_51_79_groupi_n_10339 ,csa_tree_add_51_79_groupi_n_10038 ,csa_tree_add_51_79_groupi_n_10193);
  and csa_tree_add_51_79_groupi_g35783__4733(csa_tree_add_51_79_groupi_n_10338 ,csa_tree_add_51_79_groupi_n_10036 ,csa_tree_add_51_79_groupi_n_10192);
  and csa_tree_add_51_79_groupi_g35784__6161(csa_tree_add_51_79_groupi_n_10337 ,csa_tree_add_51_79_groupi_n_10030 ,csa_tree_add_51_79_groupi_n_10181);
  and csa_tree_add_51_79_groupi_g35785__9315(csa_tree_add_51_79_groupi_n_10336 ,csa_tree_add_51_79_groupi_n_10044 ,csa_tree_add_51_79_groupi_n_10175);
  and csa_tree_add_51_79_groupi_g35786__9945(csa_tree_add_51_79_groupi_n_10335 ,csa_tree_add_51_79_groupi_n_10026 ,csa_tree_add_51_79_groupi_n_10176);
  and csa_tree_add_51_79_groupi_g35787__2883(csa_tree_add_51_79_groupi_n_10334 ,csa_tree_add_51_79_groupi_n_10052 ,csa_tree_add_51_79_groupi_n_10172);
  and csa_tree_add_51_79_groupi_g35788__2346(csa_tree_add_51_79_groupi_n_10333 ,csa_tree_add_51_79_groupi_n_9976 ,csa_tree_add_51_79_groupi_n_10179);
  and csa_tree_add_51_79_groupi_g35789__1666(csa_tree_add_51_79_groupi_n_10332 ,csa_tree_add_51_79_groupi_n_9974 ,csa_tree_add_51_79_groupi_n_10169);
  and csa_tree_add_51_79_groupi_g35790__7410(csa_tree_add_51_79_groupi_n_10331 ,csa_tree_add_51_79_groupi_n_10048 ,csa_tree_add_51_79_groupi_n_10168);
  or csa_tree_add_51_79_groupi_g35791__6417(csa_tree_add_51_79_groupi_n_10328 ,csa_tree_add_51_79_groupi_n_10041 ,csa_tree_add_51_79_groupi_n_10210);
  and csa_tree_add_51_79_groupi_g35792__5477(csa_tree_add_51_79_groupi_n_10327 ,csa_tree_add_51_79_groupi_n_10045 ,csa_tree_add_51_79_groupi_n_10195);
  and csa_tree_add_51_79_groupi_g35793__2398(csa_tree_add_51_79_groupi_n_10325 ,csa_tree_add_51_79_groupi_n_10051 ,csa_tree_add_51_79_groupi_n_10202);
  and csa_tree_add_51_79_groupi_g35794__5107(csa_tree_add_51_79_groupi_n_10323 ,csa_tree_add_51_79_groupi_n_10208 ,csa_tree_add_51_79_groupi_n_10050);
  and csa_tree_add_51_79_groupi_g35795__6260(csa_tree_add_51_79_groupi_n_10322 ,csa_tree_add_51_79_groupi_n_10211 ,csa_tree_add_51_79_groupi_n_9964);
  not csa_tree_add_51_79_groupi_g35796(csa_tree_add_51_79_groupi_n_10269 ,csa_tree_add_51_79_groupi_n_10268);
  not csa_tree_add_51_79_groupi_g35797(csa_tree_add_51_79_groupi_n_10262 ,csa_tree_add_51_79_groupi_n_10263);
  and csa_tree_add_51_79_groupi_g35798__4319(csa_tree_add_51_79_groupi_n_10261 ,csa_tree_add_51_79_groupi_n_10147 ,csa_tree_add_51_79_groupi_n_10146);
  or csa_tree_add_51_79_groupi_g35799__8428(csa_tree_add_51_79_groupi_n_10260 ,csa_tree_add_51_79_groupi_n_10142 ,csa_tree_add_51_79_groupi_n_10005);
  and csa_tree_add_51_79_groupi_g35800__5526(csa_tree_add_51_79_groupi_n_10259 ,csa_tree_add_51_79_groupi_n_10142 ,csa_tree_add_51_79_groupi_n_10005);
  or csa_tree_add_51_79_groupi_g35801__6783(csa_tree_add_51_79_groupi_n_10258 ,csa_tree_add_51_79_groupi_n_10157 ,csa_tree_add_51_79_groupi_n_10153);
  nor csa_tree_add_51_79_groupi_g35802__3680(csa_tree_add_51_79_groupi_n_10257 ,csa_tree_add_51_79_groupi_n_10219 ,csa_tree_add_51_79_groupi_n_10123);
  nor csa_tree_add_51_79_groupi_g35803__1617(csa_tree_add_51_79_groupi_n_10256 ,csa_tree_add_51_79_groupi_n_10158 ,csa_tree_add_51_79_groupi_n_10154);
  or csa_tree_add_51_79_groupi_g35804__2802(csa_tree_add_51_79_groupi_n_10255 ,csa_tree_add_51_79_groupi_n_10118 ,csa_tree_add_51_79_groupi_n_10020);
  or csa_tree_add_51_79_groupi_g35805__1705(csa_tree_add_51_79_groupi_n_10254 ,csa_tree_add_51_79_groupi_n_9940 ,csa_tree_add_51_79_groupi_n_10117);
  nor csa_tree_add_51_79_groupi_g35806__5122(csa_tree_add_51_79_groupi_n_10253 ,csa_tree_add_51_79_groupi_n_9866 ,csa_tree_add_51_79_groupi_n_10151);
  or csa_tree_add_51_79_groupi_g35807__8246(csa_tree_add_51_79_groupi_n_10252 ,csa_tree_add_51_79_groupi_n_32 ,csa_tree_add_51_79_groupi_n_10150);
  or csa_tree_add_51_79_groupi_g35808__7098(csa_tree_add_51_79_groupi_n_10251 ,csa_tree_add_51_79_groupi_n_10016 ,csa_tree_add_51_79_groupi_n_10148);
  and csa_tree_add_51_79_groupi_g35809__6131(csa_tree_add_51_79_groupi_n_10250 ,csa_tree_add_51_79_groupi_n_10016 ,csa_tree_add_51_79_groupi_n_10148);
  or csa_tree_add_51_79_groupi_g35810__1881(csa_tree_add_51_79_groupi_n_10249 ,csa_tree_add_51_79_groupi_n_10147 ,csa_tree_add_51_79_groupi_n_10146);
  or csa_tree_add_51_79_groupi_g35811__5115(csa_tree_add_51_79_groupi_n_10248 ,csa_tree_add_51_79_groupi_n_10079 ,csa_tree_add_51_79_groupi_n_10180);
  xnor csa_tree_add_51_79_groupi_g35812__7482(csa_tree_add_51_79_groupi_n_10247 ,csa_tree_add_51_79_groupi_n_10092 ,csa_tree_add_51_79_groupi_n_9935);
  xnor csa_tree_add_51_79_groupi_g35813__4733(csa_tree_add_51_79_groupi_n_10246 ,csa_tree_add_51_79_groupi_n_10064 ,csa_tree_add_51_79_groupi_n_9991);
  xnor csa_tree_add_51_79_groupi_g35814__6161(csa_tree_add_51_79_groupi_n_10245 ,csa_tree_add_51_79_groupi_n_9998 ,csa_tree_add_51_79_groupi_n_10063);
  xnor csa_tree_add_51_79_groupi_g35815__9315(csa_tree_add_51_79_groupi_n_10244 ,csa_tree_add_51_79_groupi_n_9444 ,csa_tree_add_51_79_groupi_n_10023);
  xnor csa_tree_add_51_79_groupi_g35816__9945(csa_tree_add_51_79_groupi_n_10243 ,csa_tree_add_51_79_groupi_n_10096 ,csa_tree_add_51_79_groupi_n_10068);
  xnor csa_tree_add_51_79_groupi_g35817__2883(csa_tree_add_51_79_groupi_n_10242 ,csa_tree_add_51_79_groupi_n_10070 ,csa_tree_add_51_79_groupi_n_10017);
  xnor csa_tree_add_51_79_groupi_g35818__2346(csa_tree_add_51_79_groupi_n_10241 ,csa_tree_add_51_79_groupi_n_10066 ,csa_tree_add_51_79_groupi_n_9981);
  xnor csa_tree_add_51_79_groupi_g35819__1666(csa_tree_add_51_79_groupi_n_10240 ,csa_tree_add_51_79_groupi_n_10000 ,csa_tree_add_51_79_groupi_n_9925);
  xnor csa_tree_add_51_79_groupi_g35820__7410(csa_tree_add_51_79_groupi_n_10239 ,csa_tree_add_51_79_groupi_n_10001 ,csa_tree_add_51_79_groupi_n_10060);
  xnor csa_tree_add_51_79_groupi_g35821__6417(csa_tree_add_51_79_groupi_n_10238 ,csa_tree_add_51_79_groupi_n_10002 ,csa_tree_add_51_79_groupi_n_10090);
  xnor csa_tree_add_51_79_groupi_g35822__5477(csa_tree_add_51_79_groupi_n_10237 ,csa_tree_add_51_79_groupi_n_9679 ,csa_tree_add_51_79_groupi_n_10093);
  xnor csa_tree_add_51_79_groupi_g35823__2398(csa_tree_add_51_79_groupi_n_10236 ,csa_tree_add_51_79_groupi_n_10015 ,csa_tree_add_51_79_groupi_n_10095);
  xnor csa_tree_add_51_79_groupi_g35824__5107(csa_tree_add_51_79_groupi_n_10235 ,csa_tree_add_51_79_groupi_n_10062 ,csa_tree_add_51_79_groupi_n_9993);
  xnor csa_tree_add_51_79_groupi_g35825__6260(csa_tree_add_51_79_groupi_n_10234 ,csa_tree_add_51_79_groupi_n_10079 ,csa_tree_add_51_79_groupi_n_9922);
  xnor csa_tree_add_51_79_groupi_g35826__4319(csa_tree_add_51_79_groupi_n_10233 ,csa_tree_add_51_79_groupi_n_10008 ,csa_tree_add_51_79_groupi_n_10004);
  xnor csa_tree_add_51_79_groupi_g35827__8428(csa_tree_add_51_79_groupi_n_10232 ,csa_tree_add_51_79_groupi_n_9855 ,csa_tree_add_51_79_groupi_n_10019);
  xnor csa_tree_add_51_79_groupi_g35828__5526(csa_tree_add_51_79_groupi_n_10231 ,csa_tree_add_51_79_groupi_n_9997 ,csa_tree_add_51_79_groupi_n_9995);
  xnor csa_tree_add_51_79_groupi_g35829__6783(csa_tree_add_51_79_groupi_n_10230 ,csa_tree_add_51_79_groupi_n_10006 ,csa_tree_add_51_79_groupi_n_9861);
  xnor csa_tree_add_51_79_groupi_g35830__3680(csa_tree_add_51_79_groupi_n_10229 ,csa_tree_add_51_79_groupi_n_10094 ,csa_tree_add_51_79_groupi_n_9978);
  xnor csa_tree_add_51_79_groupi_g35831__1617(csa_tree_add_51_79_groupi_n_10228 ,csa_tree_add_51_79_groupi_n_10022 ,csa_tree_add_51_79_groupi_n_10071);
  xnor csa_tree_add_51_79_groupi_g35832__2802(csa_tree_add_51_79_groupi_n_10227 ,csa_tree_add_51_79_groupi_n_9979 ,csa_tree_add_51_79_groupi_n_10018);
  xnor csa_tree_add_51_79_groupi_g35833__1705(csa_tree_add_51_79_groupi_n_10226 ,csa_tree_add_51_79_groupi_n_10012 ,csa_tree_add_51_79_groupi_n_9990);
  xnor csa_tree_add_51_79_groupi_g35834__5122(csa_tree_add_51_79_groupi_n_10225 ,csa_tree_add_51_79_groupi_n_9977 ,csa_tree_add_51_79_groupi_n_10076);
  xnor csa_tree_add_51_79_groupi_g35835__8246(csa_tree_add_51_79_groupi_n_10282 ,csa_tree_add_51_79_groupi_n_9931 ,csa_tree_add_51_79_groupi_n_9956);
  xnor csa_tree_add_51_79_groupi_g35836__7098(csa_tree_add_51_79_groupi_n_10281 ,csa_tree_add_51_79_groupi_n_9685 ,csa_tree_add_51_79_groupi_n_9949);
  xnor csa_tree_add_51_79_groupi_g35837__6131(csa_tree_add_51_79_groupi_n_10280 ,csa_tree_add_51_79_groupi_n_9994 ,csa_tree_add_51_79_groupi_n_9962);
  xnor csa_tree_add_51_79_groupi_g35838__1881(csa_tree_add_51_79_groupi_n_10279 ,csa_tree_add_51_79_groupi_n_9457 ,csa_tree_add_51_79_groupi_n_9951);
  xnor csa_tree_add_51_79_groupi_g35839__5115(csa_tree_add_51_79_groupi_n_10278 ,csa_tree_add_51_79_groupi_n_9871 ,csa_tree_add_51_79_groupi_n_9963);
  xnor csa_tree_add_51_79_groupi_g35840__7482(csa_tree_add_51_79_groupi_n_10277 ,csa_tree_add_51_79_groupi_n_9858 ,csa_tree_add_51_79_groupi_n_9961);
  xnor csa_tree_add_51_79_groupi_g35841__4733(csa_tree_add_51_79_groupi_n_10276 ,csa_tree_add_51_79_groupi_n_9680 ,csa_tree_add_51_79_groupi_n_9950);
  xnor csa_tree_add_51_79_groupi_g35842__6161(csa_tree_add_51_79_groupi_n_10275 ,csa_tree_add_51_79_groupi_n_9464 ,csa_tree_add_51_79_groupi_n_9948);
  xnor csa_tree_add_51_79_groupi_g35843__9315(csa_tree_add_51_79_groupi_n_10274 ,csa_tree_add_51_79_groupi_n_9945 ,csa_tree_add_51_79_groupi_n_9957);
  and csa_tree_add_51_79_groupi_g35844__9945(csa_tree_add_51_79_groupi_n_10273 ,csa_tree_add_51_79_groupi_n_9967 ,csa_tree_add_51_79_groupi_n_10120);
  xnor csa_tree_add_51_79_groupi_g35845__2883(csa_tree_add_51_79_groupi_n_10272 ,csa_tree_add_51_79_groupi_n_9934 ,csa_tree_add_51_79_groupi_n_9953);
  xnor csa_tree_add_51_79_groupi_g35846__2346(csa_tree_add_51_79_groupi_n_10271 ,csa_tree_add_51_79_groupi_n_9708 ,csa_tree_add_51_79_groupi_n_9955);
  xnor csa_tree_add_51_79_groupi_g35847__1666(csa_tree_add_51_79_groupi_n_10270 ,csa_tree_add_51_79_groupi_n_9913 ,csa_tree_add_51_79_groupi_n_9960);
  xnor csa_tree_add_51_79_groupi_g35848__7410(csa_tree_add_51_79_groupi_n_10268 ,csa_tree_add_51_79_groupi_n_8328 ,csa_tree_add_51_79_groupi_n_10078);
  xnor csa_tree_add_51_79_groupi_g35849__6417(csa_tree_add_51_79_groupi_n_10267 ,csa_tree_add_51_79_groupi_n_9706 ,csa_tree_add_51_79_groupi_n_9954);
  xnor csa_tree_add_51_79_groupi_g35850__5477(csa_tree_add_51_79_groupi_n_10266 ,csa_tree_add_51_79_groupi_n_9917 ,csa_tree_add_51_79_groupi_n_9952);
  xnor csa_tree_add_51_79_groupi_g35851__2398(csa_tree_add_51_79_groupi_n_10265 ,csa_tree_add_51_79_groupi_n_9362 ,csa_tree_add_51_79_groupi_n_9959);
  xnor csa_tree_add_51_79_groupi_g35852__5107(csa_tree_add_51_79_groupi_n_10264 ,csa_tree_add_51_79_groupi_n_9496 ,csa_tree_add_51_79_groupi_n_9958);
  or csa_tree_add_51_79_groupi_g35853__6260(csa_tree_add_51_79_groupi_n_10263 ,csa_tree_add_51_79_groupi_n_10042 ,csa_tree_add_51_79_groupi_n_10204);
  not csa_tree_add_51_79_groupi_g35854(csa_tree_add_51_79_groupi_n_10215 ,csa_tree_add_51_79_groupi_n_10216);
  or csa_tree_add_51_79_groupi_g35855__4319(csa_tree_add_51_79_groupi_n_10213 ,csa_tree_add_51_79_groupi_n_10063 ,csa_tree_add_51_79_groupi_n_9998);
  nor csa_tree_add_51_79_groupi_g35856__8428(csa_tree_add_51_79_groupi_n_10212 ,csa_tree_add_51_79_groupi_n_9679 ,csa_tree_add_51_79_groupi_n_10014);
  or csa_tree_add_51_79_groupi_g35857__5526(csa_tree_add_51_79_groupi_n_10211 ,csa_tree_add_51_79_groupi_n_9937 ,csa_tree_add_51_79_groupi_n_10057);
  and csa_tree_add_51_79_groupi_g35858__6783(csa_tree_add_51_79_groupi_n_10210 ,csa_tree_add_51_79_groupi_n_10058 ,csa_tree_add_51_79_groupi_n_10025);
  or csa_tree_add_51_79_groupi_g35859__3680(csa_tree_add_51_79_groupi_n_10209 ,csa_tree_add_51_79_groupi_n_9859 ,csa_tree_add_51_79_groupi_n_9985);
  or csa_tree_add_51_79_groupi_g35860__1617(csa_tree_add_51_79_groupi_n_10208 ,csa_tree_add_51_79_groupi_n_10056 ,csa_tree_add_51_79_groupi_n_10021);
  and csa_tree_add_51_79_groupi_g35861__2802(csa_tree_add_51_79_groupi_n_10207 ,csa_tree_add_51_79_groupi_n_9859 ,csa_tree_add_51_79_groupi_n_9985);
  and csa_tree_add_51_79_groupi_g35862__1705(csa_tree_add_51_79_groupi_n_10206 ,csa_tree_add_51_79_groupi_n_10072 ,csa_tree_add_51_79_groupi_n_9979);
  or csa_tree_add_51_79_groupi_g35863__5122(csa_tree_add_51_79_groupi_n_10205 ,csa_tree_add_51_79_groupi_n_10072 ,csa_tree_add_51_79_groupi_n_9979);
  nor csa_tree_add_51_79_groupi_g35864__8246(csa_tree_add_51_79_groupi_n_10204 ,csa_tree_add_51_79_groupi_n_9698 ,csa_tree_add_51_79_groupi_n_10040);
  nor csa_tree_add_51_79_groupi_g35865__7098(csa_tree_add_51_79_groupi_n_10203 ,csa_tree_add_51_79_groupi_n_9989 ,csa_tree_add_51_79_groupi_n_10010);
  or csa_tree_add_51_79_groupi_g35866__6131(csa_tree_add_51_79_groupi_n_10202 ,csa_tree_add_51_79_groupi_n_9942 ,csa_tree_add_51_79_groupi_n_10043);
  or csa_tree_add_51_79_groupi_g35867__1881(csa_tree_add_51_79_groupi_n_10201 ,csa_tree_add_51_79_groupi_n_9991 ,csa_tree_add_51_79_groupi_n_10064);
  and csa_tree_add_51_79_groupi_g35868__5115(csa_tree_add_51_79_groupi_n_10200 ,csa_tree_add_51_79_groupi_n_9991 ,csa_tree_add_51_79_groupi_n_10064);
  and csa_tree_add_51_79_groupi_g35869__7482(csa_tree_add_51_79_groupi_n_10199 ,csa_tree_add_51_79_groupi_n_9935 ,csa_tree_add_51_79_groupi_n_9983);
  or csa_tree_add_51_79_groupi_g35870__4733(csa_tree_add_51_79_groupi_n_10198 ,csa_tree_add_51_79_groupi_n_9935 ,csa_tree_add_51_79_groupi_n_9983);
  nor csa_tree_add_51_79_groupi_g35871__6161(csa_tree_add_51_79_groupi_n_10197 ,csa_tree_add_51_79_groupi_n_10069 ,csa_tree_add_51_79_groupi_n_10017);
  or csa_tree_add_51_79_groupi_g35872__9315(csa_tree_add_51_79_groupi_n_10196 ,csa_tree_add_51_79_groupi_n_10070 ,csa_tree_add_51_79_groupi_n_33);
  or csa_tree_add_51_79_groupi_g35873__9945(csa_tree_add_51_79_groupi_n_10195 ,csa_tree_add_51_79_groupi_n_9611 ,csa_tree_add_51_79_groupi_n_10039);
  or csa_tree_add_51_79_groupi_g35874__2883(csa_tree_add_51_79_groupi_n_10194 ,csa_tree_add_51_79_groupi_n_9988 ,csa_tree_add_51_79_groupi_n_10009);
  or csa_tree_add_51_79_groupi_g35875__2346(csa_tree_add_51_79_groupi_n_10193 ,csa_tree_add_51_79_groupi_n_9700 ,csa_tree_add_51_79_groupi_n_10037);
  or csa_tree_add_51_79_groupi_g35876__1666(csa_tree_add_51_79_groupi_n_10192 ,csa_tree_add_51_79_groupi_n_9701 ,csa_tree_add_51_79_groupi_n_10035);
  and csa_tree_add_51_79_groupi_g35877__7410(csa_tree_add_51_79_groupi_n_10191 ,csa_tree_add_51_79_groupi_n_10071 ,csa_tree_add_51_79_groupi_n_10074);
  or csa_tree_add_51_79_groupi_g35878__6417(csa_tree_add_51_79_groupi_n_10190 ,csa_tree_add_51_79_groupi_n_10071 ,csa_tree_add_51_79_groupi_n_10074);
  or csa_tree_add_51_79_groupi_g35879__5477(csa_tree_add_51_79_groupi_n_10189 ,csa_tree_add_51_79_groupi_n_9870 ,csa_tree_add_51_79_groupi_n_10033);
  or csa_tree_add_51_79_groupi_g35880__2398(csa_tree_add_51_79_groupi_n_10188 ,csa_tree_add_51_79_groupi_n_9922 ,csa_tree_add_51_79_groupi_n_10011);
  or csa_tree_add_51_79_groupi_g35881__5107(csa_tree_add_51_79_groupi_n_10187 ,csa_tree_add_51_79_groupi_n_10060 ,csa_tree_add_51_79_groupi_n_10001);
  and csa_tree_add_51_79_groupi_g35882__6260(csa_tree_add_51_79_groupi_n_10186 ,csa_tree_add_51_79_groupi_n_10060 ,csa_tree_add_51_79_groupi_n_10001);
  or csa_tree_add_51_79_groupi_g35883__4319(csa_tree_add_51_79_groupi_n_10185 ,csa_tree_add_51_79_groupi_n_9925 ,csa_tree_add_51_79_groupi_n_10000);
  and csa_tree_add_51_79_groupi_g35884__8428(csa_tree_add_51_79_groupi_n_10184 ,csa_tree_add_51_79_groupi_n_9925 ,csa_tree_add_51_79_groupi_n_10000);
  and csa_tree_add_51_79_groupi_g35885__5526(csa_tree_add_51_79_groupi_n_10183 ,csa_tree_add_51_79_groupi_n_9969 ,csa_tree_add_51_79_groupi_n_10087);
  and csa_tree_add_51_79_groupi_g35886__6783(csa_tree_add_51_79_groupi_n_10182 ,csa_tree_add_51_79_groupi_n_10063 ,csa_tree_add_51_79_groupi_n_9998);
  or csa_tree_add_51_79_groupi_g35887__3680(csa_tree_add_51_79_groupi_n_10181 ,csa_tree_add_51_79_groupi_n_9938 ,csa_tree_add_51_79_groupi_n_10029);
  and csa_tree_add_51_79_groupi_g35888__1617(csa_tree_add_51_79_groupi_n_10180 ,csa_tree_add_51_79_groupi_n_9922 ,csa_tree_add_51_79_groupi_n_10011);
  or csa_tree_add_51_79_groupi_g35889__2802(csa_tree_add_51_79_groupi_n_10179 ,csa_tree_add_51_79_groupi_n_9601 ,csa_tree_add_51_79_groupi_n_9975);
  and csa_tree_add_51_79_groupi_g35890__1705(csa_tree_add_51_79_groupi_n_10178 ,csa_tree_add_51_79_groupi_n_10076 ,csa_tree_add_51_79_groupi_n_9977);
  or csa_tree_add_51_79_groupi_g35891__5122(csa_tree_add_51_79_groupi_n_10177 ,csa_tree_add_51_79_groupi_n_10076 ,csa_tree_add_51_79_groupi_n_9977);
  or csa_tree_add_51_79_groupi_g35892__8246(csa_tree_add_51_79_groupi_n_10176 ,csa_tree_add_51_79_groupi_n_9704 ,csa_tree_add_51_79_groupi_n_10027);
  or csa_tree_add_51_79_groupi_g35893__7098(csa_tree_add_51_79_groupi_n_10175 ,csa_tree_add_51_79_groupi_n_9943 ,csa_tree_add_51_79_groupi_n_10031);
  or csa_tree_add_51_79_groupi_g35894__6131(csa_tree_add_51_79_groupi_n_10174 ,csa_tree_add_51_79_groupi_n_9861 ,csa_tree_add_51_79_groupi_n_10006);
  and csa_tree_add_51_79_groupi_g35895__1881(csa_tree_add_51_79_groupi_n_10173 ,csa_tree_add_51_79_groupi_n_9861 ,csa_tree_add_51_79_groupi_n_10006);
  or csa_tree_add_51_79_groupi_g35896__5115(csa_tree_add_51_79_groupi_n_10172 ,csa_tree_add_51_79_groupi_n_9936 ,csa_tree_add_51_79_groupi_n_10054);
  or csa_tree_add_51_79_groupi_g35897__7482(csa_tree_add_51_79_groupi_n_10171 ,csa_tree_add_51_79_groupi_n_9677 ,csa_tree_add_51_79_groupi_n_9994);
  and csa_tree_add_51_79_groupi_g35898__4733(csa_tree_add_51_79_groupi_n_10170 ,csa_tree_add_51_79_groupi_n_9677 ,csa_tree_add_51_79_groupi_n_9994);
  or csa_tree_add_51_79_groupi_g35899__6161(csa_tree_add_51_79_groupi_n_10169 ,csa_tree_add_51_79_groupi_n_9873 ,csa_tree_add_51_79_groupi_n_9973);
  or csa_tree_add_51_79_groupi_g35900__9315(csa_tree_add_51_79_groupi_n_10168 ,csa_tree_add_51_79_groupi_n_10080 ,csa_tree_add_51_79_groupi_n_10047);
  or csa_tree_add_51_79_groupi_g35901__9945(csa_tree_add_51_79_groupi_n_10167 ,csa_tree_add_51_79_groupi_n_9842 ,csa_tree_add_51_79_groupi_n_10023);
  and csa_tree_add_51_79_groupi_g35902__2883(csa_tree_add_51_79_groupi_n_10166 ,csa_tree_add_51_79_groupi_n_9990 ,csa_tree_add_51_79_groupi_n_10012);
  or csa_tree_add_51_79_groupi_g35903__2346(csa_tree_add_51_79_groupi_n_10165 ,csa_tree_add_51_79_groupi_n_9990 ,csa_tree_add_51_79_groupi_n_10012);
  or csa_tree_add_51_79_groupi_g35904__1666(csa_tree_add_51_79_groupi_n_10164 ,csa_tree_add_51_79_groupi_n_8329 ,csa_tree_add_51_79_groupi_n_10078);
  and csa_tree_add_51_79_groupi_g35905__7410(csa_tree_add_51_79_groupi_n_10224 ,csa_tree_add_51_79_groupi_n_9848 ,csa_tree_add_51_79_groupi_n_9972);
  and csa_tree_add_51_79_groupi_g35906__6417(csa_tree_add_51_79_groupi_n_10223 ,csa_tree_add_51_79_groupi_n_9888 ,csa_tree_add_51_79_groupi_n_10028);
  and csa_tree_add_51_79_groupi_g35907__5477(csa_tree_add_51_79_groupi_n_10222 ,csa_tree_add_51_79_groupi_n_9905 ,csa_tree_add_51_79_groupi_n_10059);
  and csa_tree_add_51_79_groupi_g35908__2398(csa_tree_add_51_79_groupi_n_10221 ,csa_tree_add_51_79_groupi_n_9837 ,csa_tree_add_51_79_groupi_n_9970);
  and csa_tree_add_51_79_groupi_g35909__5107(csa_tree_add_51_79_groupi_n_10220 ,csa_tree_add_51_79_groupi_n_9846 ,csa_tree_add_51_79_groupi_n_9971);
  and csa_tree_add_51_79_groupi_g35910__6260(csa_tree_add_51_79_groupi_n_10219 ,csa_tree_add_51_79_groupi_n_9900 ,csa_tree_add_51_79_groupi_n_10053);
  and csa_tree_add_51_79_groupi_g35911__4319(csa_tree_add_51_79_groupi_n_10218 ,csa_tree_add_51_79_groupi_n_9891 ,csa_tree_add_51_79_groupi_n_10049);
  and csa_tree_add_51_79_groupi_g35912__8428(csa_tree_add_51_79_groupi_n_10217 ,csa_tree_add_51_79_groupi_n_9880 ,csa_tree_add_51_79_groupi_n_10055);
  or csa_tree_add_51_79_groupi_g35913__5526(csa_tree_add_51_79_groupi_n_10216 ,csa_tree_add_51_79_groupi_n_9840 ,csa_tree_add_51_79_groupi_n_10046);
  and csa_tree_add_51_79_groupi_g35914__6783(csa_tree_add_51_79_groupi_n_10214 ,csa_tree_add_51_79_groupi_n_9729 ,csa_tree_add_51_79_groupi_n_10032);
  not csa_tree_add_51_79_groupi_g35915(csa_tree_add_51_79_groupi_n_10160 ,csa_tree_add_51_79_groupi_n_10159);
  not csa_tree_add_51_79_groupi_g35916(csa_tree_add_51_79_groupi_n_10158 ,csa_tree_add_51_79_groupi_n_10157);
  not csa_tree_add_51_79_groupi_g35917(csa_tree_add_51_79_groupi_n_10154 ,csa_tree_add_51_79_groupi_n_10153);
  not csa_tree_add_51_79_groupi_g35918(csa_tree_add_51_79_groupi_n_10151 ,csa_tree_add_51_79_groupi_n_10150);
  not csa_tree_add_51_79_groupi_g35919(csa_tree_add_51_79_groupi_n_10139 ,csa_tree_add_51_79_groupi_n_10138);
  not csa_tree_add_51_79_groupi_g35920(csa_tree_add_51_79_groupi_n_10137 ,csa_tree_add_51_79_groupi_n_10136);
  not csa_tree_add_51_79_groupi_g35921(csa_tree_add_51_79_groupi_n_10128 ,csa_tree_add_51_79_groupi_n_10129);
  nor csa_tree_add_51_79_groupi_g35922__3680(csa_tree_add_51_79_groupi_n_10126 ,csa_tree_add_51_79_groupi_n_10008 ,csa_tree_add_51_79_groupi_n_10003);
  or csa_tree_add_51_79_groupi_g35923__1617(csa_tree_add_51_79_groupi_n_10125 ,csa_tree_add_51_79_groupi_n_10007 ,csa_tree_add_51_79_groupi_n_10004);
  or csa_tree_add_51_79_groupi_g35924__2802(csa_tree_add_51_79_groupi_n_10124 ,csa_tree_add_51_79_groupi_n_10061 ,csa_tree_add_51_79_groupi_n_9993);
  and csa_tree_add_51_79_groupi_g35925__1705(csa_tree_add_51_79_groupi_n_10123 ,csa_tree_add_51_79_groupi_n_9997 ,csa_tree_add_51_79_groupi_n_9996);
  nor csa_tree_add_51_79_groupi_g35926__5122(csa_tree_add_51_79_groupi_n_10122 ,csa_tree_add_51_79_groupi_n_10062 ,csa_tree_add_51_79_groupi_n_9992);
  nor csa_tree_add_51_79_groupi_g35927__8246(csa_tree_add_51_79_groupi_n_10121 ,csa_tree_add_51_79_groupi_n_9997 ,csa_tree_add_51_79_groupi_n_9996);
  or csa_tree_add_51_79_groupi_g35928__7098(csa_tree_add_51_79_groupi_n_10120 ,csa_tree_add_51_79_groupi_n_9939 ,csa_tree_add_51_79_groupi_n_9966);
  or csa_tree_add_51_79_groupi_g35929__6131(csa_tree_add_51_79_groupi_n_10119 ,csa_tree_add_51_79_groupi_n_9854 ,csa_tree_add_51_79_groupi_n_9987);
  nor csa_tree_add_51_79_groupi_g35930__1881(csa_tree_add_51_79_groupi_n_10118 ,csa_tree_add_51_79_groupi_n_9855 ,csa_tree_add_51_79_groupi_n_9986);
  and csa_tree_add_51_79_groupi_g35931__5115(csa_tree_add_51_79_groupi_n_10117 ,csa_tree_add_51_79_groupi_n_9856 ,csa_tree_add_51_79_groupi_n_9984);
  or csa_tree_add_51_79_groupi_g35932__7482(csa_tree_add_51_79_groupi_n_10116 ,csa_tree_add_51_79_groupi_n_9856 ,csa_tree_add_51_79_groupi_n_9984);
  or csa_tree_add_51_79_groupi_g35933__4733(csa_tree_add_51_79_groupi_n_10115 ,csa_tree_add_51_79_groupi_n_10066 ,csa_tree_add_51_79_groupi_n_9980);
  nor csa_tree_add_51_79_groupi_g35934__6161(csa_tree_add_51_79_groupi_n_10114 ,csa_tree_add_51_79_groupi_n_10065 ,csa_tree_add_51_79_groupi_n_9981);
  or csa_tree_add_51_79_groupi_g35935__9315(csa_tree_add_51_79_groupi_n_10113 ,csa_tree_add_51_79_groupi_n_9678 ,csa_tree_add_51_79_groupi_n_10013);
  xnor csa_tree_add_51_79_groupi_g35936__9945(csa_tree_add_51_79_groupi_n_10112 ,csa_tree_add_51_79_groupi_n_9453 ,csa_tree_add_51_79_groupi_n_9929);
  xnor csa_tree_add_51_79_groupi_g35937__2883(csa_tree_add_51_79_groupi_n_10111 ,csa_tree_add_51_79_groupi_n_9799 ,csa_tree_add_51_79_groupi_n_9915);
  xnor csa_tree_add_51_79_groupi_g35938__2346(csa_tree_add_51_79_groupi_n_10110 ,csa_tree_add_51_79_groupi_n_9918 ,csa_tree_add_51_79_groupi_n_9789);
  xnor csa_tree_add_51_79_groupi_g35939__1666(csa_tree_add_51_79_groupi_n_10109 ,csa_tree_add_51_79_groupi_n_9788 ,csa_tree_add_51_79_groupi_n_9944);
  xnor csa_tree_add_51_79_groupi_g35940__7410(csa_tree_add_51_79_groupi_n_10108 ,csa_tree_add_51_79_groupi_n_9860 ,csa_tree_add_51_79_groupi_n_9923);
  xnor csa_tree_add_51_79_groupi_g35941__6417(csa_tree_add_51_79_groupi_n_10107 ,csa_tree_add_51_79_groupi_n_9947 ,csa_tree_add_51_79_groupi_n_9859);
  xnor csa_tree_add_51_79_groupi_g35942__5477(csa_tree_add_51_79_groupi_n_10106 ,csa_tree_add_51_79_groupi_n_9919 ,csa_tree_add_51_79_groupi_n_9924);
  xnor csa_tree_add_51_79_groupi_g35943__2398(csa_tree_add_51_79_groupi_n_10105 ,csa_tree_add_51_79_groupi_n_9933 ,csa_tree_add_51_79_groupi_n_9921);
  xnor csa_tree_add_51_79_groupi_g35944__5107(csa_tree_add_51_79_groupi_n_10104 ,csa_tree_add_51_79_groupi_n_9927 ,csa_tree_add_51_79_groupi_n_9868);
  xnor csa_tree_add_51_79_groupi_g35945__6260(csa_tree_add_51_79_groupi_n_10103 ,csa_tree_add_51_79_groupi_n_9692 ,csa_tree_add_51_79_groupi_n_9857);
  xnor csa_tree_add_51_79_groupi_g35946__4319(csa_tree_add_51_79_groupi_n_10102 ,csa_tree_add_51_79_groupi_n_9863 ,csa_tree_add_51_79_groupi_n_9686);
  xnor csa_tree_add_51_79_groupi_g35947__8428(csa_tree_add_51_79_groupi_n_10101 ,csa_tree_add_51_79_groupi_n_9943 ,csa_tree_add_51_79_groupi_n_8765);
  xnor csa_tree_add_51_79_groupi_g35948__5526(csa_tree_add_51_79_groupi_n_10100 ,csa_tree_add_51_79_groupi_n_9940 ,csa_tree_add_51_79_groupi_n_9856);
  xnor csa_tree_add_51_79_groupi_g35949__6783(csa_tree_add_51_79_groupi_n_10099 ,csa_tree_add_51_79_groupi_n_9853 ,csa_tree_add_51_79_groupi_n_9601);
  xnor csa_tree_add_51_79_groupi_g35950__3680(csa_tree_add_51_79_groupi_n_10098 ,csa_tree_add_51_79_groupi_n_9865 ,csa_tree_add_51_79_groupi_n_9938);
  xnor csa_tree_add_51_79_groupi_g35951__1617(csa_tree_add_51_79_groupi_n_10097 ,csa_tree_add_51_79_groupi_n_9916 ,csa_tree_add_51_79_groupi_n_9455);
  xnor csa_tree_add_51_79_groupi_g35952__2802(csa_tree_add_51_79_groupi_n_10163 ,csa_tree_add_51_79_groupi_n_9614 ,csa_tree_add_51_79_groupi_n_9821);
  xnor csa_tree_add_51_79_groupi_g35953__1705(csa_tree_add_51_79_groupi_n_10162 ,csa_tree_add_51_79_groupi_n_9695 ,csa_tree_add_51_79_groupi_n_9830);
  xnor csa_tree_add_51_79_groupi_g35954__5122(csa_tree_add_51_79_groupi_n_10161 ,csa_tree_add_51_79_groupi_n_9500 ,csa_tree_add_51_79_groupi_n_9834);
  xnor csa_tree_add_51_79_groupi_g35955__8246(csa_tree_add_51_79_groupi_n_10159 ,csa_tree_add_51_79_groupi_n_9705 ,csa_tree_add_51_79_groupi_n_9828);
  xnor csa_tree_add_51_79_groupi_g35956__7098(csa_tree_add_51_79_groupi_n_10157 ,csa_tree_add_51_79_groupi_n_9587 ,csa_tree_add_51_79_groupi_n_9833);
  xnor csa_tree_add_51_79_groupi_g35957__6131(csa_tree_add_51_79_groupi_n_10156 ,csa_tree_add_51_79_groupi_n_9466 ,csa_tree_add_51_79_groupi_n_9827);
  xnor csa_tree_add_51_79_groupi_g35958__1881(csa_tree_add_51_79_groupi_n_10155 ,csa_tree_add_51_79_groupi_n_9508 ,csa_tree_add_51_79_groupi_n_9826);
  xnor csa_tree_add_51_79_groupi_g35959__5115(csa_tree_add_51_79_groupi_n_10153 ,csa_tree_add_51_79_groupi_n_9805 ,csa_tree_add_51_79_groupi_n_9832);
  xnor csa_tree_add_51_79_groupi_g35960__7482(csa_tree_add_51_79_groupi_n_10152 ,csa_tree_add_51_79_groupi_n_9586 ,csa_tree_add_51_79_groupi_n_9807);
  xnor csa_tree_add_51_79_groupi_g35961__4733(csa_tree_add_51_79_groupi_n_10150 ,csa_tree_add_51_79_groupi_n_9402 ,csa_tree_add_51_79_groupi_n_9825);
  xnor csa_tree_add_51_79_groupi_g35962__6161(csa_tree_add_51_79_groupi_n_10149 ,csa_tree_add_51_79_groupi_n_9696 ,csa_tree_add_51_79_groupi_n_9831);
  xnor csa_tree_add_51_79_groupi_g35963__9315(csa_tree_add_51_79_groupi_n_10148 ,csa_tree_add_51_79_groupi_n_9451 ,csa_tree_add_51_79_groupi_n_9824);
  xnor csa_tree_add_51_79_groupi_g35964__9945(csa_tree_add_51_79_groupi_n_10147 ,csa_tree_add_51_79_groupi_n_9505 ,csa_tree_add_51_79_groupi_n_9823);
  xnor csa_tree_add_51_79_groupi_g35965__2883(csa_tree_add_51_79_groupi_n_10146 ,csa_tree_add_51_79_groupi_n_9699 ,csa_tree_add_51_79_groupi_n_9822);
  xnor csa_tree_add_51_79_groupi_g35966__2346(csa_tree_add_51_79_groupi_n_10145 ,csa_tree_add_51_79_groupi_n_9872 ,csa_tree_add_51_79_groupi_n_9820);
  xnor csa_tree_add_51_79_groupi_g35967__1666(csa_tree_add_51_79_groupi_n_10144 ,csa_tree_add_51_79_groupi_n_9482 ,csa_tree_add_51_79_groupi_n_9817);
  xnor csa_tree_add_51_79_groupi_g35968__7410(csa_tree_add_51_79_groupi_n_10143 ,csa_tree_add_51_79_groupi_n_9697 ,csa_tree_add_51_79_groupi_n_9829);
  xnor csa_tree_add_51_79_groupi_g35969__6417(csa_tree_add_51_79_groupi_n_10142 ,csa_tree_add_51_79_groupi_n_9602 ,csa_tree_add_51_79_groupi_n_9816);
  xnor csa_tree_add_51_79_groupi_g35970__5477(csa_tree_add_51_79_groupi_n_10141 ,csa_tree_add_51_79_groupi_n_9481 ,csa_tree_add_51_79_groupi_n_9819);
  xnor csa_tree_add_51_79_groupi_g35971__2398(csa_tree_add_51_79_groupi_n_10140 ,csa_tree_add_51_79_groupi_n_9606 ,csa_tree_add_51_79_groupi_n_9818);
  xnor csa_tree_add_51_79_groupi_g35972__5107(csa_tree_add_51_79_groupi_n_10138 ,csa_tree_add_51_79_groupi_n_9801 ,csa_tree_add_51_79_groupi_n_9812);
  xnor csa_tree_add_51_79_groupi_g35973__6260(csa_tree_add_51_79_groupi_n_10136 ,csa_tree_add_51_79_groupi_n_9439 ,csa_tree_add_51_79_groupi_n_9835);
  xnor csa_tree_add_51_79_groupi_g35974__4319(csa_tree_add_51_79_groupi_n_10135 ,csa_tree_add_51_79_groupi_n_9515 ,csa_tree_add_51_79_groupi_n_9814);
  xnor csa_tree_add_51_79_groupi_g35975__8428(csa_tree_add_51_79_groupi_n_10134 ,csa_tree_add_51_79_groupi_n_9688 ,csa_tree_add_51_79_groupi_n_9806);
  xnor csa_tree_add_51_79_groupi_g35976__5526(csa_tree_add_51_79_groupi_n_10133 ,csa_tree_add_51_79_groupi_n_9461 ,csa_tree_add_51_79_groupi_n_9813);
  xnor csa_tree_add_51_79_groupi_g35977__6783(csa_tree_add_51_79_groupi_n_10132 ,csa_tree_add_51_79_groupi_n_9604 ,csa_tree_add_51_79_groupi_n_9808);
  xnor csa_tree_add_51_79_groupi_g35978__3680(csa_tree_add_51_79_groupi_n_10131 ,csa_tree_add_51_79_groupi_n_9456 ,csa_tree_add_51_79_groupi_n_9811);
  xnor csa_tree_add_51_79_groupi_g35979__1617(csa_tree_add_51_79_groupi_n_10130 ,csa_tree_add_51_79_groupi_n_9702 ,csa_tree_add_51_79_groupi_n_9810);
  xnor csa_tree_add_51_79_groupi_g35980__2802(csa_tree_add_51_79_groupi_n_10129 ,csa_tree_add_51_79_groupi_n_9302 ,csa_tree_add_51_79_groupi_n_9815);
  xnor csa_tree_add_51_79_groupi_g35981__1705(csa_tree_add_51_79_groupi_n_10127 ,csa_tree_add_51_79_groupi_n_9612 ,csa_tree_add_51_79_groupi_n_9809);
  not csa_tree_add_51_79_groupi_g35982(csa_tree_add_51_79_groupi_n_10086 ,csa_tree_add_51_79_groupi_n_10085);
  not csa_tree_add_51_79_groupi_g35983(csa_tree_add_51_79_groupi_n_10069 ,csa_tree_add_51_79_groupi_n_10070);
  not csa_tree_add_51_79_groupi_g35984(csa_tree_add_51_79_groupi_n_10067 ,csa_tree_add_51_79_groupi_n_10068);
  not csa_tree_add_51_79_groupi_g35985(csa_tree_add_51_79_groupi_n_10065 ,csa_tree_add_51_79_groupi_n_10066);
  not csa_tree_add_51_79_groupi_g35986(csa_tree_add_51_79_groupi_n_10062 ,csa_tree_add_51_79_groupi_n_10061);
  or csa_tree_add_51_79_groupi_g35987__5122(csa_tree_add_51_79_groupi_n_10059 ,csa_tree_add_51_79_groupi_n_9946 ,csa_tree_add_51_79_groupi_n_9901);
  or csa_tree_add_51_79_groupi_g35988__8246(csa_tree_add_51_79_groupi_n_10058 ,csa_tree_add_51_79_groupi_n_9933 ,csa_tree_add_51_79_groupi_n_9920);
  and csa_tree_add_51_79_groupi_g35989__7098(csa_tree_add_51_79_groupi_n_10057 ,csa_tree_add_51_79_groupi_n_9923 ,csa_tree_add_51_79_groupi_n_9860);
  and csa_tree_add_51_79_groupi_g35990__6131(csa_tree_add_51_79_groupi_n_10056 ,csa_tree_add_51_79_groupi_n_9924 ,csa_tree_add_51_79_groupi_n_9919);
  or csa_tree_add_51_79_groupi_g35991__1881(csa_tree_add_51_79_groupi_n_10055 ,csa_tree_add_51_79_groupi_n_9800 ,csa_tree_add_51_79_groupi_n_9881);
  and csa_tree_add_51_79_groupi_g35992__5115(csa_tree_add_51_79_groupi_n_10054 ,csa_tree_add_51_79_groupi_n_9789 ,csa_tree_add_51_79_groupi_n_9918);
  or csa_tree_add_51_79_groupi_g35993__7482(csa_tree_add_51_79_groupi_n_10053 ,csa_tree_add_51_79_groupi_n_9709 ,csa_tree_add_51_79_groupi_n_9894);
  or csa_tree_add_51_79_groupi_g35994__4733(csa_tree_add_51_79_groupi_n_10052 ,csa_tree_add_51_79_groupi_n_9789 ,csa_tree_add_51_79_groupi_n_9918);
  or csa_tree_add_51_79_groupi_g35995__6161(csa_tree_add_51_79_groupi_n_10051 ,csa_tree_add_51_79_groupi_n_9452 ,csa_tree_add_51_79_groupi_n_9929);
  or csa_tree_add_51_79_groupi_g35996(csa_tree_add_51_79_groupi_n_10050 ,csa_tree_add_51_79_groupi_n_9924 ,csa_tree_add_51_79_groupi_n_9919);
  or csa_tree_add_51_79_groupi_g35997(csa_tree_add_51_79_groupi_n_10049 ,csa_tree_add_51_79_groupi_n_9871 ,csa_tree_add_51_79_groupi_n_9886);
  or csa_tree_add_51_79_groupi_g35998(csa_tree_add_51_79_groupi_n_10048 ,csa_tree_add_51_79_groupi_n_9686 ,csa_tree_add_51_79_groupi_n_9863);
  and csa_tree_add_51_79_groupi_g35999(csa_tree_add_51_79_groupi_n_10047 ,csa_tree_add_51_79_groupi_n_9686 ,csa_tree_add_51_79_groupi_n_9863);
  and csa_tree_add_51_79_groupi_g36000(csa_tree_add_51_79_groupi_n_10046 ,csa_tree_add_51_79_groupi_n_9944 ,csa_tree_add_51_79_groupi_n_9841);
  or csa_tree_add_51_79_groupi_g36001(csa_tree_add_51_79_groupi_n_10045 ,csa_tree_add_51_79_groupi_n_9689 ,csa_tree_add_51_79_groupi_n_9913);
  or csa_tree_add_51_79_groupi_g36002(csa_tree_add_51_79_groupi_n_10044 ,csa_tree_add_51_79_groupi_n_8765 ,csa_tree_add_51_79_groupi_n_31);
  nor csa_tree_add_51_79_groupi_g36003(csa_tree_add_51_79_groupi_n_10043 ,csa_tree_add_51_79_groupi_n_9453 ,csa_tree_add_51_79_groupi_n_9928);
  nor csa_tree_add_51_79_groupi_g36004(csa_tree_add_51_79_groupi_n_10042 ,csa_tree_add_51_79_groupi_n_9934 ,csa_tree_add_51_79_groupi_n_9674);
  nor csa_tree_add_51_79_groupi_g36005(csa_tree_add_51_79_groupi_n_10041 ,csa_tree_add_51_79_groupi_n_9932 ,csa_tree_add_51_79_groupi_n_9921);
  and csa_tree_add_51_79_groupi_g36006(csa_tree_add_51_79_groupi_n_10040 ,csa_tree_add_51_79_groupi_n_9934 ,csa_tree_add_51_79_groupi_n_9674);
  and csa_tree_add_51_79_groupi_g36007(csa_tree_add_51_79_groupi_n_10039 ,csa_tree_add_51_79_groupi_n_9689 ,csa_tree_add_51_79_groupi_n_9913);
  or csa_tree_add_51_79_groupi_g36008(csa_tree_add_51_79_groupi_n_10038 ,csa_tree_add_51_79_groupi_n_9684 ,csa_tree_add_51_79_groupi_n_9858);
  and csa_tree_add_51_79_groupi_g36009(csa_tree_add_51_79_groupi_n_10037 ,csa_tree_add_51_79_groupi_n_9684 ,csa_tree_add_51_79_groupi_n_9858);
  or csa_tree_add_51_79_groupi_g36010(csa_tree_add_51_79_groupi_n_10036 ,csa_tree_add_51_79_groupi_n_9917 ,csa_tree_add_51_79_groupi_n_9693);
  and csa_tree_add_51_79_groupi_g36011(csa_tree_add_51_79_groupi_n_10035 ,csa_tree_add_51_79_groupi_n_9917 ,csa_tree_add_51_79_groupi_n_9693);
  or csa_tree_add_51_79_groupi_g36012(csa_tree_add_51_79_groupi_n_10034 ,csa_tree_add_51_79_groupi_n_9455 ,csa_tree_add_51_79_groupi_n_9916);
  and csa_tree_add_51_79_groupi_g36013(csa_tree_add_51_79_groupi_n_10033 ,csa_tree_add_51_79_groupi_n_9455 ,csa_tree_add_51_79_groupi_n_9916);
  or csa_tree_add_51_79_groupi_g36014(csa_tree_add_51_79_groupi_n_10032 ,csa_tree_add_51_79_groupi_n_9872 ,csa_tree_add_51_79_groupi_n_9728);
  and csa_tree_add_51_79_groupi_g36015(csa_tree_add_51_79_groupi_n_10031 ,csa_tree_add_51_79_groupi_n_8765 ,csa_tree_add_51_79_groupi_n_31);
  or csa_tree_add_51_79_groupi_g36016(csa_tree_add_51_79_groupi_n_10030 ,csa_tree_add_51_79_groupi_n_9865 ,csa_tree_add_51_79_groupi_n_9930);
  and csa_tree_add_51_79_groupi_g36017(csa_tree_add_51_79_groupi_n_10029 ,csa_tree_add_51_79_groupi_n_9865 ,csa_tree_add_51_79_groupi_n_9930);
  or csa_tree_add_51_79_groupi_g36018(csa_tree_add_51_79_groupi_n_10028 ,csa_tree_add_51_79_groupi_n_9706 ,csa_tree_add_51_79_groupi_n_9889);
  and csa_tree_add_51_79_groupi_g36019(csa_tree_add_51_79_groupi_n_10027 ,csa_tree_add_51_79_groupi_n_9589 ,csa_tree_add_51_79_groupi_n_9931);
  or csa_tree_add_51_79_groupi_g36020(csa_tree_add_51_79_groupi_n_10026 ,csa_tree_add_51_79_groupi_n_9589 ,csa_tree_add_51_79_groupi_n_9931);
  and csa_tree_add_51_79_groupi_g36021(csa_tree_add_51_79_groupi_n_10096 ,csa_tree_add_51_79_groupi_n_9785 ,csa_tree_add_51_79_groupi_n_9911);
  and csa_tree_add_51_79_groupi_g36022(csa_tree_add_51_79_groupi_n_10095 ,csa_tree_add_51_79_groupi_n_9740 ,csa_tree_add_51_79_groupi_n_9877);
  and csa_tree_add_51_79_groupi_g36023(csa_tree_add_51_79_groupi_n_10094 ,csa_tree_add_51_79_groupi_n_9751 ,csa_tree_add_51_79_groupi_n_9912);
  and csa_tree_add_51_79_groupi_g36024(csa_tree_add_51_79_groupi_n_10093 ,csa_tree_add_51_79_groupi_n_9731 ,csa_tree_add_51_79_groupi_n_9879);
  and csa_tree_add_51_79_groupi_g36025(csa_tree_add_51_79_groupi_n_10092 ,csa_tree_add_51_79_groupi_n_9750 ,csa_tree_add_51_79_groupi_n_9882);
  and csa_tree_add_51_79_groupi_g36026(csa_tree_add_51_79_groupi_n_10091 ,csa_tree_add_51_79_groupi_n_9727 ,csa_tree_add_51_79_groupi_n_9884);
  and csa_tree_add_51_79_groupi_g36027(csa_tree_add_51_79_groupi_n_10090 ,csa_tree_add_51_79_groupi_n_9733 ,csa_tree_add_51_79_groupi_n_9910);
  or csa_tree_add_51_79_groupi_g36028(csa_tree_add_51_79_groupi_n_10089 ,csa_tree_add_51_79_groupi_n_9662 ,csa_tree_add_51_79_groupi_n_9899);
  and csa_tree_add_51_79_groupi_g36029(csa_tree_add_51_79_groupi_n_10088 ,csa_tree_add_51_79_groupi_n_9651 ,csa_tree_add_51_79_groupi_n_9875);
  or csa_tree_add_51_79_groupi_g36030(csa_tree_add_51_79_groupi_n_10087 ,csa_tree_add_51_79_groupi_n_9779 ,csa_tree_add_51_79_groupi_n_9907);
  or csa_tree_add_51_79_groupi_g36031(csa_tree_add_51_79_groupi_n_10085 ,csa_tree_add_51_79_groupi_n_9668 ,csa_tree_add_51_79_groupi_n_9878);
  and csa_tree_add_51_79_groupi_g36032(csa_tree_add_51_79_groupi_n_10084 ,csa_tree_add_51_79_groupi_n_9660 ,csa_tree_add_51_79_groupi_n_9885);
  and csa_tree_add_51_79_groupi_g36033(csa_tree_add_51_79_groupi_n_10083 ,csa_tree_add_51_79_groupi_n_9717 ,csa_tree_add_51_79_groupi_n_9896);
  and csa_tree_add_51_79_groupi_g36034(csa_tree_add_51_79_groupi_n_10082 ,csa_tree_add_51_79_groupi_n_9715 ,csa_tree_add_51_79_groupi_n_9897);
  and csa_tree_add_51_79_groupi_g36035(csa_tree_add_51_79_groupi_n_10081 ,csa_tree_add_51_79_groupi_n_9713 ,csa_tree_add_51_79_groupi_n_9902);
  and csa_tree_add_51_79_groupi_g36036(csa_tree_add_51_79_groupi_n_10080 ,csa_tree_add_51_79_groupi_n_9711 ,csa_tree_add_51_79_groupi_n_9903);
  and csa_tree_add_51_79_groupi_g36037(csa_tree_add_51_79_groupi_n_10079 ,csa_tree_add_51_79_groupi_n_9666 ,csa_tree_add_51_79_groupi_n_9904);
  and csa_tree_add_51_79_groupi_g36038(csa_tree_add_51_79_groupi_n_10078 ,csa_tree_add_51_79_groupi_n_8948 ,csa_tree_add_51_79_groupi_n_9906);
  and csa_tree_add_51_79_groupi_g36039(csa_tree_add_51_79_groupi_n_10077 ,csa_tree_add_51_79_groupi_n_9672 ,csa_tree_add_51_79_groupi_n_9908);
  and csa_tree_add_51_79_groupi_g36040(csa_tree_add_51_79_groupi_n_10076 ,csa_tree_add_51_79_groupi_n_9669 ,csa_tree_add_51_79_groupi_n_9909);
  and csa_tree_add_51_79_groupi_g36041(csa_tree_add_51_79_groupi_n_10075 ,csa_tree_add_51_79_groupi_n_9565 ,csa_tree_add_51_79_groupi_n_9893);
  and csa_tree_add_51_79_groupi_g36042(csa_tree_add_51_79_groupi_n_10074 ,csa_tree_add_51_79_groupi_n_9722 ,csa_tree_add_51_79_groupi_n_9890);
  and csa_tree_add_51_79_groupi_g36043(csa_tree_add_51_79_groupi_n_10073 ,csa_tree_add_51_79_groupi_n_9725 ,csa_tree_add_51_79_groupi_n_9887);
  and csa_tree_add_51_79_groupi_g36044(csa_tree_add_51_79_groupi_n_10072 ,csa_tree_add_51_79_groupi_n_9757 ,csa_tree_add_51_79_groupi_n_9851);
  and csa_tree_add_51_79_groupi_g36045(csa_tree_add_51_79_groupi_n_10071 ,csa_tree_add_51_79_groupi_n_9657 ,csa_tree_add_51_79_groupi_n_9852);
  and csa_tree_add_51_79_groupi_g36046(csa_tree_add_51_79_groupi_n_10070 ,csa_tree_add_51_79_groupi_n_9742 ,csa_tree_add_51_79_groupi_n_9874);
  or csa_tree_add_51_79_groupi_g36047(csa_tree_add_51_79_groupi_n_10068 ,csa_tree_add_51_79_groupi_n_9781 ,csa_tree_add_51_79_groupi_n_9850);
  and csa_tree_add_51_79_groupi_g36048(csa_tree_add_51_79_groupi_n_10066 ,csa_tree_add_51_79_groupi_n_9746 ,csa_tree_add_51_79_groupi_n_9876);
  and csa_tree_add_51_79_groupi_g36049(csa_tree_add_51_79_groupi_n_10064 ,csa_tree_add_51_79_groupi_n_9720 ,csa_tree_add_51_79_groupi_n_9883);
  and csa_tree_add_51_79_groupi_g36050(csa_tree_add_51_79_groupi_n_10063 ,csa_tree_add_51_79_groupi_n_9762 ,csa_tree_add_51_79_groupi_n_9892);
  or csa_tree_add_51_79_groupi_g36051(csa_tree_add_51_79_groupi_n_10061 ,csa_tree_add_51_79_groupi_n_9764 ,csa_tree_add_51_79_groupi_n_9895);
  and csa_tree_add_51_79_groupi_g36052(csa_tree_add_51_79_groupi_n_10060 ,csa_tree_add_51_79_groupi_n_9771 ,csa_tree_add_51_79_groupi_n_9898);
  not csa_tree_add_51_79_groupi_g36053(csa_tree_add_51_79_groupi_n_10020 ,csa_tree_add_51_79_groupi_n_10019);
  not csa_tree_add_51_79_groupi_g36054(csa_tree_add_51_79_groupi_n_10017 ,csa_tree_add_51_79_groupi_n_33);
  not csa_tree_add_51_79_groupi_g36055(csa_tree_add_51_79_groupi_n_10016 ,csa_tree_add_51_79_groupi_n_10015);
  not csa_tree_add_51_79_groupi_g36056(csa_tree_add_51_79_groupi_n_10014 ,csa_tree_add_51_79_groupi_n_10013);
  not csa_tree_add_51_79_groupi_g36057(csa_tree_add_51_79_groupi_n_10010 ,csa_tree_add_51_79_groupi_n_10009);
  not csa_tree_add_51_79_groupi_g36058(csa_tree_add_51_79_groupi_n_10008 ,csa_tree_add_51_79_groupi_n_10007);
  not csa_tree_add_51_79_groupi_g36059(csa_tree_add_51_79_groupi_n_10004 ,csa_tree_add_51_79_groupi_n_10003);
  not csa_tree_add_51_79_groupi_g36060(csa_tree_add_51_79_groupi_n_9996 ,csa_tree_add_51_79_groupi_n_9995);
  not csa_tree_add_51_79_groupi_g36061(csa_tree_add_51_79_groupi_n_9993 ,csa_tree_add_51_79_groupi_n_9992);
  not csa_tree_add_51_79_groupi_g36062(csa_tree_add_51_79_groupi_n_9988 ,csa_tree_add_51_79_groupi_n_9989);
  not csa_tree_add_51_79_groupi_g36063(csa_tree_add_51_79_groupi_n_9987 ,csa_tree_add_51_79_groupi_n_9986);
  not csa_tree_add_51_79_groupi_g36064(csa_tree_add_51_79_groupi_n_9981 ,csa_tree_add_51_79_groupi_n_9980);
  or csa_tree_add_51_79_groupi_g36065(csa_tree_add_51_79_groupi_n_9976 ,csa_tree_add_51_79_groupi_n_9853 ,csa_tree_add_51_79_groupi_n_9864);
  and csa_tree_add_51_79_groupi_g36066(csa_tree_add_51_79_groupi_n_9975 ,csa_tree_add_51_79_groupi_n_9853 ,csa_tree_add_51_79_groupi_n_9864);
  or csa_tree_add_51_79_groupi_g36067(csa_tree_add_51_79_groupi_n_9974 ,csa_tree_add_51_79_groupi_n_9857 ,csa_tree_add_51_79_groupi_n_9692);
  and csa_tree_add_51_79_groupi_g36068(csa_tree_add_51_79_groupi_n_9973 ,csa_tree_add_51_79_groupi_n_9857 ,csa_tree_add_51_79_groupi_n_9692);
  or csa_tree_add_51_79_groupi_g36069(csa_tree_add_51_79_groupi_n_9972 ,csa_tree_add_51_79_groupi_n_9516 ,csa_tree_add_51_79_groupi_n_9847);
  or csa_tree_add_51_79_groupi_g36070(csa_tree_add_51_79_groupi_n_9971 ,csa_tree_add_51_79_groupi_n_9703 ,csa_tree_add_51_79_groupi_n_9845);
  or csa_tree_add_51_79_groupi_g36071(csa_tree_add_51_79_groupi_n_9970 ,csa_tree_add_51_79_groupi_n_9598 ,csa_tree_add_51_79_groupi_n_9836);
  or csa_tree_add_51_79_groupi_g36072(csa_tree_add_51_79_groupi_n_9969 ,csa_tree_add_51_79_groupi_n_9798 ,csa_tree_add_51_79_groupi_n_9915);
  nor csa_tree_add_51_79_groupi_g36073(csa_tree_add_51_79_groupi_n_9968 ,csa_tree_add_51_79_groupi_n_9799 ,csa_tree_add_51_79_groupi_n_9914);
  or csa_tree_add_51_79_groupi_g36074(csa_tree_add_51_79_groupi_n_9967 ,csa_tree_add_51_79_groupi_n_9926 ,csa_tree_add_51_79_groupi_n_9867);
  nor csa_tree_add_51_79_groupi_g36075(csa_tree_add_51_79_groupi_n_9966 ,csa_tree_add_51_79_groupi_n_9927 ,csa_tree_add_51_79_groupi_n_9868);
  xnor csa_tree_add_51_79_groupi_g36076(out1[1] ,csa_tree_add_51_79_groupi_n_7592 ,csa_tree_add_51_79_groupi_n_9644);
  or csa_tree_add_51_79_groupi_g36077(csa_tree_add_51_79_groupi_n_9964 ,csa_tree_add_51_79_groupi_n_9923 ,csa_tree_add_51_79_groupi_n_9860);
  xnor csa_tree_add_51_79_groupi_g36078(csa_tree_add_51_79_groupi_n_9963 ,csa_tree_add_51_79_groupi_n_9681 ,csa_tree_add_51_79_groupi_n_9796);
  xnor csa_tree_add_51_79_groupi_g36079(csa_tree_add_51_79_groupi_n_9962 ,csa_tree_add_51_79_groupi_n_9677 ,csa_tree_add_51_79_groupi_n_9802);
  xnor csa_tree_add_51_79_groupi_g36080(csa_tree_add_51_79_groupi_n_9961 ,csa_tree_add_51_79_groupi_n_9700 ,csa_tree_add_51_79_groupi_n_9684);
  xnor csa_tree_add_51_79_groupi_g36081(csa_tree_add_51_79_groupi_n_9960 ,csa_tree_add_51_79_groupi_n_9689 ,csa_tree_add_51_79_groupi_n_9611);
  xnor csa_tree_add_51_79_groupi_g36082(csa_tree_add_51_79_groupi_n_9959 ,csa_tree_add_51_79_groupi_n_9803 ,csa_tree_add_51_79_groupi_n_9363);
  xnor csa_tree_add_51_79_groupi_g36083(csa_tree_add_51_79_groupi_n_9958 ,csa_tree_add_51_79_groupi_n_9516 ,csa_tree_add_51_79_groupi_n_9691);
  xnor csa_tree_add_51_79_groupi_g36084(csa_tree_add_51_79_groupi_n_9957 ,csa_tree_add_51_79_groupi_n_9683 ,csa_tree_add_51_79_groupi_n_9592);
  xor csa_tree_add_51_79_groupi_g36085(csa_tree_add_51_79_groupi_n_9956 ,csa_tree_add_51_79_groupi_n_9704 ,csa_tree_add_51_79_groupi_n_9589);
  xnor csa_tree_add_51_79_groupi_g36086(csa_tree_add_51_79_groupi_n_9955 ,csa_tree_add_51_79_groupi_n_9594 ,csa_tree_add_51_79_groupi_n_9791);
  xnor csa_tree_add_51_79_groupi_g36087(csa_tree_add_51_79_groupi_n_9954 ,csa_tree_add_51_79_groupi_n_9582 ,csa_tree_add_51_79_groupi_n_9797);
  xnor csa_tree_add_51_79_groupi_g36088(csa_tree_add_51_79_groupi_n_9953 ,csa_tree_add_51_79_groupi_n_9674 ,csa_tree_add_51_79_groupi_n_9698);
  xnor csa_tree_add_51_79_groupi_g36089(csa_tree_add_51_79_groupi_n_9952 ,csa_tree_add_51_79_groupi_n_9693 ,csa_tree_add_51_79_groupi_n_9701);
  xnor csa_tree_add_51_79_groupi_g36090(csa_tree_add_51_79_groupi_n_9951 ,csa_tree_add_51_79_groupi_n_9475 ,csa_tree_add_51_79_groupi_n_9694);
  xnor csa_tree_add_51_79_groupi_g36091(csa_tree_add_51_79_groupi_n_9950 ,csa_tree_add_51_79_groupi_n_9682 ,csa_tree_add_51_79_groupi_n_9800);
  xnor csa_tree_add_51_79_groupi_g36092(csa_tree_add_51_79_groupi_n_9949 ,csa_tree_add_51_79_groupi_n_9703 ,csa_tree_add_51_79_groupi_n_9690);
  xnor csa_tree_add_51_79_groupi_g36093(csa_tree_add_51_79_groupi_n_9948 ,csa_tree_add_51_79_groupi_n_9707 ,csa_tree_add_51_79_groupi_n_9465);
  or csa_tree_add_51_79_groupi_g36094(csa_tree_add_51_79_groupi_n_10025 ,csa_tree_add_51_79_groupi_n_9664 ,csa_tree_add_51_79_groupi_n_9839);
  and csa_tree_add_51_79_groupi_g36095(csa_tree_add_51_79_groupi_n_10024 ,csa_tree_add_51_79_groupi_n_9661 ,csa_tree_add_51_79_groupi_n_9849);
  xnor csa_tree_add_51_79_groupi_g36096(csa_tree_add_51_79_groupi_n_10023 ,csa_tree_add_51_79_groupi_n_9447 ,csa_tree_add_51_79_groupi_n_9641);
  xnor csa_tree_add_51_79_groupi_g36097(csa_tree_add_51_79_groupi_n_10022 ,csa_tree_add_51_79_groupi_n_9463 ,csa_tree_add_51_79_groupi_n_9632);
  xnor csa_tree_add_51_79_groupi_g36098(csa_tree_add_51_79_groupi_n_10021 ,csa_tree_add_51_79_groupi_n_9368 ,csa_tree_add_51_79_groupi_n_9633);
  or csa_tree_add_51_79_groupi_g36099(csa_tree_add_51_79_groupi_n_10019 ,csa_tree_add_51_79_groupi_n_9656 ,csa_tree_add_51_79_groupi_n_9838);
  xnor csa_tree_add_51_79_groupi_g36100(csa_tree_add_51_79_groupi_n_10018 ,csa_tree_add_51_79_groupi_n_9297 ,csa_tree_add_51_79_groupi_n_9620);
  xnor csa_tree_add_51_79_groupi_g36102(csa_tree_add_51_79_groupi_n_10015 ,csa_tree_add_51_79_groupi_n_9391 ,csa_tree_add_51_79_groupi_n_9624);
  xnor csa_tree_add_51_79_groupi_g36103(csa_tree_add_51_79_groupi_n_10013 ,csa_tree_add_51_79_groupi_n_9502 ,csa_tree_add_51_79_groupi_n_9640);
  xnor csa_tree_add_51_79_groupi_g36104(csa_tree_add_51_79_groupi_n_10012 ,csa_tree_add_51_79_groupi_n_9303 ,csa_tree_add_51_79_groupi_n_9629);
  xnor csa_tree_add_51_79_groupi_g36105(csa_tree_add_51_79_groupi_n_10011 ,csa_tree_add_51_79_groupi_n_9396 ,csa_tree_add_51_79_groupi_n_9622);
  xnor csa_tree_add_51_79_groupi_g36106(csa_tree_add_51_79_groupi_n_10009 ,csa_tree_add_51_79_groupi_n_9300 ,csa_tree_add_51_79_groupi_n_9621);
  xnor csa_tree_add_51_79_groupi_g36107(csa_tree_add_51_79_groupi_n_10007 ,csa_tree_add_51_79_groupi_n_9294 ,csa_tree_add_51_79_groupi_n_9639);
  xnor csa_tree_add_51_79_groupi_g36108(csa_tree_add_51_79_groupi_n_10006 ,csa_tree_add_51_79_groupi_n_9509 ,csa_tree_add_51_79_groupi_n_9619);
  xnor csa_tree_add_51_79_groupi_g36109(csa_tree_add_51_79_groupi_n_10005 ,csa_tree_add_51_79_groupi_n_9397 ,csa_tree_add_51_79_groupi_n_9618);
  xnor csa_tree_add_51_79_groupi_g36110(csa_tree_add_51_79_groupi_n_10003 ,csa_tree_add_51_79_groupi_n_9249 ,csa_tree_add_51_79_groupi_n_9638);
  xnor csa_tree_add_51_79_groupi_g36111(csa_tree_add_51_79_groupi_n_10002 ,csa_tree_add_51_79_groupi_n_9250 ,csa_tree_add_51_79_groupi_n_9617);
  xnor csa_tree_add_51_79_groupi_g36112(csa_tree_add_51_79_groupi_n_10001 ,csa_tree_add_51_79_groupi_n_9264 ,csa_tree_add_51_79_groupi_n_9615);
  xnor csa_tree_add_51_79_groupi_g36113(csa_tree_add_51_79_groupi_n_10000 ,csa_tree_add_51_79_groupi_n_9398 ,csa_tree_add_51_79_groupi_n_9616);
  xnor csa_tree_add_51_79_groupi_g36114(csa_tree_add_51_79_groupi_n_9999 ,csa_tree_add_51_79_groupi_n_9804 ,csa_tree_add_51_79_groupi_n_9000);
  xnor csa_tree_add_51_79_groupi_g36115(csa_tree_add_51_79_groupi_n_9998 ,csa_tree_add_51_79_groupi_n_9389 ,csa_tree_add_51_79_groupi_n_9623);
  xnor csa_tree_add_51_79_groupi_g36116(csa_tree_add_51_79_groupi_n_9997 ,csa_tree_add_51_79_groupi_n_9400 ,csa_tree_add_51_79_groupi_n_9636);
  xnor csa_tree_add_51_79_groupi_g36117(csa_tree_add_51_79_groupi_n_9995 ,csa_tree_add_51_79_groupi_n_9595 ,csa_tree_add_51_79_groupi_n_9634);
  xnor csa_tree_add_51_79_groupi_g36118(csa_tree_add_51_79_groupi_n_9994 ,csa_tree_add_51_79_groupi_n_9373 ,csa_tree_add_51_79_groupi_n_9625);
  xnor csa_tree_add_51_79_groupi_g36119(csa_tree_add_51_79_groupi_n_9992 ,csa_tree_add_51_79_groupi_n_9075 ,csa_tree_add_51_79_groupi_n_9635);
  xnor csa_tree_add_51_79_groupi_g36120(csa_tree_add_51_79_groupi_n_9991 ,csa_tree_add_51_79_groupi_n_9282 ,csa_tree_add_51_79_groupi_n_9637);
  and csa_tree_add_51_79_groupi_g36121(csa_tree_add_51_79_groupi_n_9990 ,csa_tree_add_51_79_groupi_n_9653 ,csa_tree_add_51_79_groupi_n_9844);
  xnor csa_tree_add_51_79_groupi_g36122(csa_tree_add_51_79_groupi_n_9989 ,csa_tree_add_51_79_groupi_n_9377 ,csa_tree_add_51_79_groupi_n_9643);
  xnor csa_tree_add_51_79_groupi_g36123(csa_tree_add_51_79_groupi_n_9986 ,csa_tree_add_51_79_groupi_n_9305 ,csa_tree_add_51_79_groupi_n_9631);
  xnor csa_tree_add_51_79_groupi_g36124(csa_tree_add_51_79_groupi_n_9985 ,csa_tree_add_51_79_groupi_n_9275 ,csa_tree_add_51_79_groupi_n_9648);
  xnor csa_tree_add_51_79_groupi_g36125(csa_tree_add_51_79_groupi_n_9984 ,csa_tree_add_51_79_groupi_n_9251 ,csa_tree_add_51_79_groupi_n_9630);
  xnor csa_tree_add_51_79_groupi_g36126(csa_tree_add_51_79_groupi_n_9983 ,csa_tree_add_51_79_groupi_n_9266 ,csa_tree_add_51_79_groupi_n_9647);
  xnor csa_tree_add_51_79_groupi_g36127(csa_tree_add_51_79_groupi_n_9982 ,csa_tree_add_51_79_groupi_n_9514 ,csa_tree_add_51_79_groupi_n_9626);
  xnor csa_tree_add_51_79_groupi_g36128(csa_tree_add_51_79_groupi_n_9980 ,csa_tree_add_51_79_groupi_n_9360 ,csa_tree_add_51_79_groupi_n_9628);
  xnor csa_tree_add_51_79_groupi_g36129(csa_tree_add_51_79_groupi_n_9979 ,csa_tree_add_51_79_groupi_n_9259 ,csa_tree_add_51_79_groupi_n_9642);
  xnor csa_tree_add_51_79_groupi_g36130(csa_tree_add_51_79_groupi_n_9978 ,csa_tree_add_51_79_groupi_n_9395 ,csa_tree_add_51_79_groupi_n_9645);
  xnor csa_tree_add_51_79_groupi_g36131(csa_tree_add_51_79_groupi_n_9977 ,csa_tree_add_51_79_groupi_n_9283 ,csa_tree_add_51_79_groupi_n_9627);
  not csa_tree_add_51_79_groupi_g36132(csa_tree_add_51_79_groupi_n_9946 ,csa_tree_add_51_79_groupi_n_9945);
  not csa_tree_add_51_79_groupi_g36133(csa_tree_add_51_79_groupi_n_9942 ,csa_tree_add_51_79_groupi_n_9941);
  not csa_tree_add_51_79_groupi_g36134(csa_tree_add_51_79_groupi_n_9933 ,csa_tree_add_51_79_groupi_n_9932);
  not csa_tree_add_51_79_groupi_g36135(csa_tree_add_51_79_groupi_n_9928 ,csa_tree_add_51_79_groupi_n_9929);
  not csa_tree_add_51_79_groupi_g36136(csa_tree_add_51_79_groupi_n_9927 ,csa_tree_add_51_79_groupi_n_9926);
  not csa_tree_add_51_79_groupi_g36137(csa_tree_add_51_79_groupi_n_9920 ,csa_tree_add_51_79_groupi_n_9921);
  not csa_tree_add_51_79_groupi_g36138(csa_tree_add_51_79_groupi_n_9915 ,csa_tree_add_51_79_groupi_n_9914);
  or csa_tree_add_51_79_groupi_g36139(csa_tree_add_51_79_groupi_n_9912 ,csa_tree_add_51_79_groupi_n_9613 ,csa_tree_add_51_79_groupi_n_9747);
  or csa_tree_add_51_79_groupi_g36140(csa_tree_add_51_79_groupi_n_9911 ,csa_tree_add_51_79_groupi_n_9596 ,csa_tree_add_51_79_groupi_n_9784);
  or csa_tree_add_51_79_groupi_g36141(csa_tree_add_51_79_groupi_n_9910 ,csa_tree_add_51_79_groupi_n_9197 ,csa_tree_add_51_79_groupi_n_9732);
  or csa_tree_add_51_79_groupi_g36142(csa_tree_add_51_79_groupi_n_9909 ,csa_tree_add_51_79_groupi_n_8968 ,csa_tree_add_51_79_groupi_n_9670);
  or csa_tree_add_51_79_groupi_g36143(csa_tree_add_51_79_groupi_n_9908 ,csa_tree_add_51_79_groupi_n_9386 ,csa_tree_add_51_79_groupi_n_9671);
  nor csa_tree_add_51_79_groupi_g36144(csa_tree_add_51_79_groupi_n_9907 ,csa_tree_add_51_79_groupi_n_9600 ,csa_tree_add_51_79_groupi_n_9778);
  or csa_tree_add_51_79_groupi_g36145(csa_tree_add_51_79_groupi_n_9906 ,csa_tree_add_51_79_groupi_n_8949 ,csa_tree_add_51_79_groupi_n_9804);
  or csa_tree_add_51_79_groupi_g36146(csa_tree_add_51_79_groupi_n_9905 ,csa_tree_add_51_79_groupi_n_9592 ,csa_tree_add_51_79_groupi_n_9683);
  or csa_tree_add_51_79_groupi_g36147(csa_tree_add_51_79_groupi_n_9904 ,csa_tree_add_51_79_groupi_n_9307 ,csa_tree_add_51_79_groupi_n_9665);
  or csa_tree_add_51_79_groupi_g36148(csa_tree_add_51_79_groupi_n_9903 ,csa_tree_add_51_79_groupi_n_9388 ,csa_tree_add_51_79_groupi_n_9710);
  or csa_tree_add_51_79_groupi_g36149(csa_tree_add_51_79_groupi_n_9902 ,csa_tree_add_51_79_groupi_n_9302 ,csa_tree_add_51_79_groupi_n_9712);
  and csa_tree_add_51_79_groupi_g36150(csa_tree_add_51_79_groupi_n_9901 ,csa_tree_add_51_79_groupi_n_9592 ,csa_tree_add_51_79_groupi_n_9683);
  or csa_tree_add_51_79_groupi_g36151(csa_tree_add_51_79_groupi_n_9900 ,csa_tree_add_51_79_groupi_n_9593 ,csa_tree_add_51_79_groupi_n_9791);
  and csa_tree_add_51_79_groupi_g36152(csa_tree_add_51_79_groupi_n_9899 ,csa_tree_add_51_79_groupi_n_9673 ,csa_tree_add_51_79_groupi_n_9695);
  or csa_tree_add_51_79_groupi_g36153(csa_tree_add_51_79_groupi_n_9898 ,csa_tree_add_51_79_groupi_n_9606 ,csa_tree_add_51_79_groupi_n_9769);
  or csa_tree_add_51_79_groupi_g36154(csa_tree_add_51_79_groupi_n_9897 ,csa_tree_add_51_79_groupi_n_9702 ,csa_tree_add_51_79_groupi_n_9714);
  or csa_tree_add_51_79_groupi_g36155(csa_tree_add_51_79_groupi_n_9896 ,csa_tree_add_51_79_groupi_n_9599 ,csa_tree_add_51_79_groupi_n_9716);
  nor csa_tree_add_51_79_groupi_g36156(csa_tree_add_51_79_groupi_n_9895 ,csa_tree_add_51_79_groupi_n_9607 ,csa_tree_add_51_79_groupi_n_9763);
  nor csa_tree_add_51_79_groupi_g36157(csa_tree_add_51_79_groupi_n_9894 ,csa_tree_add_51_79_groupi_n_9594 ,csa_tree_add_51_79_groupi_n_9790);
  or csa_tree_add_51_79_groupi_g36158(csa_tree_add_51_79_groupi_n_9893 ,csa_tree_add_51_79_groupi_n_9803 ,csa_tree_add_51_79_groupi_n_9569);
  or csa_tree_add_51_79_groupi_g36159(csa_tree_add_51_79_groupi_n_9892 ,csa_tree_add_51_79_groupi_n_9515 ,csa_tree_add_51_79_groupi_n_9761);
  or csa_tree_add_51_79_groupi_g36160(csa_tree_add_51_79_groupi_n_9891 ,csa_tree_add_51_79_groupi_n_9796 ,csa_tree_add_51_79_groupi_n_9681);
  or csa_tree_add_51_79_groupi_g36161(csa_tree_add_51_79_groupi_n_9890 ,csa_tree_add_51_79_groupi_n_9608 ,csa_tree_add_51_79_groupi_n_9721);
  and csa_tree_add_51_79_groupi_g36162(csa_tree_add_51_79_groupi_n_9889 ,csa_tree_add_51_79_groupi_n_9797 ,csa_tree_add_51_79_groupi_n_9582);
  or csa_tree_add_51_79_groupi_g36163(csa_tree_add_51_79_groupi_n_9888 ,csa_tree_add_51_79_groupi_n_9797 ,csa_tree_add_51_79_groupi_n_9582);
  or csa_tree_add_51_79_groupi_g36164(csa_tree_add_51_79_groupi_n_9887 ,csa_tree_add_51_79_groupi_n_9707 ,csa_tree_add_51_79_groupi_n_9724);
  and csa_tree_add_51_79_groupi_g36165(csa_tree_add_51_79_groupi_n_9886 ,csa_tree_add_51_79_groupi_n_9796 ,csa_tree_add_51_79_groupi_n_9681);
  or csa_tree_add_51_79_groupi_g36166(csa_tree_add_51_79_groupi_n_9885 ,csa_tree_add_51_79_groupi_n_9659 ,csa_tree_add_51_79_groupi_n_9699);
  or csa_tree_add_51_79_groupi_g36167(csa_tree_add_51_79_groupi_n_9884 ,csa_tree_add_51_79_groupi_n_9602 ,csa_tree_add_51_79_groupi_n_9726);
  or csa_tree_add_51_79_groupi_g36168(csa_tree_add_51_79_groupi_n_9883 ,csa_tree_add_51_79_groupi_n_9801 ,csa_tree_add_51_79_groupi_n_9719);
  or csa_tree_add_51_79_groupi_g36169(csa_tree_add_51_79_groupi_n_9882 ,csa_tree_add_51_79_groupi_n_9612 ,csa_tree_add_51_79_groupi_n_9749);
  and csa_tree_add_51_79_groupi_g36170(csa_tree_add_51_79_groupi_n_9881 ,csa_tree_add_51_79_groupi_n_9682 ,csa_tree_add_51_79_groupi_n_9680);
  or csa_tree_add_51_79_groupi_g36171(csa_tree_add_51_79_groupi_n_9880 ,csa_tree_add_51_79_groupi_n_9682 ,csa_tree_add_51_79_groupi_n_9680);
  or csa_tree_add_51_79_groupi_g36172(csa_tree_add_51_79_groupi_n_9879 ,csa_tree_add_51_79_groupi_n_9614 ,csa_tree_add_51_79_groupi_n_9730);
  and csa_tree_add_51_79_groupi_g36173(csa_tree_add_51_79_groupi_n_9878 ,csa_tree_add_51_79_groupi_n_9667 ,csa_tree_add_51_79_groupi_n_9697);
  or csa_tree_add_51_79_groupi_g36174(csa_tree_add_51_79_groupi_n_9877 ,csa_tree_add_51_79_groupi_n_9739 ,csa_tree_add_51_79_groupi_n_9705);
  or csa_tree_add_51_79_groupi_g36175(csa_tree_add_51_79_groupi_n_9876 ,csa_tree_add_51_79_groupi_n_9605 ,csa_tree_add_51_79_groupi_n_9745);
  or csa_tree_add_51_79_groupi_g36176(csa_tree_add_51_79_groupi_n_9875 ,csa_tree_add_51_79_groupi_n_9696 ,csa_tree_add_51_79_groupi_n_9650);
  or csa_tree_add_51_79_groupi_g36177(csa_tree_add_51_79_groupi_n_9874 ,csa_tree_add_51_79_groupi_n_9597 ,csa_tree_add_51_79_groupi_n_9741);
  and csa_tree_add_51_79_groupi_g36178(csa_tree_add_51_79_groupi_n_9947 ,csa_tree_add_51_79_groupi_n_9538 ,csa_tree_add_51_79_groupi_n_9735);
  or csa_tree_add_51_79_groupi_g36179(csa_tree_add_51_79_groupi_n_9945 ,csa_tree_add_51_79_groupi_n_9423 ,csa_tree_add_51_79_groupi_n_9734);
  or csa_tree_add_51_79_groupi_g36180(csa_tree_add_51_79_groupi_n_9944 ,csa_tree_add_51_79_groupi_n_9420 ,csa_tree_add_51_79_groupi_n_9772);
  and csa_tree_add_51_79_groupi_g36181(csa_tree_add_51_79_groupi_n_9943 ,csa_tree_add_51_79_groupi_n_9577 ,csa_tree_add_51_79_groupi_n_9783);
  or csa_tree_add_51_79_groupi_g36182(csa_tree_add_51_79_groupi_n_9941 ,csa_tree_add_51_79_groupi_n_9520 ,csa_tree_add_51_79_groupi_n_9744);
  and csa_tree_add_51_79_groupi_g36183(csa_tree_add_51_79_groupi_n_9940 ,csa_tree_add_51_79_groupi_n_9529 ,csa_tree_add_51_79_groupi_n_9755);
  and csa_tree_add_51_79_groupi_g36184(csa_tree_add_51_79_groupi_n_9939 ,csa_tree_add_51_79_groupi_n_9533 ,csa_tree_add_51_79_groupi_n_9754);
  and csa_tree_add_51_79_groupi_g36185(csa_tree_add_51_79_groupi_n_9938 ,csa_tree_add_51_79_groupi_n_9541 ,csa_tree_add_51_79_groupi_n_9758);
  and csa_tree_add_51_79_groupi_g36186(csa_tree_add_51_79_groupi_n_9937 ,csa_tree_add_51_79_groupi_n_9561 ,csa_tree_add_51_79_groupi_n_9775);
  and csa_tree_add_51_79_groupi_g36187(csa_tree_add_51_79_groupi_n_9936 ,csa_tree_add_51_79_groupi_n_9563 ,csa_tree_add_51_79_groupi_n_9776);
  and csa_tree_add_51_79_groupi_g36188(csa_tree_add_51_79_groupi_n_9935 ,csa_tree_add_51_79_groupi_n_9523 ,csa_tree_add_51_79_groupi_n_9748);
  and csa_tree_add_51_79_groupi_g36189(csa_tree_add_51_79_groupi_n_9934 ,csa_tree_add_51_79_groupi_n_9553 ,csa_tree_add_51_79_groupi_n_9737);
  and csa_tree_add_51_79_groupi_g36190(csa_tree_add_51_79_groupi_n_9932 ,csa_tree_add_51_79_groupi_n_9525 ,csa_tree_add_51_79_groupi_n_9782);
  and csa_tree_add_51_79_groupi_g36191(csa_tree_add_51_79_groupi_n_9931 ,csa_tree_add_51_79_groupi_n_9518 ,csa_tree_add_51_79_groupi_n_9743);
  and csa_tree_add_51_79_groupi_g36192(csa_tree_add_51_79_groupi_n_9930 ,csa_tree_add_51_79_groupi_n_9543 ,csa_tree_add_51_79_groupi_n_9759);
  and csa_tree_add_51_79_groupi_g36193(csa_tree_add_51_79_groupi_n_9929 ,csa_tree_add_51_79_groupi_n_9544 ,csa_tree_add_51_79_groupi_n_9753);
  and csa_tree_add_51_79_groupi_g36194(csa_tree_add_51_79_groupi_n_9926 ,csa_tree_add_51_79_groupi_n_9545 ,csa_tree_add_51_79_groupi_n_9756);
  and csa_tree_add_51_79_groupi_g36195(csa_tree_add_51_79_groupi_n_9925 ,csa_tree_add_51_79_groupi_n_9551 ,csa_tree_add_51_79_groupi_n_9767);
  and csa_tree_add_51_79_groupi_g36196(csa_tree_add_51_79_groupi_n_9924 ,csa_tree_add_51_79_groupi_n_9552 ,csa_tree_add_51_79_groupi_n_9768);
  and csa_tree_add_51_79_groupi_g36197(csa_tree_add_51_79_groupi_n_9923 ,csa_tree_add_51_79_groupi_n_9559 ,csa_tree_add_51_79_groupi_n_9774);
  and csa_tree_add_51_79_groupi_g36198(csa_tree_add_51_79_groupi_n_9922 ,csa_tree_add_51_79_groupi_n_9531 ,csa_tree_add_51_79_groupi_n_9736);
  and csa_tree_add_51_79_groupi_g36199(csa_tree_add_51_79_groupi_n_9921 ,csa_tree_add_51_79_groupi_n_9573 ,csa_tree_add_51_79_groupi_n_9773);
  and csa_tree_add_51_79_groupi_g36200(csa_tree_add_51_79_groupi_n_9919 ,csa_tree_add_51_79_groupi_n_9579 ,csa_tree_add_51_79_groupi_n_9718);
  and csa_tree_add_51_79_groupi_g36201(csa_tree_add_51_79_groupi_n_9918 ,csa_tree_add_51_79_groupi_n_9566 ,csa_tree_add_51_79_groupi_n_9777);
  and csa_tree_add_51_79_groupi_g36202(csa_tree_add_51_79_groupi_n_9917 ,csa_tree_add_51_79_groupi_n_9433 ,csa_tree_add_51_79_groupi_n_9723);
  and csa_tree_add_51_79_groupi_g36203(csa_tree_add_51_79_groupi_n_9916 ,csa_tree_add_51_79_groupi_n_9435 ,csa_tree_add_51_79_groupi_n_9752);
  and csa_tree_add_51_79_groupi_g36204(csa_tree_add_51_79_groupi_n_9914 ,csa_tree_add_51_79_groupi_n_9571 ,csa_tree_add_51_79_groupi_n_9780);
  and csa_tree_add_51_79_groupi_g36205(csa_tree_add_51_79_groupi_n_9913 ,csa_tree_add_51_79_groupi_n_9517 ,csa_tree_add_51_79_groupi_n_9738);
  not csa_tree_add_51_79_groupi_g36206(csa_tree_add_51_79_groupi_n_9868 ,csa_tree_add_51_79_groupi_n_9867);
  not csa_tree_add_51_79_groupi_g36207(csa_tree_add_51_79_groupi_n_9866 ,csa_tree_add_51_79_groupi_n_32);
  not csa_tree_add_51_79_groupi_g36208(csa_tree_add_51_79_groupi_n_9855 ,csa_tree_add_51_79_groupi_n_9854);
  or csa_tree_add_51_79_groupi_g36209(csa_tree_add_51_79_groupi_n_9852 ,csa_tree_add_51_79_groupi_n_9610 ,csa_tree_add_51_79_groupi_n_9654);
  or csa_tree_add_51_79_groupi_g36210(csa_tree_add_51_79_groupi_n_9851 ,csa_tree_add_51_79_groupi_n_9603 ,csa_tree_add_51_79_groupi_n_9760);
  and csa_tree_add_51_79_groupi_g36211(csa_tree_add_51_79_groupi_n_9850 ,csa_tree_add_51_79_groupi_n_9805 ,csa_tree_add_51_79_groupi_n_9786);
  or csa_tree_add_51_79_groupi_g36212(csa_tree_add_51_79_groupi_n_9849 ,csa_tree_add_51_79_groupi_n_9694 ,csa_tree_add_51_79_groupi_n_9649);
  or csa_tree_add_51_79_groupi_g36213(csa_tree_add_51_79_groupi_n_9848 ,csa_tree_add_51_79_groupi_n_9496 ,csa_tree_add_51_79_groupi_n_9691);
  and csa_tree_add_51_79_groupi_g36214(csa_tree_add_51_79_groupi_n_9847 ,csa_tree_add_51_79_groupi_n_9496 ,csa_tree_add_51_79_groupi_n_9691);
  or csa_tree_add_51_79_groupi_g36215(csa_tree_add_51_79_groupi_n_9846 ,csa_tree_add_51_79_groupi_n_9685 ,csa_tree_add_51_79_groupi_n_9690);
  and csa_tree_add_51_79_groupi_g36216(csa_tree_add_51_79_groupi_n_9845 ,csa_tree_add_51_79_groupi_n_9685 ,csa_tree_add_51_79_groupi_n_9690);
  or csa_tree_add_51_79_groupi_g36217(csa_tree_add_51_79_groupi_n_9844 ,csa_tree_add_51_79_groupi_n_9402 ,csa_tree_add_51_79_groupi_n_9652);
  or csa_tree_add_51_79_groupi_g36218(csa_tree_add_51_79_groupi_n_9843 ,csa_tree_add_51_79_groupi_n_9793 ,csa_tree_add_51_79_groupi_n_9443);
  nor csa_tree_add_51_79_groupi_g36219(csa_tree_add_51_79_groupi_n_9842 ,csa_tree_add_51_79_groupi_n_9792 ,csa_tree_add_51_79_groupi_n_9444);
  or csa_tree_add_51_79_groupi_g36220(csa_tree_add_51_79_groupi_n_9841 ,csa_tree_add_51_79_groupi_n_9787 ,csa_tree_add_51_79_groupi_n_9675);
  nor csa_tree_add_51_79_groupi_g36221(csa_tree_add_51_79_groupi_n_9840 ,csa_tree_add_51_79_groupi_n_9788 ,csa_tree_add_51_79_groupi_n_9676);
  nor csa_tree_add_51_79_groupi_g36222(csa_tree_add_51_79_groupi_n_9839 ,csa_tree_add_51_79_groupi_n_9511 ,csa_tree_add_51_79_groupi_n_9663);
  nor csa_tree_add_51_79_groupi_g36223(csa_tree_add_51_79_groupi_n_9838 ,csa_tree_add_51_79_groupi_n_9513 ,csa_tree_add_51_79_groupi_n_9655);
  or csa_tree_add_51_79_groupi_g36224(csa_tree_add_51_79_groupi_n_9837 ,csa_tree_add_51_79_groupi_n_9687 ,csa_tree_add_51_79_groupi_n_9484);
  nor csa_tree_add_51_79_groupi_g36225(csa_tree_add_51_79_groupi_n_9836 ,csa_tree_add_51_79_groupi_n_9688 ,csa_tree_add_51_79_groupi_n_9485);
  xnor csa_tree_add_51_79_groupi_g36226(csa_tree_add_51_79_groupi_n_9835 ,csa_tree_add_51_79_groupi_n_9486 ,csa_tree_add_51_79_groupi_n_9597);
  xnor csa_tree_add_51_79_groupi_g36227(csa_tree_add_51_79_groupi_n_9834 ,csa_tree_add_51_79_groupi_n_9613 ,csa_tree_add_51_79_groupi_n_9498);
  xnor csa_tree_add_51_79_groupi_g36228(csa_tree_add_51_79_groupi_n_9833 ,csa_tree_add_51_79_groupi_n_9483 ,csa_tree_add_51_79_groupi_n_9596);
  xnor csa_tree_add_51_79_groupi_g36229(csa_tree_add_51_79_groupi_n_9832 ,csa_tree_add_51_79_groupi_n_9474 ,csa_tree_add_51_79_groupi_n_9449);
  xnor csa_tree_add_51_79_groupi_g36230(csa_tree_add_51_79_groupi_n_9831 ,csa_tree_add_51_79_groupi_n_9491 ,csa_tree_add_51_79_groupi_n_9488);
  xnor csa_tree_add_51_79_groupi_g36231(csa_tree_add_51_79_groupi_n_9830 ,csa_tree_add_51_79_groupi_n_9462 ,csa_tree_add_51_79_groupi_n_9458);
  xnor csa_tree_add_51_79_groupi_g36232(csa_tree_add_51_79_groupi_n_9829 ,csa_tree_add_51_79_groupi_n_9504 ,csa_tree_add_51_79_groupi_n_9591);
  xnor csa_tree_add_51_79_groupi_g36233(csa_tree_add_51_79_groupi_n_9828 ,csa_tree_add_51_79_groupi_n_9296 ,csa_tree_add_51_79_groupi_n_9469);
  xnor csa_tree_add_51_79_groupi_g36234(csa_tree_add_51_79_groupi_n_9827 ,csa_tree_add_51_79_groupi_n_9082 ,csa_tree_add_51_79_groupi_n_9510);
  xnor csa_tree_add_51_79_groupi_g36235(csa_tree_add_51_79_groupi_n_9826 ,csa_tree_add_51_79_groupi_n_9610 ,csa_tree_add_51_79_groupi_n_9273);
  xnor csa_tree_add_51_79_groupi_g36236(csa_tree_add_51_79_groupi_n_9825 ,csa_tree_add_51_79_groupi_n_9495 ,csa_tree_add_51_79_groupi_n_9493);
  xnor csa_tree_add_51_79_groupi_g36237(csa_tree_add_51_79_groupi_n_9824 ,csa_tree_add_51_79_groupi_n_9279 ,csa_tree_add_51_79_groupi_n_9607);
  xnor csa_tree_add_51_79_groupi_g36238(csa_tree_add_51_79_groupi_n_9823 ,csa_tree_add_51_79_groupi_n_9506 ,csa_tree_add_51_79_groupi_n_9512);
  xnor csa_tree_add_51_79_groupi_g36239(csa_tree_add_51_79_groupi_n_9822 ,csa_tree_add_51_79_groupi_n_9584 ,csa_tree_add_51_79_groupi_n_9446);
  xnor csa_tree_add_51_79_groupi_g36240(csa_tree_add_51_79_groupi_n_9821 ,csa_tree_add_51_79_groupi_n_9479 ,csa_tree_add_51_79_groupi_n_9585);
  xnor csa_tree_add_51_79_groupi_g36241(csa_tree_add_51_79_groupi_n_9820 ,csa_tree_add_51_79_groupi_n_9477 ,csa_tree_add_51_79_groupi_n_9478);
  xnor csa_tree_add_51_79_groupi_g36242(csa_tree_add_51_79_groupi_n_9819 ,csa_tree_add_51_79_groupi_n_9480 ,csa_tree_add_51_79_groupi_n_9197);
  xnor csa_tree_add_51_79_groupi_g36243(csa_tree_add_51_79_groupi_n_9818 ,csa_tree_add_51_79_groupi_n_9476 ,csa_tree_add_51_79_groupi_n_9581);
  xnor csa_tree_add_51_79_groupi_g36244(csa_tree_add_51_79_groupi_n_9817 ,csa_tree_add_51_79_groupi_n_9379 ,csa_tree_add_51_79_groupi_n_9603);
  xnor csa_tree_add_51_79_groupi_g36245(csa_tree_add_51_79_groupi_n_9816 ,csa_tree_add_51_79_groupi_n_9471 ,csa_tree_add_51_79_groupi_n_9472);
  xnor csa_tree_add_51_79_groupi_g36246(csa_tree_add_51_79_groupi_n_9815 ,csa_tree_add_51_79_groupi_n_9450 ,csa_tree_add_51_79_groupi_n_9375);
  xnor csa_tree_add_51_79_groupi_g36247(csa_tree_add_51_79_groupi_n_9814 ,csa_tree_add_51_79_groupi_n_9470 ,csa_tree_add_51_79_groupi_n_9380);
  xnor csa_tree_add_51_79_groupi_g36248(csa_tree_add_51_79_groupi_n_9813 ,csa_tree_add_51_79_groupi_n_9608 ,csa_tree_add_51_79_groupi_n_9358);
  xnor csa_tree_add_51_79_groupi_g36249(csa_tree_add_51_79_groupi_n_9812 ,csa_tree_add_51_79_groupi_n_9459 ,csa_tree_add_51_79_groupi_n_9460);
  xnor csa_tree_add_51_79_groupi_g36250(csa_tree_add_51_79_groupi_n_9811 ,csa_tree_add_51_79_groupi_n_9599 ,csa_tree_add_51_79_groupi_n_9376);
  xnor csa_tree_add_51_79_groupi_g36251(csa_tree_add_51_79_groupi_n_9810 ,csa_tree_add_51_79_groupi_n_9588 ,csa_tree_add_51_79_groupi_n_9454);
  xnor csa_tree_add_51_79_groupi_g36252(csa_tree_add_51_79_groupi_n_9809 ,csa_tree_add_51_79_groupi_n_9441 ,csa_tree_add_51_79_groupi_n_9442);
  xnor csa_tree_add_51_79_groupi_g36253(csa_tree_add_51_79_groupi_n_9808 ,csa_tree_add_51_79_groupi_n_9440 ,csa_tree_add_51_79_groupi_n_9181);
  xor csa_tree_add_51_79_groupi_g36254(csa_tree_add_51_79_groupi_n_9807 ,csa_tree_add_51_79_groupi_n_9438 ,csa_tree_add_51_79_groupi_n_9600);
  xnor csa_tree_add_51_79_groupi_g36255(csa_tree_add_51_79_groupi_n_9806 ,csa_tree_add_51_79_groupi_n_9485 ,csa_tree_add_51_79_groupi_n_9598);
  xnor csa_tree_add_51_79_groupi_g36256(csa_tree_add_51_79_groupi_n_9873 ,csa_tree_add_51_79_groupi_n_9298 ,csa_tree_add_51_79_groupi_n_9408);
  xnor csa_tree_add_51_79_groupi_g36257(csa_tree_add_51_79_groupi_n_9872 ,csa_tree_add_51_79_groupi_n_8770 ,csa_tree_add_51_79_groupi_n_9412);
  xnor csa_tree_add_51_79_groupi_g36258(csa_tree_add_51_79_groupi_n_9871 ,csa_tree_add_51_79_groupi_n_9085 ,csa_tree_add_51_79_groupi_n_9417);
  xnor csa_tree_add_51_79_groupi_g36259(csa_tree_add_51_79_groupi_n_9870 ,csa_tree_add_51_79_groupi_n_8795 ,csa_tree_add_51_79_groupi_n_9407);
  and csa_tree_add_51_79_groupi_g36260(csa_tree_add_51_79_groupi_n_9869 ,csa_tree_add_51_79_groupi_n_9427 ,csa_tree_add_51_79_groupi_n_9770);
  xnor csa_tree_add_51_79_groupi_g36261(csa_tree_add_51_79_groupi_n_9867 ,csa_tree_add_51_79_groupi_n_9278 ,csa_tree_add_51_79_groupi_n_9416);
  xnor csa_tree_add_51_79_groupi_g36263(csa_tree_add_51_79_groupi_n_9865 ,csa_tree_add_51_79_groupi_n_9203 ,csa_tree_add_51_79_groupi_n_9409);
  xnor csa_tree_add_51_79_groupi_g36264(csa_tree_add_51_79_groupi_n_9864 ,csa_tree_add_51_79_groupi_n_8750 ,csa_tree_add_51_79_groupi_n_9418);
  xnor csa_tree_add_51_79_groupi_g36265(csa_tree_add_51_79_groupi_n_9863 ,csa_tree_add_51_79_groupi_n_9489 ,csa_tree_add_51_79_groupi_n_9406);
  and csa_tree_add_51_79_groupi_g36266(csa_tree_add_51_79_groupi_n_9862 ,csa_tree_add_51_79_groupi_n_9429 ,csa_tree_add_51_79_groupi_n_9766);
  and csa_tree_add_51_79_groupi_g36267(csa_tree_add_51_79_groupi_n_9861 ,csa_tree_add_51_79_groupi_n_9431 ,csa_tree_add_51_79_groupi_n_9765);
  xnor csa_tree_add_51_79_groupi_g36268(csa_tree_add_51_79_groupi_n_9860 ,csa_tree_add_51_79_groupi_n_9401 ,csa_tree_add_51_79_groupi_n_9419);
  xnor csa_tree_add_51_79_groupi_g36270(csa_tree_add_51_79_groupi_n_9859 ,csa_tree_add_51_79_groupi_n_9202 ,csa_tree_add_51_79_groupi_n_9404);
  xnor csa_tree_add_51_79_groupi_g36271(csa_tree_add_51_79_groupi_n_9858 ,csa_tree_add_51_79_groupi_n_9286 ,csa_tree_add_51_79_groupi_n_9405);
  xnor csa_tree_add_51_79_groupi_g36272(csa_tree_add_51_79_groupi_n_9857 ,csa_tree_add_51_79_groupi_n_9176 ,csa_tree_add_51_79_groupi_n_9415);
  xnor csa_tree_add_51_79_groupi_g36273(csa_tree_add_51_79_groupi_n_9856 ,csa_tree_add_51_79_groupi_n_8742 ,csa_tree_add_51_79_groupi_n_9414);
  and csa_tree_add_51_79_groupi_g36274(csa_tree_add_51_79_groupi_n_9854 ,csa_tree_add_51_79_groupi_n_9536 ,csa_tree_add_51_79_groupi_n_9658);
  xnor csa_tree_add_51_79_groupi_g36275(csa_tree_add_51_79_groupi_n_9853 ,csa_tree_add_51_79_groupi_n_8755 ,csa_tree_add_51_79_groupi_n_9410);
  not csa_tree_add_51_79_groupi_g36276(csa_tree_add_51_79_groupi_n_9799 ,csa_tree_add_51_79_groupi_n_9798);
  not csa_tree_add_51_79_groupi_g36277(csa_tree_add_51_79_groupi_n_9794 ,csa_tree_add_51_79_groupi_n_9795);
  not csa_tree_add_51_79_groupi_g36278(csa_tree_add_51_79_groupi_n_9792 ,csa_tree_add_51_79_groupi_n_9793);
  not csa_tree_add_51_79_groupi_g36279(csa_tree_add_51_79_groupi_n_9791 ,csa_tree_add_51_79_groupi_n_9790);
  not csa_tree_add_51_79_groupi_g36280(csa_tree_add_51_79_groupi_n_9788 ,csa_tree_add_51_79_groupi_n_9787);
  or csa_tree_add_51_79_groupi_g36281(csa_tree_add_51_79_groupi_n_9786 ,csa_tree_add_51_79_groupi_n_9473 ,csa_tree_add_51_79_groupi_n_9449);
  or csa_tree_add_51_79_groupi_g36282(csa_tree_add_51_79_groupi_n_9785 ,csa_tree_add_51_79_groupi_n_9587 ,csa_tree_add_51_79_groupi_n_9483);
  and csa_tree_add_51_79_groupi_g36283(csa_tree_add_51_79_groupi_n_9784 ,csa_tree_add_51_79_groupi_n_9587 ,csa_tree_add_51_79_groupi_n_9483);
  or csa_tree_add_51_79_groupi_g36284(csa_tree_add_51_79_groupi_n_9783 ,csa_tree_add_51_79_groupi_n_8969 ,csa_tree_add_51_79_groupi_n_9558);
  or csa_tree_add_51_79_groupi_g36285(csa_tree_add_51_79_groupi_n_9782 ,csa_tree_add_51_79_groupi_n_8963 ,csa_tree_add_51_79_groupi_n_9574);
  nor csa_tree_add_51_79_groupi_g36286(csa_tree_add_51_79_groupi_n_9781 ,csa_tree_add_51_79_groupi_n_9474 ,csa_tree_add_51_79_groupi_n_9448);
  or csa_tree_add_51_79_groupi_g36287(csa_tree_add_51_79_groupi_n_9780 ,csa_tree_add_51_79_groupi_n_9305 ,csa_tree_add_51_79_groupi_n_9570);
  and csa_tree_add_51_79_groupi_g36288(csa_tree_add_51_79_groupi_n_9779 ,csa_tree_add_51_79_groupi_n_9586 ,csa_tree_add_51_79_groupi_n_9438);
  nor csa_tree_add_51_79_groupi_g36289(csa_tree_add_51_79_groupi_n_9778 ,csa_tree_add_51_79_groupi_n_9586 ,csa_tree_add_51_79_groupi_n_9438);
  or csa_tree_add_51_79_groupi_g36290(csa_tree_add_51_79_groupi_n_9777 ,csa_tree_add_51_79_groupi_n_9392 ,csa_tree_add_51_79_groupi_n_9564);
  or csa_tree_add_51_79_groupi_g36291(csa_tree_add_51_79_groupi_n_9776 ,csa_tree_add_51_79_groupi_n_9398 ,csa_tree_add_51_79_groupi_n_9562);
  or csa_tree_add_51_79_groupi_g36292(csa_tree_add_51_79_groupi_n_9775 ,csa_tree_add_51_79_groupi_n_9199 ,csa_tree_add_51_79_groupi_n_9560);
  or csa_tree_add_51_79_groupi_g36293(csa_tree_add_51_79_groupi_n_9774 ,csa_tree_add_51_79_groupi_n_9389 ,csa_tree_add_51_79_groupi_n_9557);
  or csa_tree_add_51_79_groupi_g36294(csa_tree_add_51_79_groupi_n_9773 ,csa_tree_add_51_79_groupi_n_9395 ,csa_tree_add_51_79_groupi_n_9556);
  and csa_tree_add_51_79_groupi_g36295(csa_tree_add_51_79_groupi_n_9772 ,csa_tree_add_51_79_groupi_n_9391 ,csa_tree_add_51_79_groupi_n_9421);
  or csa_tree_add_51_79_groupi_g36296(csa_tree_add_51_79_groupi_n_9771 ,csa_tree_add_51_79_groupi_n_9581 ,csa_tree_add_51_79_groupi_n_9476);
  or csa_tree_add_51_79_groupi_g36297(csa_tree_add_51_79_groupi_n_9770 ,csa_tree_add_51_79_groupi_n_9426 ,csa_tree_add_51_79_groupi_n_9514);
  and csa_tree_add_51_79_groupi_g36298(csa_tree_add_51_79_groupi_n_9769 ,csa_tree_add_51_79_groupi_n_9581 ,csa_tree_add_51_79_groupi_n_9476);
  or csa_tree_add_51_79_groupi_g36299(csa_tree_add_51_79_groupi_n_9768 ,csa_tree_add_51_79_groupi_n_9200 ,csa_tree_add_51_79_groupi_n_9547);
  or csa_tree_add_51_79_groupi_g36300(csa_tree_add_51_79_groupi_n_9767 ,csa_tree_add_51_79_groupi_n_9509 ,csa_tree_add_51_79_groupi_n_9550);
  or csa_tree_add_51_79_groupi_g36301(csa_tree_add_51_79_groupi_n_9766 ,csa_tree_add_51_79_groupi_n_9303 ,csa_tree_add_51_79_groupi_n_9428);
  or csa_tree_add_51_79_groupi_g36302(csa_tree_add_51_79_groupi_n_9765 ,csa_tree_add_51_79_groupi_n_9397 ,csa_tree_add_51_79_groupi_n_9430);
  and csa_tree_add_51_79_groupi_g36303(csa_tree_add_51_79_groupi_n_9764 ,csa_tree_add_51_79_groupi_n_9279 ,csa_tree_add_51_79_groupi_n_9451);
  nor csa_tree_add_51_79_groupi_g36304(csa_tree_add_51_79_groupi_n_9763 ,csa_tree_add_51_79_groupi_n_9279 ,csa_tree_add_51_79_groupi_n_9451);
  or csa_tree_add_51_79_groupi_g36305(csa_tree_add_51_79_groupi_n_9762 ,csa_tree_add_51_79_groupi_n_9380 ,csa_tree_add_51_79_groupi_n_9470);
  and csa_tree_add_51_79_groupi_g36306(csa_tree_add_51_79_groupi_n_9761 ,csa_tree_add_51_79_groupi_n_9380 ,csa_tree_add_51_79_groupi_n_9470);
  and csa_tree_add_51_79_groupi_g36307(csa_tree_add_51_79_groupi_n_9760 ,csa_tree_add_51_79_groupi_n_9482 ,csa_tree_add_51_79_groupi_n_9379);
  or csa_tree_add_51_79_groupi_g36308(csa_tree_add_51_79_groupi_n_9759 ,csa_tree_add_51_79_groupi_n_9390 ,csa_tree_add_51_79_groupi_n_9542);
  or csa_tree_add_51_79_groupi_g36309(csa_tree_add_51_79_groupi_n_9758 ,csa_tree_add_51_79_groupi_n_9299 ,csa_tree_add_51_79_groupi_n_9539);
  or csa_tree_add_51_79_groupi_g36310(csa_tree_add_51_79_groupi_n_9757 ,csa_tree_add_51_79_groupi_n_9482 ,csa_tree_add_51_79_groupi_n_9379);
  or csa_tree_add_51_79_groupi_g36311(csa_tree_add_51_79_groupi_n_9756 ,csa_tree_add_51_79_groupi_n_9393 ,csa_tree_add_51_79_groupi_n_9534);
  or csa_tree_add_51_79_groupi_g36312(csa_tree_add_51_79_groupi_n_9755 ,csa_tree_add_51_79_groupi_n_9301 ,csa_tree_add_51_79_groupi_n_9526);
  or csa_tree_add_51_79_groupi_g36313(csa_tree_add_51_79_groupi_n_9754 ,csa_tree_add_51_79_groupi_n_9385 ,csa_tree_add_51_79_groupi_n_9528);
  or csa_tree_add_51_79_groupi_g36314(csa_tree_add_51_79_groupi_n_9753 ,csa_tree_add_51_79_groupi_n_9400 ,csa_tree_add_51_79_groupi_n_9519);
  or csa_tree_add_51_79_groupi_g36315(csa_tree_add_51_79_groupi_n_9752 ,csa_tree_add_51_79_groupi_n_8966 ,csa_tree_add_51_79_groupi_n_9434);
  or csa_tree_add_51_79_groupi_g36316(csa_tree_add_51_79_groupi_n_9751 ,csa_tree_add_51_79_groupi_n_9497 ,csa_tree_add_51_79_groupi_n_9499);
  or csa_tree_add_51_79_groupi_g36317(csa_tree_add_51_79_groupi_n_9750 ,csa_tree_add_51_79_groupi_n_9442 ,csa_tree_add_51_79_groupi_n_9441);
  and csa_tree_add_51_79_groupi_g36318(csa_tree_add_51_79_groupi_n_9749 ,csa_tree_add_51_79_groupi_n_9442 ,csa_tree_add_51_79_groupi_n_9441);
  or csa_tree_add_51_79_groupi_g36319(csa_tree_add_51_79_groupi_n_9748 ,csa_tree_add_51_79_groupi_n_9396 ,csa_tree_add_51_79_groupi_n_9522);
  nor csa_tree_add_51_79_groupi_g36320(csa_tree_add_51_79_groupi_n_9747 ,csa_tree_add_51_79_groupi_n_9498 ,csa_tree_add_51_79_groupi_n_9500);
  or csa_tree_add_51_79_groupi_g36321(csa_tree_add_51_79_groupi_n_9746 ,csa_tree_add_51_79_groupi_n_9181 ,csa_tree_add_51_79_groupi_n_9440);
  and csa_tree_add_51_79_groupi_g36322(csa_tree_add_51_79_groupi_n_9745 ,csa_tree_add_51_79_groupi_n_9181 ,csa_tree_add_51_79_groupi_n_9440);
  and csa_tree_add_51_79_groupi_g36323(csa_tree_add_51_79_groupi_n_9744 ,csa_tree_add_51_79_groupi_n_9595 ,csa_tree_add_51_79_groupi_n_9524);
  or csa_tree_add_51_79_groupi_g36324(csa_tree_add_51_79_groupi_n_9743 ,csa_tree_add_51_79_groupi_n_9308 ,csa_tree_add_51_79_groupi_n_9521);
  or csa_tree_add_51_79_groupi_g36325(csa_tree_add_51_79_groupi_n_9742 ,csa_tree_add_51_79_groupi_n_9439 ,csa_tree_add_51_79_groupi_n_9486);
  and csa_tree_add_51_79_groupi_g36326(csa_tree_add_51_79_groupi_n_9741 ,csa_tree_add_51_79_groupi_n_9439 ,csa_tree_add_51_79_groupi_n_9486);
  or csa_tree_add_51_79_groupi_g36327(csa_tree_add_51_79_groupi_n_9740 ,csa_tree_add_51_79_groupi_n_9296 ,csa_tree_add_51_79_groupi_n_9468);
  nor csa_tree_add_51_79_groupi_g36328(csa_tree_add_51_79_groupi_n_9739 ,csa_tree_add_51_79_groupi_n_9295 ,csa_tree_add_51_79_groupi_n_9469);
  or csa_tree_add_51_79_groupi_g36329(csa_tree_add_51_79_groupi_n_9738 ,csa_tree_add_51_79_groupi_n_9306 ,csa_tree_add_51_79_groupi_n_9530);
  or csa_tree_add_51_79_groupi_g36330(csa_tree_add_51_79_groupi_n_9737 ,csa_tree_add_51_79_groupi_n_9205 ,csa_tree_add_51_79_groupi_n_9554);
  or csa_tree_add_51_79_groupi_g36331(csa_tree_add_51_79_groupi_n_9736 ,csa_tree_add_51_79_groupi_n_9383 ,csa_tree_add_51_79_groupi_n_9546);
  or csa_tree_add_51_79_groupi_g36332(csa_tree_add_51_79_groupi_n_9735 ,csa_tree_add_51_79_groupi_n_9384 ,csa_tree_add_51_79_groupi_n_9580);
  nor csa_tree_add_51_79_groupi_g36333(csa_tree_add_51_79_groupi_n_9734 ,csa_tree_add_51_79_groupi_n_9387 ,csa_tree_add_51_79_groupi_n_9422);
  or csa_tree_add_51_79_groupi_g36334(csa_tree_add_51_79_groupi_n_9733 ,csa_tree_add_51_79_groupi_n_9481 ,csa_tree_add_51_79_groupi_n_9480);
  and csa_tree_add_51_79_groupi_g36335(csa_tree_add_51_79_groupi_n_9732 ,csa_tree_add_51_79_groupi_n_9481 ,csa_tree_add_51_79_groupi_n_9480);
  or csa_tree_add_51_79_groupi_g36336(csa_tree_add_51_79_groupi_n_9731 ,csa_tree_add_51_79_groupi_n_9585 ,csa_tree_add_51_79_groupi_n_9479);
  and csa_tree_add_51_79_groupi_g36337(csa_tree_add_51_79_groupi_n_9730 ,csa_tree_add_51_79_groupi_n_9585 ,csa_tree_add_51_79_groupi_n_9479);
  or csa_tree_add_51_79_groupi_g36338(csa_tree_add_51_79_groupi_n_9729 ,csa_tree_add_51_79_groupi_n_9478 ,csa_tree_add_51_79_groupi_n_9477);
  and csa_tree_add_51_79_groupi_g36339(csa_tree_add_51_79_groupi_n_9728 ,csa_tree_add_51_79_groupi_n_9478 ,csa_tree_add_51_79_groupi_n_9477);
  or csa_tree_add_51_79_groupi_g36340(csa_tree_add_51_79_groupi_n_9727 ,csa_tree_add_51_79_groupi_n_9472 ,csa_tree_add_51_79_groupi_n_9471);
  and csa_tree_add_51_79_groupi_g36341(csa_tree_add_51_79_groupi_n_9726 ,csa_tree_add_51_79_groupi_n_9472 ,csa_tree_add_51_79_groupi_n_9471);
  or csa_tree_add_51_79_groupi_g36342(csa_tree_add_51_79_groupi_n_9725 ,csa_tree_add_51_79_groupi_n_9465 ,csa_tree_add_51_79_groupi_n_9464);
  and csa_tree_add_51_79_groupi_g36343(csa_tree_add_51_79_groupi_n_9724 ,csa_tree_add_51_79_groupi_n_9465 ,csa_tree_add_51_79_groupi_n_9464);
  or csa_tree_add_51_79_groupi_g36344(csa_tree_add_51_79_groupi_n_9723 ,csa_tree_add_51_79_groupi_n_9297 ,csa_tree_add_51_79_groupi_n_9432);
  or csa_tree_add_51_79_groupi_g36345(csa_tree_add_51_79_groupi_n_9722 ,csa_tree_add_51_79_groupi_n_9358 ,csa_tree_add_51_79_groupi_n_9461);
  and csa_tree_add_51_79_groupi_g36346(csa_tree_add_51_79_groupi_n_9721 ,csa_tree_add_51_79_groupi_n_9358 ,csa_tree_add_51_79_groupi_n_9461);
  or csa_tree_add_51_79_groupi_g36347(csa_tree_add_51_79_groupi_n_9720 ,csa_tree_add_51_79_groupi_n_9460 ,csa_tree_add_51_79_groupi_n_9459);
  and csa_tree_add_51_79_groupi_g36348(csa_tree_add_51_79_groupi_n_9719 ,csa_tree_add_51_79_groupi_n_9460 ,csa_tree_add_51_79_groupi_n_9459);
  or csa_tree_add_51_79_groupi_g36349(csa_tree_add_51_79_groupi_n_9718 ,csa_tree_add_51_79_groupi_n_9403 ,csa_tree_add_51_79_groupi_n_9437);
  or csa_tree_add_51_79_groupi_g36350(csa_tree_add_51_79_groupi_n_9717 ,csa_tree_add_51_79_groupi_n_9376 ,csa_tree_add_51_79_groupi_n_9456);
  and csa_tree_add_51_79_groupi_g36351(csa_tree_add_51_79_groupi_n_9716 ,csa_tree_add_51_79_groupi_n_9376 ,csa_tree_add_51_79_groupi_n_9456);
  or csa_tree_add_51_79_groupi_g36352(csa_tree_add_51_79_groupi_n_9715 ,csa_tree_add_51_79_groupi_n_9454 ,csa_tree_add_51_79_groupi_n_9588);
  and csa_tree_add_51_79_groupi_g36353(csa_tree_add_51_79_groupi_n_9714 ,csa_tree_add_51_79_groupi_n_9454 ,csa_tree_add_51_79_groupi_n_9588);
  or csa_tree_add_51_79_groupi_g36354(csa_tree_add_51_79_groupi_n_9713 ,csa_tree_add_51_79_groupi_n_9375 ,csa_tree_add_51_79_groupi_n_9450);
  and csa_tree_add_51_79_groupi_g36355(csa_tree_add_51_79_groupi_n_9712 ,csa_tree_add_51_79_groupi_n_9375 ,csa_tree_add_51_79_groupi_n_9450);
  or csa_tree_add_51_79_groupi_g36356(csa_tree_add_51_79_groupi_n_9711 ,csa_tree_add_51_79_groupi_n_8775 ,csa_tree_add_51_79_groupi_n_9447);
  and csa_tree_add_51_79_groupi_g36357(csa_tree_add_51_79_groupi_n_9710 ,csa_tree_add_51_79_groupi_n_8775 ,csa_tree_add_51_79_groupi_n_9447);
  or csa_tree_add_51_79_groupi_g36358(csa_tree_add_51_79_groupi_n_9805 ,csa_tree_add_51_79_groupi_n_9245 ,csa_tree_add_51_79_groupi_n_9575);
  and csa_tree_add_51_79_groupi_g36359(csa_tree_add_51_79_groupi_n_9804 ,csa_tree_add_51_79_groupi_n_9311 ,csa_tree_add_51_79_groupi_n_9436);
  and csa_tree_add_51_79_groupi_g36360(csa_tree_add_51_79_groupi_n_9803 ,csa_tree_add_51_79_groupi_n_9344 ,csa_tree_add_51_79_groupi_n_9568);
  and csa_tree_add_51_79_groupi_g36361(csa_tree_add_51_79_groupi_n_9802 ,csa_tree_add_51_79_groupi_n_9340 ,csa_tree_add_51_79_groupi_n_9555);
  and csa_tree_add_51_79_groupi_g36362(csa_tree_add_51_79_groupi_n_9801 ,csa_tree_add_51_79_groupi_n_9060 ,csa_tree_add_51_79_groupi_n_9527);
  and csa_tree_add_51_79_groupi_g36363(csa_tree_add_51_79_groupi_n_9800 ,csa_tree_add_51_79_groupi_n_9332 ,csa_tree_add_51_79_groupi_n_9548);
  or csa_tree_add_51_79_groupi_g36364(csa_tree_add_51_79_groupi_n_9798 ,csa_tree_add_51_79_groupi_n_9353 ,csa_tree_add_51_79_groupi_n_9572);
  and csa_tree_add_51_79_groupi_g36365(csa_tree_add_51_79_groupi_n_9797 ,csa_tree_add_51_79_groupi_n_9314 ,csa_tree_add_51_79_groupi_n_9537);
  and csa_tree_add_51_79_groupi_g36366(csa_tree_add_51_79_groupi_n_9796 ,csa_tree_add_51_79_groupi_n_9322 ,csa_tree_add_51_79_groupi_n_9540);
  or csa_tree_add_51_79_groupi_g36367(csa_tree_add_51_79_groupi_n_9795 ,csa_tree_add_51_79_groupi_n_9239 ,csa_tree_add_51_79_groupi_n_9535);
  and csa_tree_add_51_79_groupi_g36368(csa_tree_add_51_79_groupi_n_9793 ,csa_tree_add_51_79_groupi_n_9092 ,csa_tree_add_51_79_groupi_n_9578);
  or csa_tree_add_51_79_groupi_g36369(csa_tree_add_51_79_groupi_n_9790 ,csa_tree_add_51_79_groupi_n_9329 ,csa_tree_add_51_79_groupi_n_9549);
  and csa_tree_add_51_79_groupi_g36370(csa_tree_add_51_79_groupi_n_9789 ,csa_tree_add_51_79_groupi_n_9350 ,csa_tree_add_51_79_groupi_n_9567);
  or csa_tree_add_51_79_groupi_g36371(csa_tree_add_51_79_groupi_n_9787 ,csa_tree_add_51_79_groupi_n_9247 ,csa_tree_add_51_79_groupi_n_9576);
  not csa_tree_add_51_79_groupi_g36372(csa_tree_add_51_79_groupi_n_9709 ,csa_tree_add_51_79_groupi_n_9708);
  not csa_tree_add_51_79_groupi_g36373(csa_tree_add_51_79_groupi_n_9688 ,csa_tree_add_51_79_groupi_n_9687);
  not csa_tree_add_51_79_groupi_g36374(csa_tree_add_51_79_groupi_n_9679 ,csa_tree_add_51_79_groupi_n_9678);
  not csa_tree_add_51_79_groupi_g36375(csa_tree_add_51_79_groupi_n_9675 ,csa_tree_add_51_79_groupi_n_9676);
  or csa_tree_add_51_79_groupi_g36376(csa_tree_add_51_79_groupi_n_9673 ,csa_tree_add_51_79_groupi_n_9462 ,csa_tree_add_51_79_groupi_n_9458);
  or csa_tree_add_51_79_groupi_g36377(csa_tree_add_51_79_groupi_n_9672 ,csa_tree_add_51_79_groupi_n_9276 ,csa_tree_add_51_79_groupi_n_9463);
  and csa_tree_add_51_79_groupi_g36378(csa_tree_add_51_79_groupi_n_9671 ,csa_tree_add_51_79_groupi_n_9276 ,csa_tree_add_51_79_groupi_n_9463);
  and csa_tree_add_51_79_groupi_g36379(csa_tree_add_51_79_groupi_n_9670 ,csa_tree_add_51_79_groupi_n_9079 ,csa_tree_add_51_79_groupi_n_9489);
  or csa_tree_add_51_79_groupi_g36380(csa_tree_add_51_79_groupi_n_9669 ,csa_tree_add_51_79_groupi_n_9079 ,csa_tree_add_51_79_groupi_n_9489);
  nor csa_tree_add_51_79_groupi_g36381(csa_tree_add_51_79_groupi_n_9668 ,csa_tree_add_51_79_groupi_n_9503 ,csa_tree_add_51_79_groupi_n_9591);
  or csa_tree_add_51_79_groupi_g36382(csa_tree_add_51_79_groupi_n_9667 ,csa_tree_add_51_79_groupi_n_9504 ,csa_tree_add_51_79_groupi_n_9590);
  or csa_tree_add_51_79_groupi_g36383(csa_tree_add_51_79_groupi_n_9666 ,csa_tree_add_51_79_groupi_n_9292 ,csa_tree_add_51_79_groupi_n_9501);
  nor csa_tree_add_51_79_groupi_g36384(csa_tree_add_51_79_groupi_n_9665 ,csa_tree_add_51_79_groupi_n_9293 ,csa_tree_add_51_79_groupi_n_9502);
  nor csa_tree_add_51_79_groupi_g36385(csa_tree_add_51_79_groupi_n_9664 ,csa_tree_add_51_79_groupi_n_9082 ,csa_tree_add_51_79_groupi_n_9467);
  and csa_tree_add_51_79_groupi_g36386(csa_tree_add_51_79_groupi_n_9663 ,csa_tree_add_51_79_groupi_n_9082 ,csa_tree_add_51_79_groupi_n_9467);
  and csa_tree_add_51_79_groupi_g36387(csa_tree_add_51_79_groupi_n_9662 ,csa_tree_add_51_79_groupi_n_9462 ,csa_tree_add_51_79_groupi_n_9458);
  or csa_tree_add_51_79_groupi_g36388(csa_tree_add_51_79_groupi_n_9661 ,csa_tree_add_51_79_groupi_n_9475 ,csa_tree_add_51_79_groupi_n_9457);
  or csa_tree_add_51_79_groupi_g36389(csa_tree_add_51_79_groupi_n_9660 ,csa_tree_add_51_79_groupi_n_9584 ,csa_tree_add_51_79_groupi_n_9445);
  nor csa_tree_add_51_79_groupi_g36390(csa_tree_add_51_79_groupi_n_9659 ,csa_tree_add_51_79_groupi_n_9583 ,csa_tree_add_51_79_groupi_n_9446);
  or csa_tree_add_51_79_groupi_g36391(csa_tree_add_51_79_groupi_n_9658 ,csa_tree_add_51_79_groupi_n_9532 ,csa_tree_add_51_79_groupi_n_9609);
  or csa_tree_add_51_79_groupi_g36392(csa_tree_add_51_79_groupi_n_9657 ,csa_tree_add_51_79_groupi_n_9507 ,csa_tree_add_51_79_groupi_n_9272);
  nor csa_tree_add_51_79_groupi_g36393(csa_tree_add_51_79_groupi_n_9656 ,csa_tree_add_51_79_groupi_n_9506 ,csa_tree_add_51_79_groupi_n_9505);
  and csa_tree_add_51_79_groupi_g36394(csa_tree_add_51_79_groupi_n_9655 ,csa_tree_add_51_79_groupi_n_9506 ,csa_tree_add_51_79_groupi_n_9505);
  nor csa_tree_add_51_79_groupi_g36395(csa_tree_add_51_79_groupi_n_9654 ,csa_tree_add_51_79_groupi_n_9508 ,csa_tree_add_51_79_groupi_n_9273);
  or csa_tree_add_51_79_groupi_g36396(csa_tree_add_51_79_groupi_n_9653 ,csa_tree_add_51_79_groupi_n_9494 ,csa_tree_add_51_79_groupi_n_9492);
  nor csa_tree_add_51_79_groupi_g36397(csa_tree_add_51_79_groupi_n_9652 ,csa_tree_add_51_79_groupi_n_9495 ,csa_tree_add_51_79_groupi_n_9493);
  or csa_tree_add_51_79_groupi_g36398(csa_tree_add_51_79_groupi_n_9651 ,csa_tree_add_51_79_groupi_n_9491 ,csa_tree_add_51_79_groupi_n_9487);
  nor csa_tree_add_51_79_groupi_g36399(csa_tree_add_51_79_groupi_n_9650 ,csa_tree_add_51_79_groupi_n_9490 ,csa_tree_add_51_79_groupi_n_9488);
  and csa_tree_add_51_79_groupi_g36400(csa_tree_add_51_79_groupi_n_9649 ,csa_tree_add_51_79_groupi_n_9475 ,csa_tree_add_51_79_groupi_n_9457);
  xor csa_tree_add_51_79_groupi_g36401(csa_tree_add_51_79_groupi_n_9648 ,csa_tree_add_51_79_groupi_n_9393 ,csa_tree_add_51_79_groupi_n_9193);
  xnor csa_tree_add_51_79_groupi_g36402(csa_tree_add_51_79_groupi_n_9647 ,csa_tree_add_51_79_groupi_n_9257 ,csa_tree_add_51_79_groupi_n_9200);
  xnor csa_tree_add_51_79_groupi_g36403(csa_tree_add_51_79_groupi_n_9646 ,csa_tree_add_51_79_groupi_n_9365 ,csa_tree_add_51_79_groupi_n_9356);
  xnor csa_tree_add_51_79_groupi_g36404(csa_tree_add_51_79_groupi_n_9645 ,csa_tree_add_51_79_groupi_n_9367 ,csa_tree_add_51_79_groupi_n_9359);
  xnor csa_tree_add_51_79_groupi_g36405(csa_tree_add_51_79_groupi_n_9644 ,csa_tree_add_51_79_groupi_n_8777 ,csa_tree_add_51_79_groupi_n_9304);
  xor csa_tree_add_51_79_groupi_g36406(csa_tree_add_51_79_groupi_n_9643 ,csa_tree_add_51_79_groupi_n_9308 ,csa_tree_add_51_79_groupi_n_9191);
  xnor csa_tree_add_51_79_groupi_g36407(csa_tree_add_51_79_groupi_n_9642 ,csa_tree_add_51_79_groupi_n_9199 ,csa_tree_add_51_79_groupi_n_9366);
  xnor csa_tree_add_51_79_groupi_g36408(csa_tree_add_51_79_groupi_n_9641 ,csa_tree_add_51_79_groupi_n_9388 ,csa_tree_add_51_79_groupi_n_8775);
  xnor csa_tree_add_51_79_groupi_g36409(csa_tree_add_51_79_groupi_n_9640 ,csa_tree_add_51_79_groupi_n_9293 ,csa_tree_add_51_79_groupi_n_9307);
  xor csa_tree_add_51_79_groupi_g36410(csa_tree_add_51_79_groupi_n_9639 ,csa_tree_add_51_79_groupi_n_9306 ,csa_tree_add_51_79_groupi_n_9190);
  xnor csa_tree_add_51_79_groupi_g36411(csa_tree_add_51_79_groupi_n_9638 ,csa_tree_add_51_79_groupi_n_9384 ,csa_tree_add_51_79_groupi_n_9369);
  xnor csa_tree_add_51_79_groupi_g36412(csa_tree_add_51_79_groupi_n_9637 ,csa_tree_add_51_79_groupi_n_9390 ,csa_tree_add_51_79_groupi_n_9378);
  xnor csa_tree_add_51_79_groupi_g36413(csa_tree_add_51_79_groupi_n_9636 ,csa_tree_add_51_79_groupi_n_9268 ,csa_tree_add_51_79_groupi_n_9195);
  xnor csa_tree_add_51_79_groupi_g36414(csa_tree_add_51_79_groupi_n_9635 ,csa_tree_add_51_79_groupi_n_9187 ,csa_tree_add_51_79_groupi_n_9394);
  xnor csa_tree_add_51_79_groupi_g36415(csa_tree_add_51_79_groupi_n_9634 ,csa_tree_add_51_79_groupi_n_9372 ,csa_tree_add_51_79_groupi_n_9185);
  xnor csa_tree_add_51_79_groupi_g36416(csa_tree_add_51_79_groupi_n_9633 ,csa_tree_add_51_79_groupi_n_9387 ,csa_tree_add_51_79_groupi_n_9288);
  xnor csa_tree_add_51_79_groupi_g36417(csa_tree_add_51_79_groupi_n_9632 ,csa_tree_add_51_79_groupi_n_9276 ,csa_tree_add_51_79_groupi_n_9386);
  xnor csa_tree_add_51_79_groupi_g36418(csa_tree_add_51_79_groupi_n_9631 ,csa_tree_add_51_79_groupi_n_9261 ,csa_tree_add_51_79_groupi_n_9281);
  xnor csa_tree_add_51_79_groupi_g36419(csa_tree_add_51_79_groupi_n_9630 ,csa_tree_add_51_79_groupi_n_9285 ,csa_tree_add_51_79_groupi_n_9403);
  xnor csa_tree_add_51_79_groupi_g36420(csa_tree_add_51_79_groupi_n_9629 ,csa_tree_add_51_79_groupi_n_9258 ,csa_tree_add_51_79_groupi_n_9284);
  xnor csa_tree_add_51_79_groupi_g36421(csa_tree_add_51_79_groupi_n_9628 ,csa_tree_add_51_79_groupi_n_9271 ,csa_tree_add_51_79_groupi_n_9385);
  xnor csa_tree_add_51_79_groupi_g36422(csa_tree_add_51_79_groupi_n_9627 ,csa_tree_add_51_79_groupi_n_9255 ,csa_tree_add_51_79_groupi_n_8966);
  xnor csa_tree_add_51_79_groupi_g36423(csa_tree_add_51_79_groupi_n_9626 ,csa_tree_add_51_79_groupi_n_9252 ,csa_tree_add_51_79_groupi_n_9291);
  xnor csa_tree_add_51_79_groupi_g36424(csa_tree_add_51_79_groupi_n_9625 ,csa_tree_add_51_79_groupi_n_9299 ,csa_tree_add_51_79_groupi_n_8733);
  xnor csa_tree_add_51_79_groupi_g36425(csa_tree_add_51_79_groupi_n_9624 ,csa_tree_add_51_79_groupi_n_9069 ,csa_tree_add_51_79_groupi_n_9357);
  xnor csa_tree_add_51_79_groupi_g36426(csa_tree_add_51_79_groupi_n_9623 ,csa_tree_add_51_79_groupi_n_9374 ,csa_tree_add_51_79_groupi_n_9382);
  xnor csa_tree_add_51_79_groupi_g36427(csa_tree_add_51_79_groupi_n_9622 ,csa_tree_add_51_79_groupi_n_9370 ,csa_tree_add_51_79_groupi_n_9265);
  xnor csa_tree_add_51_79_groupi_g36428(csa_tree_add_51_79_groupi_n_9621 ,csa_tree_add_51_79_groupi_n_9254 ,csa_tree_add_51_79_groupi_n_9270);
  xnor csa_tree_add_51_79_groupi_g36429(csa_tree_add_51_79_groupi_n_9620 ,csa_tree_add_51_79_groupi_n_9290 ,csa_tree_add_51_79_groupi_n_8761);
  xnor csa_tree_add_51_79_groupi_g36430(csa_tree_add_51_79_groupi_n_9619 ,csa_tree_add_51_79_groupi_n_9289 ,csa_tree_add_51_79_groupi_n_9256);
  xnor csa_tree_add_51_79_groupi_g36431(csa_tree_add_51_79_groupi_n_9618 ,csa_tree_add_51_79_groupi_n_9267 ,csa_tree_add_51_79_groupi_n_9083);
  xnor csa_tree_add_51_79_groupi_g36432(csa_tree_add_51_79_groupi_n_9617 ,csa_tree_add_51_79_groupi_n_9383 ,csa_tree_add_51_79_groupi_n_9381);
  xnor csa_tree_add_51_79_groupi_g36433(csa_tree_add_51_79_groupi_n_9616 ,csa_tree_add_51_79_groupi_n_9287 ,csa_tree_add_51_79_groupi_n_9263);
  xnor csa_tree_add_51_79_groupi_g36434(csa_tree_add_51_79_groupi_n_9615 ,csa_tree_add_51_79_groupi_n_9392 ,csa_tree_add_51_79_groupi_n_9361);
  xnor csa_tree_add_51_79_groupi_g36435(csa_tree_add_51_79_groupi_n_9708 ,csa_tree_add_51_79_groupi_n_8792 ,csa_tree_add_51_79_groupi_n_9219);
  xnor csa_tree_add_51_79_groupi_g36436(csa_tree_add_51_79_groupi_n_9707 ,csa_tree_add_51_79_groupi_n_8423 ,csa_tree_add_51_79_groupi_n_9210);
  xnor csa_tree_add_51_79_groupi_g36437(csa_tree_add_51_79_groupi_n_9706 ,csa_tree_add_51_79_groupi_n_8964 ,csa_tree_add_51_79_groupi_n_9209);
  xnor csa_tree_add_51_79_groupi_g36438(csa_tree_add_51_79_groupi_n_9705 ,csa_tree_add_51_79_groupi_n_8823 ,csa_tree_add_51_79_groupi_n_9233);
  xnor csa_tree_add_51_79_groupi_g36439(csa_tree_add_51_79_groupi_n_9704 ,csa_tree_add_51_79_groupi_n_8798 ,csa_tree_add_51_79_groupi_n_9216);
  xnor csa_tree_add_51_79_groupi_g36440(csa_tree_add_51_79_groupi_n_9703 ,csa_tree_add_51_79_groupi_n_9399 ,csa_tree_add_51_79_groupi_n_9232);
  xnor csa_tree_add_51_79_groupi_g36441(csa_tree_add_51_79_groupi_n_9702 ,csa_tree_add_51_79_groupi_n_8785 ,csa_tree_add_51_79_groupi_n_9234);
  xnor csa_tree_add_51_79_groupi_g36442(csa_tree_add_51_79_groupi_n_9701 ,csa_tree_add_51_79_groupi_n_8784 ,csa_tree_add_51_79_groupi_n_9223);
  xnor csa_tree_add_51_79_groupi_g36443(csa_tree_add_51_79_groupi_n_9700 ,csa_tree_add_51_79_groupi_n_8804 ,csa_tree_add_51_79_groupi_n_9221);
  xnor csa_tree_add_51_79_groupi_g36444(csa_tree_add_51_79_groupi_n_9699 ,csa_tree_add_51_79_groupi_n_8796 ,csa_tree_add_51_79_groupi_n_9227);
  xnor csa_tree_add_51_79_groupi_g36445(csa_tree_add_51_79_groupi_n_9698 ,csa_tree_add_51_79_groupi_n_9204 ,csa_tree_add_51_79_groupi_n_9236);
  xnor csa_tree_add_51_79_groupi_g36446(csa_tree_add_51_79_groupi_n_9697 ,csa_tree_add_51_79_groupi_n_8758 ,csa_tree_add_51_79_groupi_n_9225);
  xnor csa_tree_add_51_79_groupi_g36447(csa_tree_add_51_79_groupi_n_9696 ,csa_tree_add_51_79_groupi_n_8802 ,csa_tree_add_51_79_groupi_n_9231);
  xnor csa_tree_add_51_79_groupi_g36448(csa_tree_add_51_79_groupi_n_9695 ,csa_tree_add_51_79_groupi_n_9198 ,csa_tree_add_51_79_groupi_n_9228);
  and csa_tree_add_51_79_groupi_g36449(csa_tree_add_51_79_groupi_n_9694 ,csa_tree_add_51_79_groupi_n_9243 ,csa_tree_add_51_79_groupi_n_9425);
  xnor csa_tree_add_51_79_groupi_g36450(csa_tree_add_51_79_groupi_n_9693 ,csa_tree_add_51_79_groupi_n_8772 ,csa_tree_add_51_79_groupi_n_9213);
  xnor csa_tree_add_51_79_groupi_g36451(csa_tree_add_51_79_groupi_n_9692 ,csa_tree_add_51_79_groupi_n_8803 ,csa_tree_add_51_79_groupi_n_9208);
  xnor csa_tree_add_51_79_groupi_g36452(csa_tree_add_51_79_groupi_n_9691 ,csa_tree_add_51_79_groupi_n_8642 ,csa_tree_add_51_79_groupi_n_9222);
  xnor csa_tree_add_51_79_groupi_g36453(csa_tree_add_51_79_groupi_n_9690 ,csa_tree_add_51_79_groupi_n_8723 ,csa_tree_add_51_79_groupi_n_9229);
  xnor csa_tree_add_51_79_groupi_g36454(csa_tree_add_51_79_groupi_n_9689 ,csa_tree_add_51_79_groupi_n_8817 ,csa_tree_add_51_79_groupi_n_9226);
  xnor csa_tree_add_51_79_groupi_g36455(csa_tree_add_51_79_groupi_n_9687 ,csa_tree_add_51_79_groupi_n_8479 ,csa_tree_add_51_79_groupi_n_9215);
  xnor csa_tree_add_51_79_groupi_g36456(csa_tree_add_51_79_groupi_n_9686 ,csa_tree_add_51_79_groupi_n_8780 ,csa_tree_add_51_79_groupi_n_9207);
  and csa_tree_add_51_79_groupi_g36457(csa_tree_add_51_79_groupi_n_9685 ,csa_tree_add_51_79_groupi_n_9240 ,csa_tree_add_51_79_groupi_n_9424);
  xnor csa_tree_add_51_79_groupi_g36458(csa_tree_add_51_79_groupi_n_9684 ,csa_tree_add_51_79_groupi_n_8726 ,csa_tree_add_51_79_groupi_n_9235);
  xnor csa_tree_add_51_79_groupi_g36459(csa_tree_add_51_79_groupi_n_9683 ,csa_tree_add_51_79_groupi_n_9201 ,csa_tree_add_51_79_groupi_n_9217);
  xnor csa_tree_add_51_79_groupi_g36460(csa_tree_add_51_79_groupi_n_9682 ,csa_tree_add_51_79_groupi_n_8764 ,csa_tree_add_51_79_groupi_n_9212);
  xnor csa_tree_add_51_79_groupi_g36461(csa_tree_add_51_79_groupi_n_9681 ,csa_tree_add_51_79_groupi_n_8728 ,csa_tree_add_51_79_groupi_n_9230);
  xnor csa_tree_add_51_79_groupi_g36462(csa_tree_add_51_79_groupi_n_9680 ,csa_tree_add_51_79_groupi_n_8756 ,csa_tree_add_51_79_groupi_n_9211);
  xnor csa_tree_add_51_79_groupi_g36463(csa_tree_add_51_79_groupi_n_9678 ,csa_tree_add_51_79_groupi_n_8960 ,csa_tree_add_51_79_groupi_n_9220);
  xnor csa_tree_add_51_79_groupi_g36464(csa_tree_add_51_79_groupi_n_9677 ,csa_tree_add_51_79_groupi_n_8743 ,csa_tree_add_51_79_groupi_n_9218);
  xnor csa_tree_add_51_79_groupi_g36465(csa_tree_add_51_79_groupi_n_9676 ,csa_tree_add_51_79_groupi_n_9262 ,csa_tree_add_51_79_groupi_n_9214);
  xor csa_tree_add_51_79_groupi_g36466(csa_tree_add_51_79_groupi_n_9674 ,csa_tree_add_51_79_groupi_n_8738 ,csa_tree_add_51_79_groupi_n_9224);
  not csa_tree_add_51_79_groupi_g36468(csa_tree_add_51_79_groupi_n_9605 ,csa_tree_add_51_79_groupi_n_9604);
  not csa_tree_add_51_79_groupi_g36469(csa_tree_add_51_79_groupi_n_9593 ,csa_tree_add_51_79_groupi_n_9594);
  not csa_tree_add_51_79_groupi_g36470(csa_tree_add_51_79_groupi_n_9591 ,csa_tree_add_51_79_groupi_n_9590);
  not csa_tree_add_51_79_groupi_g36471(csa_tree_add_51_79_groupi_n_9584 ,csa_tree_add_51_79_groupi_n_9583);
  and csa_tree_add_51_79_groupi_g36472(csa_tree_add_51_79_groupi_n_9580 ,csa_tree_add_51_79_groupi_n_9369 ,csa_tree_add_51_79_groupi_n_9249);
  or csa_tree_add_51_79_groupi_g36473(csa_tree_add_51_79_groupi_n_9579 ,csa_tree_add_51_79_groupi_n_9251 ,csa_tree_add_51_79_groupi_n_9285);
  or csa_tree_add_51_79_groupi_g36474(csa_tree_add_51_79_groupi_n_9578 ,csa_tree_add_51_79_groupi_n_9099 ,csa_tree_add_51_79_groupi_n_9304);
  or csa_tree_add_51_79_groupi_g36475(csa_tree_add_51_79_groupi_n_9577 ,csa_tree_add_51_79_groupi_n_8152 ,csa_tree_add_51_79_groupi_n_9262);
  nor csa_tree_add_51_79_groupi_g36476(csa_tree_add_51_79_groupi_n_9576 ,csa_tree_add_51_79_groupi_n_8635 ,csa_tree_add_51_79_groupi_n_9246);
  nor csa_tree_add_51_79_groupi_g36477(csa_tree_add_51_79_groupi_n_9575 ,csa_tree_add_51_79_groupi_n_8810 ,csa_tree_add_51_79_groupi_n_9244);
  nor csa_tree_add_51_79_groupi_g36478(csa_tree_add_51_79_groupi_n_9574 ,csa_tree_add_51_79_groupi_n_9183 ,csa_tree_add_51_79_groupi_n_9278);
  or csa_tree_add_51_79_groupi_g36479(csa_tree_add_51_79_groupi_n_9573 ,csa_tree_add_51_79_groupi_n_9359 ,csa_tree_add_51_79_groupi_n_9367);
  and csa_tree_add_51_79_groupi_g36480(csa_tree_add_51_79_groupi_n_9572 ,csa_tree_add_51_79_groupi_n_9348 ,csa_tree_add_51_79_groupi_n_9085);
  or csa_tree_add_51_79_groupi_g36481(csa_tree_add_51_79_groupi_n_9571 ,csa_tree_add_51_79_groupi_n_9261 ,csa_tree_add_51_79_groupi_n_9280);
  nor csa_tree_add_51_79_groupi_g36482(csa_tree_add_51_79_groupi_n_9570 ,csa_tree_add_51_79_groupi_n_9260 ,csa_tree_add_51_79_groupi_n_9281);
  and csa_tree_add_51_79_groupi_g36483(csa_tree_add_51_79_groupi_n_9569 ,csa_tree_add_51_79_groupi_n_9363 ,csa_tree_add_51_79_groupi_n_9362);
  or csa_tree_add_51_79_groupi_g36484(csa_tree_add_51_79_groupi_n_9568 ,csa_tree_add_51_79_groupi_n_8795 ,csa_tree_add_51_79_groupi_n_9347);
  or csa_tree_add_51_79_groupi_g36485(csa_tree_add_51_79_groupi_n_9567 ,csa_tree_add_51_79_groupi_n_9345 ,csa_tree_add_51_79_groupi_n_9401);
  or csa_tree_add_51_79_groupi_g36486(csa_tree_add_51_79_groupi_n_9566 ,csa_tree_add_51_79_groupi_n_9264 ,csa_tree_add_51_79_groupi_n_9361);
  or csa_tree_add_51_79_groupi_g36487(csa_tree_add_51_79_groupi_n_9565 ,csa_tree_add_51_79_groupi_n_9363 ,csa_tree_add_51_79_groupi_n_9362);
  and csa_tree_add_51_79_groupi_g36488(csa_tree_add_51_79_groupi_n_9564 ,csa_tree_add_51_79_groupi_n_9264 ,csa_tree_add_51_79_groupi_n_9361);
  or csa_tree_add_51_79_groupi_g36489(csa_tree_add_51_79_groupi_n_9563 ,csa_tree_add_51_79_groupi_n_9263 ,csa_tree_add_51_79_groupi_n_9287);
  and csa_tree_add_51_79_groupi_g36490(csa_tree_add_51_79_groupi_n_9562 ,csa_tree_add_51_79_groupi_n_9263 ,csa_tree_add_51_79_groupi_n_9287);
  or csa_tree_add_51_79_groupi_g36491(csa_tree_add_51_79_groupi_n_9561 ,csa_tree_add_51_79_groupi_n_9366 ,csa_tree_add_51_79_groupi_n_9259);
  and csa_tree_add_51_79_groupi_g36492(csa_tree_add_51_79_groupi_n_9560 ,csa_tree_add_51_79_groupi_n_9366 ,csa_tree_add_51_79_groupi_n_9259);
  or csa_tree_add_51_79_groupi_g36493(csa_tree_add_51_79_groupi_n_9559 ,csa_tree_add_51_79_groupi_n_9382 ,csa_tree_add_51_79_groupi_n_9374);
  and csa_tree_add_51_79_groupi_g36494(csa_tree_add_51_79_groupi_n_9558 ,csa_tree_add_51_79_groupi_n_8152 ,csa_tree_add_51_79_groupi_n_9262);
  and csa_tree_add_51_79_groupi_g36495(csa_tree_add_51_79_groupi_n_9557 ,csa_tree_add_51_79_groupi_n_9382 ,csa_tree_add_51_79_groupi_n_9374);
  and csa_tree_add_51_79_groupi_g36496(csa_tree_add_51_79_groupi_n_9556 ,csa_tree_add_51_79_groupi_n_9359 ,csa_tree_add_51_79_groupi_n_9367);
  or csa_tree_add_51_79_groupi_g36497(csa_tree_add_51_79_groupi_n_9555 ,csa_tree_add_51_79_groupi_n_9298 ,csa_tree_add_51_79_groupi_n_9342);
  and csa_tree_add_51_79_groupi_g36498(csa_tree_add_51_79_groupi_n_9554 ,csa_tree_add_51_79_groupi_n_9188 ,csa_tree_add_51_79_groupi_n_9286);
  or csa_tree_add_51_79_groupi_g36499(csa_tree_add_51_79_groupi_n_9553 ,csa_tree_add_51_79_groupi_n_9188 ,csa_tree_add_51_79_groupi_n_9286);
  or csa_tree_add_51_79_groupi_g36500(csa_tree_add_51_79_groupi_n_9552 ,csa_tree_add_51_79_groupi_n_9266 ,csa_tree_add_51_79_groupi_n_9257);
  or csa_tree_add_51_79_groupi_g36501(csa_tree_add_51_79_groupi_n_9551 ,csa_tree_add_51_79_groupi_n_9256 ,csa_tree_add_51_79_groupi_n_9289);
  and csa_tree_add_51_79_groupi_g36502(csa_tree_add_51_79_groupi_n_9550 ,csa_tree_add_51_79_groupi_n_9256 ,csa_tree_add_51_79_groupi_n_9289);
  nor csa_tree_add_51_79_groupi_g36503(csa_tree_add_51_79_groupi_n_9549 ,csa_tree_add_51_79_groupi_n_9202 ,csa_tree_add_51_79_groupi_n_9326);
  or csa_tree_add_51_79_groupi_g36504(csa_tree_add_51_79_groupi_n_9548 ,csa_tree_add_51_79_groupi_n_9203 ,csa_tree_add_51_79_groupi_n_9333);
  and csa_tree_add_51_79_groupi_g36505(csa_tree_add_51_79_groupi_n_9547 ,csa_tree_add_51_79_groupi_n_9266 ,csa_tree_add_51_79_groupi_n_9257);
  and csa_tree_add_51_79_groupi_g36506(csa_tree_add_51_79_groupi_n_9546 ,csa_tree_add_51_79_groupi_n_9381 ,csa_tree_add_51_79_groupi_n_9250);
  or csa_tree_add_51_79_groupi_g36507(csa_tree_add_51_79_groupi_n_9545 ,csa_tree_add_51_79_groupi_n_9193 ,csa_tree_add_51_79_groupi_n_9274);
  or csa_tree_add_51_79_groupi_g36508(csa_tree_add_51_79_groupi_n_9544 ,csa_tree_add_51_79_groupi_n_9195 ,csa_tree_add_51_79_groupi_n_9268);
  or csa_tree_add_51_79_groupi_g36509(csa_tree_add_51_79_groupi_n_9543 ,csa_tree_add_51_79_groupi_n_9282 ,csa_tree_add_51_79_groupi_n_9378);
  and csa_tree_add_51_79_groupi_g36510(csa_tree_add_51_79_groupi_n_9542 ,csa_tree_add_51_79_groupi_n_9282 ,csa_tree_add_51_79_groupi_n_9378);
  or csa_tree_add_51_79_groupi_g36511(csa_tree_add_51_79_groupi_n_9541 ,csa_tree_add_51_79_groupi_n_8733 ,csa_tree_add_51_79_groupi_n_9373);
  or csa_tree_add_51_79_groupi_g36512(csa_tree_add_51_79_groupi_n_9540 ,csa_tree_add_51_79_groupi_n_8970 ,csa_tree_add_51_79_groupi_n_9317);
  and csa_tree_add_51_79_groupi_g36513(csa_tree_add_51_79_groupi_n_9539 ,csa_tree_add_51_79_groupi_n_8733 ,csa_tree_add_51_79_groupi_n_9373);
  or csa_tree_add_51_79_groupi_g36514(csa_tree_add_51_79_groupi_n_9538 ,csa_tree_add_51_79_groupi_n_9369 ,csa_tree_add_51_79_groupi_n_9249);
  or csa_tree_add_51_79_groupi_g36515(csa_tree_add_51_79_groupi_n_9537 ,csa_tree_add_51_79_groupi_n_8805 ,csa_tree_add_51_79_groupi_n_9312);
  or csa_tree_add_51_79_groupi_g36516(csa_tree_add_51_79_groupi_n_9536 ,csa_tree_add_51_79_groupi_n_9364 ,csa_tree_add_51_79_groupi_n_9356);
  and csa_tree_add_51_79_groupi_g36517(csa_tree_add_51_79_groupi_n_9535 ,csa_tree_add_51_79_groupi_n_9394 ,csa_tree_add_51_79_groupi_n_9238);
  nor csa_tree_add_51_79_groupi_g36518(csa_tree_add_51_79_groupi_n_9534 ,csa_tree_add_51_79_groupi_n_9192 ,csa_tree_add_51_79_groupi_n_9275);
  or csa_tree_add_51_79_groupi_g36519(csa_tree_add_51_79_groupi_n_9533 ,csa_tree_add_51_79_groupi_n_9271 ,csa_tree_add_51_79_groupi_n_9360);
  nor csa_tree_add_51_79_groupi_g36520(csa_tree_add_51_79_groupi_n_9532 ,csa_tree_add_51_79_groupi_n_9365 ,csa_tree_add_51_79_groupi_n_9355);
  or csa_tree_add_51_79_groupi_g36521(csa_tree_add_51_79_groupi_n_9531 ,csa_tree_add_51_79_groupi_n_9381 ,csa_tree_add_51_79_groupi_n_9250);
  and csa_tree_add_51_79_groupi_g36522(csa_tree_add_51_79_groupi_n_9530 ,csa_tree_add_51_79_groupi_n_9190 ,csa_tree_add_51_79_groupi_n_9294);
  or csa_tree_add_51_79_groupi_g36523(csa_tree_add_51_79_groupi_n_9529 ,csa_tree_add_51_79_groupi_n_9254 ,csa_tree_add_51_79_groupi_n_9269);
  and csa_tree_add_51_79_groupi_g36524(csa_tree_add_51_79_groupi_n_9528 ,csa_tree_add_51_79_groupi_n_9271 ,csa_tree_add_51_79_groupi_n_9360);
  or csa_tree_add_51_79_groupi_g36525(csa_tree_add_51_79_groupi_n_9527 ,csa_tree_add_51_79_groupi_n_9399 ,csa_tree_add_51_79_groupi_n_9059);
  nor csa_tree_add_51_79_groupi_g36526(csa_tree_add_51_79_groupi_n_9526 ,csa_tree_add_51_79_groupi_n_9253 ,csa_tree_add_51_79_groupi_n_9270);
  or csa_tree_add_51_79_groupi_g36527(csa_tree_add_51_79_groupi_n_9525 ,csa_tree_add_51_79_groupi_n_9182 ,csa_tree_add_51_79_groupi_n_9277);
  or csa_tree_add_51_79_groupi_g36528(csa_tree_add_51_79_groupi_n_9524 ,csa_tree_add_51_79_groupi_n_9184 ,csa_tree_add_51_79_groupi_n_9371);
  or csa_tree_add_51_79_groupi_g36529(csa_tree_add_51_79_groupi_n_9523 ,csa_tree_add_51_79_groupi_n_9265 ,csa_tree_add_51_79_groupi_n_9370);
  and csa_tree_add_51_79_groupi_g36530(csa_tree_add_51_79_groupi_n_9522 ,csa_tree_add_51_79_groupi_n_9265 ,csa_tree_add_51_79_groupi_n_9370);
  and csa_tree_add_51_79_groupi_g36531(csa_tree_add_51_79_groupi_n_9521 ,csa_tree_add_51_79_groupi_n_9191 ,csa_tree_add_51_79_groupi_n_9377);
  nor csa_tree_add_51_79_groupi_g36532(csa_tree_add_51_79_groupi_n_9520 ,csa_tree_add_51_79_groupi_n_9185 ,csa_tree_add_51_79_groupi_n_9372);
  and csa_tree_add_51_79_groupi_g36533(csa_tree_add_51_79_groupi_n_9519 ,csa_tree_add_51_79_groupi_n_9195 ,csa_tree_add_51_79_groupi_n_9268);
  or csa_tree_add_51_79_groupi_g36534(csa_tree_add_51_79_groupi_n_9518 ,csa_tree_add_51_79_groupi_n_9191 ,csa_tree_add_51_79_groupi_n_9377);
  or csa_tree_add_51_79_groupi_g36535(csa_tree_add_51_79_groupi_n_9517 ,csa_tree_add_51_79_groupi_n_9190 ,csa_tree_add_51_79_groupi_n_9294);
  and csa_tree_add_51_79_groupi_g36536(csa_tree_add_51_79_groupi_n_9614 ,csa_tree_add_51_79_groupi_n_9158 ,csa_tree_add_51_79_groupi_n_9335);
  and csa_tree_add_51_79_groupi_g36537(csa_tree_add_51_79_groupi_n_9613 ,csa_tree_add_51_79_groupi_n_9107 ,csa_tree_add_51_79_groupi_n_9316);
  and csa_tree_add_51_79_groupi_g36538(csa_tree_add_51_79_groupi_n_9612 ,csa_tree_add_51_79_groupi_n_9108 ,csa_tree_add_51_79_groupi_n_9315);
  and csa_tree_add_51_79_groupi_g36539(csa_tree_add_51_79_groupi_n_9611 ,csa_tree_add_51_79_groupi_n_9100 ,csa_tree_add_51_79_groupi_n_9324);
  and csa_tree_add_51_79_groupi_g36540(csa_tree_add_51_79_groupi_n_9610 ,csa_tree_add_51_79_groupi_n_9116 ,csa_tree_add_51_79_groupi_n_9310);
  and csa_tree_add_51_79_groupi_g36541(csa_tree_add_51_79_groupi_n_9609 ,csa_tree_add_51_79_groupi_n_9119 ,csa_tree_add_51_79_groupi_n_9354);
  and csa_tree_add_51_79_groupi_g36542(csa_tree_add_51_79_groupi_n_9608 ,csa_tree_add_51_79_groupi_n_9132 ,csa_tree_add_51_79_groupi_n_9334);
  and csa_tree_add_51_79_groupi_g36543(csa_tree_add_51_79_groupi_n_9607 ,csa_tree_add_51_79_groupi_n_9136 ,csa_tree_add_51_79_groupi_n_9325);
  and csa_tree_add_51_79_groupi_g36544(csa_tree_add_51_79_groupi_n_9606 ,csa_tree_add_51_79_groupi_n_9144 ,csa_tree_add_51_79_groupi_n_9328);
  or csa_tree_add_51_79_groupi_g36545(csa_tree_add_51_79_groupi_n_9604 ,csa_tree_add_51_79_groupi_n_9097 ,csa_tree_add_51_79_groupi_n_9319);
  and csa_tree_add_51_79_groupi_g36546(csa_tree_add_51_79_groupi_n_9603 ,csa_tree_add_51_79_groupi_n_9173 ,csa_tree_add_51_79_groupi_n_9336);
  and csa_tree_add_51_79_groupi_g36547(csa_tree_add_51_79_groupi_n_9602 ,csa_tree_add_51_79_groupi_n_9066 ,csa_tree_add_51_79_groupi_n_9337);
  and csa_tree_add_51_79_groupi_g36548(csa_tree_add_51_79_groupi_n_9601 ,csa_tree_add_51_79_groupi_n_9064 ,csa_tree_add_51_79_groupi_n_9338);
  and csa_tree_add_51_79_groupi_g36549(csa_tree_add_51_79_groupi_n_9600 ,csa_tree_add_51_79_groupi_n_9163 ,csa_tree_add_51_79_groupi_n_9343);
  and csa_tree_add_51_79_groupi_g36550(csa_tree_add_51_79_groupi_n_9599 ,csa_tree_add_51_79_groupi_n_9056 ,csa_tree_add_51_79_groupi_n_9349);
  and csa_tree_add_51_79_groupi_g36551(csa_tree_add_51_79_groupi_n_9598 ,csa_tree_add_51_79_groupi_n_9048 ,csa_tree_add_51_79_groupi_n_9242);
  and csa_tree_add_51_79_groupi_g36552(csa_tree_add_51_79_groupi_n_9597 ,csa_tree_add_51_79_groupi_n_9090 ,csa_tree_add_51_79_groupi_n_9321);
  and csa_tree_add_51_79_groupi_g36553(csa_tree_add_51_79_groupi_n_9596 ,csa_tree_add_51_79_groupi_n_9141 ,csa_tree_add_51_79_groupi_n_9352);
  or csa_tree_add_51_79_groupi_g36554(csa_tree_add_51_79_groupi_n_9595 ,csa_tree_add_51_79_groupi_n_9087 ,csa_tree_add_51_79_groupi_n_9323);
  or csa_tree_add_51_79_groupi_g36555(csa_tree_add_51_79_groupi_n_9594 ,csa_tree_add_51_79_groupi_n_9145 ,csa_tree_add_51_79_groupi_n_9331);
  and csa_tree_add_51_79_groupi_g36556(csa_tree_add_51_79_groupi_n_9592 ,csa_tree_add_51_79_groupi_n_9159 ,csa_tree_add_51_79_groupi_n_9341);
  or csa_tree_add_51_79_groupi_g36557(csa_tree_add_51_79_groupi_n_9590 ,csa_tree_add_51_79_groupi_n_9088 ,csa_tree_add_51_79_groupi_n_9327);
  and csa_tree_add_51_79_groupi_g36558(csa_tree_add_51_79_groupi_n_9589 ,csa_tree_add_51_79_groupi_n_9043 ,csa_tree_add_51_79_groupi_n_9318);
  and csa_tree_add_51_79_groupi_g36559(csa_tree_add_51_79_groupi_n_9588 ,csa_tree_add_51_79_groupi_n_9054 ,csa_tree_add_51_79_groupi_n_9237);
  and csa_tree_add_51_79_groupi_g36560(csa_tree_add_51_79_groupi_n_9587 ,csa_tree_add_51_79_groupi_n_8955 ,csa_tree_add_51_79_groupi_n_9309);
  or csa_tree_add_51_79_groupi_g36561(csa_tree_add_51_79_groupi_n_9586 ,csa_tree_add_51_79_groupi_n_9166 ,csa_tree_add_51_79_groupi_n_9346);
  and csa_tree_add_51_79_groupi_g36562(csa_tree_add_51_79_groupi_n_9585 ,csa_tree_add_51_79_groupi_n_9170 ,csa_tree_add_51_79_groupi_n_9351);
  or csa_tree_add_51_79_groupi_g36563(csa_tree_add_51_79_groupi_n_9583 ,csa_tree_add_51_79_groupi_n_9124 ,csa_tree_add_51_79_groupi_n_9313);
  and csa_tree_add_51_79_groupi_g36564(csa_tree_add_51_79_groupi_n_9582 ,csa_tree_add_51_79_groupi_n_9062 ,csa_tree_add_51_79_groupi_n_9339);
  and csa_tree_add_51_79_groupi_g36565(csa_tree_add_51_79_groupi_n_9581 ,csa_tree_add_51_79_groupi_n_9171 ,csa_tree_add_51_79_groupi_n_9330);
  not csa_tree_add_51_79_groupi_g36566(csa_tree_add_51_79_groupi_n_9513 ,csa_tree_add_51_79_groupi_n_9512);
  not csa_tree_add_51_79_groupi_g36567(csa_tree_add_51_79_groupi_n_9511 ,csa_tree_add_51_79_groupi_n_9510);
  not csa_tree_add_51_79_groupi_g36568(csa_tree_add_51_79_groupi_n_9508 ,csa_tree_add_51_79_groupi_n_9507);
  not csa_tree_add_51_79_groupi_g36569(csa_tree_add_51_79_groupi_n_9503 ,csa_tree_add_51_79_groupi_n_9504);
  not csa_tree_add_51_79_groupi_g36570(csa_tree_add_51_79_groupi_n_9501 ,csa_tree_add_51_79_groupi_n_9502);
  not csa_tree_add_51_79_groupi_g36571(csa_tree_add_51_79_groupi_n_9499 ,csa_tree_add_51_79_groupi_n_9500);
  not csa_tree_add_51_79_groupi_g36572(csa_tree_add_51_79_groupi_n_9498 ,csa_tree_add_51_79_groupi_n_9497);
  not csa_tree_add_51_79_groupi_g36573(csa_tree_add_51_79_groupi_n_9495 ,csa_tree_add_51_79_groupi_n_9494);
  not csa_tree_add_51_79_groupi_g36574(csa_tree_add_51_79_groupi_n_9493 ,csa_tree_add_51_79_groupi_n_9492);
  not csa_tree_add_51_79_groupi_g36575(csa_tree_add_51_79_groupi_n_9491 ,csa_tree_add_51_79_groupi_n_9490);
  not csa_tree_add_51_79_groupi_g36576(csa_tree_add_51_79_groupi_n_9488 ,csa_tree_add_51_79_groupi_n_9487);
  not csa_tree_add_51_79_groupi_g36577(csa_tree_add_51_79_groupi_n_9485 ,csa_tree_add_51_79_groupi_n_9484);
  not csa_tree_add_51_79_groupi_g36578(csa_tree_add_51_79_groupi_n_9474 ,csa_tree_add_51_79_groupi_n_9473);
  not csa_tree_add_51_79_groupi_g36579(csa_tree_add_51_79_groupi_n_9468 ,csa_tree_add_51_79_groupi_n_9469);
  not csa_tree_add_51_79_groupi_g36580(csa_tree_add_51_79_groupi_n_9467 ,csa_tree_add_51_79_groupi_n_9466);
  not csa_tree_add_51_79_groupi_g36581(csa_tree_add_51_79_groupi_n_9453 ,csa_tree_add_51_79_groupi_n_9452);
  not csa_tree_add_51_79_groupi_g36582(csa_tree_add_51_79_groupi_n_9448 ,csa_tree_add_51_79_groupi_n_9449);
  not csa_tree_add_51_79_groupi_g36583(csa_tree_add_51_79_groupi_n_9446 ,csa_tree_add_51_79_groupi_n_9445);
  not csa_tree_add_51_79_groupi_g36584(csa_tree_add_51_79_groupi_n_9443 ,csa_tree_add_51_79_groupi_n_9444);
  and csa_tree_add_51_79_groupi_g36585(csa_tree_add_51_79_groupi_n_9437 ,csa_tree_add_51_79_groupi_n_9251 ,csa_tree_add_51_79_groupi_n_9285);
  or csa_tree_add_51_79_groupi_g36586(csa_tree_add_51_79_groupi_n_9436 ,csa_tree_add_51_79_groupi_n_9320 ,csa_tree_add_51_79_groupi_n_8967);
  or csa_tree_add_51_79_groupi_g36587(csa_tree_add_51_79_groupi_n_9435 ,csa_tree_add_51_79_groupi_n_9255 ,csa_tree_add_51_79_groupi_n_9283);
  and csa_tree_add_51_79_groupi_g36588(csa_tree_add_51_79_groupi_n_9434 ,csa_tree_add_51_79_groupi_n_9255 ,csa_tree_add_51_79_groupi_n_9283);
  or csa_tree_add_51_79_groupi_g36589(csa_tree_add_51_79_groupi_n_9433 ,csa_tree_add_51_79_groupi_n_8761 ,csa_tree_add_51_79_groupi_n_9290);
  and csa_tree_add_51_79_groupi_g36590(csa_tree_add_51_79_groupi_n_9432 ,csa_tree_add_51_79_groupi_n_8761 ,csa_tree_add_51_79_groupi_n_9290);
  or csa_tree_add_51_79_groupi_g36591(csa_tree_add_51_79_groupi_n_9431 ,csa_tree_add_51_79_groupi_n_9083 ,csa_tree_add_51_79_groupi_n_9267);
  and csa_tree_add_51_79_groupi_g36592(csa_tree_add_51_79_groupi_n_9430 ,csa_tree_add_51_79_groupi_n_9083 ,csa_tree_add_51_79_groupi_n_9267);
  or csa_tree_add_51_79_groupi_g36593(csa_tree_add_51_79_groupi_n_9429 ,csa_tree_add_51_79_groupi_n_9284 ,csa_tree_add_51_79_groupi_n_9258);
  and csa_tree_add_51_79_groupi_g36594(csa_tree_add_51_79_groupi_n_9428 ,csa_tree_add_51_79_groupi_n_9284 ,csa_tree_add_51_79_groupi_n_9258);
  or csa_tree_add_51_79_groupi_g36595(csa_tree_add_51_79_groupi_n_9427 ,csa_tree_add_51_79_groupi_n_9291 ,csa_tree_add_51_79_groupi_n_9252);
  and csa_tree_add_51_79_groupi_g36596(csa_tree_add_51_79_groupi_n_9426 ,csa_tree_add_51_79_groupi_n_9291 ,csa_tree_add_51_79_groupi_n_9252);
  or csa_tree_add_51_79_groupi_g36597(csa_tree_add_51_79_groupi_n_9425 ,csa_tree_add_51_79_groupi_n_8806 ,csa_tree_add_51_79_groupi_n_9248);
  or csa_tree_add_51_79_groupi_g36598(csa_tree_add_51_79_groupi_n_9424 ,csa_tree_add_51_79_groupi_n_9206 ,csa_tree_add_51_79_groupi_n_9241);
  and csa_tree_add_51_79_groupi_g36599(csa_tree_add_51_79_groupi_n_9423 ,csa_tree_add_51_79_groupi_n_9368 ,csa_tree_add_51_79_groupi_n_9288);
  nor csa_tree_add_51_79_groupi_g36600(csa_tree_add_51_79_groupi_n_9422 ,csa_tree_add_51_79_groupi_n_9368 ,csa_tree_add_51_79_groupi_n_9288);
  or csa_tree_add_51_79_groupi_g36601(csa_tree_add_51_79_groupi_n_9421 ,csa_tree_add_51_79_groupi_n_9069 ,csa_tree_add_51_79_groupi_n_9357);
  and csa_tree_add_51_79_groupi_g36602(csa_tree_add_51_79_groupi_n_9420 ,csa_tree_add_51_79_groupi_n_9069 ,csa_tree_add_51_79_groupi_n_9357);
  xnor csa_tree_add_51_79_groupi_g36603(csa_tree_add_51_79_groupi_n_9419 ,csa_tree_add_51_79_groupi_n_9180 ,csa_tree_add_51_79_groupi_n_9179);
  xnor csa_tree_add_51_79_groupi_g36604(csa_tree_add_51_79_groupi_n_9418 ,csa_tree_add_51_79_groupi_n_8806 ,csa_tree_add_51_79_groupi_n_9070);
  xnor csa_tree_add_51_79_groupi_g36605(csa_tree_add_51_79_groupi_n_9417 ,csa_tree_add_51_79_groupi_n_8962 ,csa_tree_add_51_79_groupi_n_9175);
  xnor csa_tree_add_51_79_groupi_g36606(csa_tree_add_51_79_groupi_n_9416 ,csa_tree_add_51_79_groupi_n_8963 ,csa_tree_add_51_79_groupi_n_9183);
  xnor csa_tree_add_51_79_groupi_g36607(csa_tree_add_51_79_groupi_n_9415 ,csa_tree_add_51_79_groupi_n_8805 ,csa_tree_add_51_79_groupi_n_9080);
  xnor csa_tree_add_51_79_groupi_g36608(csa_tree_add_51_79_groupi_n_9414 ,csa_tree_add_51_79_groupi_n_9194 ,csa_tree_add_51_79_groupi_n_8970);
  xnor csa_tree_add_51_79_groupi_g36609(csa_tree_add_51_79_groupi_n_9413 ,csa_tree_add_51_79_groupi_n_9077 ,csa_tree_add_51_79_groupi_n_8788);
  xnor csa_tree_add_51_79_groupi_g36610(csa_tree_add_51_79_groupi_n_9412 ,csa_tree_add_51_79_groupi_n_8810 ,csa_tree_add_51_79_groupi_n_9071);
  xnor csa_tree_add_51_79_groupi_g36611(csa_tree_add_51_79_groupi_n_9411 ,csa_tree_add_51_79_groupi_n_7819 ,csa_tree_add_51_79_groupi_n_9178);
  xnor csa_tree_add_51_79_groupi_g36612(csa_tree_add_51_79_groupi_n_9410 ,csa_tree_add_51_79_groupi_n_8747 ,csa_tree_add_51_79_groupi_n_9086);
  xnor csa_tree_add_51_79_groupi_g36613(csa_tree_add_51_79_groupi_n_9409 ,csa_tree_add_51_79_groupi_n_9081 ,csa_tree_add_51_79_groupi_n_8744);
  xnor csa_tree_add_51_79_groupi_g36614(csa_tree_add_51_79_groupi_n_9408 ,csa_tree_add_51_79_groupi_n_9189 ,csa_tree_add_51_79_groupi_n_9072);
  xnor csa_tree_add_51_79_groupi_g36615(csa_tree_add_51_79_groupi_n_9407 ,csa_tree_add_51_79_groupi_n_8791 ,csa_tree_add_51_79_groupi_n_9073);
  xnor csa_tree_add_51_79_groupi_g36616(csa_tree_add_51_79_groupi_n_9406 ,csa_tree_add_51_79_groupi_n_9079 ,csa_tree_add_51_79_groupi_n_8968);
  xnor csa_tree_add_51_79_groupi_g36617(csa_tree_add_51_79_groupi_n_9405 ,csa_tree_add_51_79_groupi_n_9188 ,csa_tree_add_51_79_groupi_n_9205);
  xnor csa_tree_add_51_79_groupi_g36618(csa_tree_add_51_79_groupi_n_9404 ,csa_tree_add_51_79_groupi_n_8614 ,csa_tree_add_51_79_groupi_n_9084);
  xnor csa_tree_add_51_79_groupi_g36619(csa_tree_add_51_79_groupi_n_9516 ,csa_tree_add_51_79_groupi_n_8436 ,csa_tree_add_51_79_groupi_n_8980);
  xnor csa_tree_add_51_79_groupi_g36620(csa_tree_add_51_79_groupi_n_9515 ,csa_tree_add_51_79_groupi_n_8634 ,csa_tree_add_51_79_groupi_n_8972);
  xnor csa_tree_add_51_79_groupi_g36621(csa_tree_add_51_79_groupi_n_9514 ,csa_tree_add_51_79_groupi_n_8434 ,csa_tree_add_51_79_groupi_n_8985);
  xnor csa_tree_add_51_79_groupi_g36622(csa_tree_add_51_79_groupi_n_9512 ,csa_tree_add_51_79_groupi_n_8470 ,csa_tree_add_51_79_groupi_n_9009);
  xnor csa_tree_add_51_79_groupi_g36623(csa_tree_add_51_79_groupi_n_9510 ,csa_tree_add_51_79_groupi_n_8403 ,csa_tree_add_51_79_groupi_n_8974);
  xnor csa_tree_add_51_79_groupi_g36624(csa_tree_add_51_79_groupi_n_9509 ,csa_tree_add_51_79_groupi_n_8652 ,csa_tree_add_51_79_groupi_n_8991);
  xnor csa_tree_add_51_79_groupi_g36625(csa_tree_add_51_79_groupi_n_9507 ,csa_tree_add_51_79_groupi_n_8178 ,csa_tree_add_51_79_groupi_n_9012);
  xnor csa_tree_add_51_79_groupi_g36626(csa_tree_add_51_79_groupi_n_9506 ,csa_tree_add_51_79_groupi_n_8633 ,csa_tree_add_51_79_groupi_n_9011);
  xnor csa_tree_add_51_79_groupi_g36627(csa_tree_add_51_79_groupi_n_9505 ,csa_tree_add_51_79_groupi_n_8484 ,csa_tree_add_51_79_groupi_n_9010);
  xnor csa_tree_add_51_79_groupi_g36628(csa_tree_add_51_79_groupi_n_9504 ,csa_tree_add_51_79_groupi_n_8398 ,csa_tree_add_51_79_groupi_n_9022);
  xnor csa_tree_add_51_79_groupi_g36629(csa_tree_add_51_79_groupi_n_9502 ,csa_tree_add_51_79_groupi_n_8420 ,csa_tree_add_51_79_groupi_n_8976);
  xnor csa_tree_add_51_79_groupi_g36630(csa_tree_add_51_79_groupi_n_9500 ,csa_tree_add_51_79_groupi_n_8406 ,csa_tree_add_51_79_groupi_n_9029);
  xnor csa_tree_add_51_79_groupi_g36631(csa_tree_add_51_79_groupi_n_9497 ,csa_tree_add_51_79_groupi_n_8628 ,csa_tree_add_51_79_groupi_n_9007);
  xnor csa_tree_add_51_79_groupi_g36632(csa_tree_add_51_79_groupi_n_9496 ,csa_tree_add_51_79_groupi_n_8502 ,csa_tree_add_51_79_groupi_n_9006);
  xnor csa_tree_add_51_79_groupi_g36633(csa_tree_add_51_79_groupi_n_9494 ,csa_tree_add_51_79_groupi_n_8185 ,csa_tree_add_51_79_groupi_n_9005);
  xnor csa_tree_add_51_79_groupi_g36634(csa_tree_add_51_79_groupi_n_9492 ,csa_tree_add_51_79_groupi_n_8031 ,csa_tree_add_51_79_groupi_n_9004);
  xnor csa_tree_add_51_79_groupi_g36635(csa_tree_add_51_79_groupi_n_9490 ,csa_tree_add_51_79_groupi_n_8386 ,csa_tree_add_51_79_groupi_n_9003);
  xnor csa_tree_add_51_79_groupi_g36636(csa_tree_add_51_79_groupi_n_9489 ,csa_tree_add_51_79_groupi_n_8457 ,csa_tree_add_51_79_groupi_n_9002);
  xnor csa_tree_add_51_79_groupi_g36637(csa_tree_add_51_79_groupi_n_9487 ,csa_tree_add_51_79_groupi_n_8469 ,csa_tree_add_51_79_groupi_n_9008);
  xnor csa_tree_add_51_79_groupi_g36638(csa_tree_add_51_79_groupi_n_9486 ,csa_tree_add_51_79_groupi_n_8503 ,csa_tree_add_51_79_groupi_n_9024);
  xnor csa_tree_add_51_79_groupi_g36639(csa_tree_add_51_79_groupi_n_9484 ,csa_tree_add_51_79_groupi_n_8499 ,csa_tree_add_51_79_groupi_n_9020);
  xnor csa_tree_add_51_79_groupi_g36640(csa_tree_add_51_79_groupi_n_9483 ,csa_tree_add_51_79_groupi_n_8486 ,csa_tree_add_51_79_groupi_n_9019);
  xnor csa_tree_add_51_79_groupi_g36641(csa_tree_add_51_79_groupi_n_9482 ,csa_tree_add_51_79_groupi_n_8016 ,csa_tree_add_51_79_groupi_n_9001);
  xnor csa_tree_add_51_79_groupi_g36642(csa_tree_add_51_79_groupi_n_9481 ,csa_tree_add_51_79_groupi_n_8490 ,csa_tree_add_51_79_groupi_n_8975);
  xnor csa_tree_add_51_79_groupi_g36643(csa_tree_add_51_79_groupi_n_9480 ,csa_tree_add_51_79_groupi_n_8494 ,csa_tree_add_51_79_groupi_n_8999);
  xnor csa_tree_add_51_79_groupi_g36644(csa_tree_add_51_79_groupi_n_9479 ,csa_tree_add_51_79_groupi_n_9196 ,csa_tree_add_51_79_groupi_n_8998);
  xnor csa_tree_add_51_79_groupi_g36645(csa_tree_add_51_79_groupi_n_9478 ,csa_tree_add_51_79_groupi_n_8604 ,csa_tree_add_51_79_groupi_n_8997);
  xnor csa_tree_add_51_79_groupi_g36646(csa_tree_add_51_79_groupi_n_9477 ,csa_tree_add_51_79_groupi_n_8372 ,csa_tree_add_51_79_groupi_n_8996);
  xnor csa_tree_add_51_79_groupi_g36647(csa_tree_add_51_79_groupi_n_9476 ,csa_tree_add_51_79_groupi_n_8407 ,csa_tree_add_51_79_groupi_n_8994);
  xnor csa_tree_add_51_79_groupi_g36648(csa_tree_add_51_79_groupi_n_9475 ,csa_tree_add_51_79_groupi_n_8653 ,csa_tree_add_51_79_groupi_n_8993);
  xnor csa_tree_add_51_79_groupi_g36649(csa_tree_add_51_79_groupi_n_9473 ,csa_tree_add_51_79_groupi_n_8618 ,csa_tree_add_51_79_groupi_n_9018);
  xnor csa_tree_add_51_79_groupi_g36650(csa_tree_add_51_79_groupi_n_9472 ,csa_tree_add_51_79_groupi_n_8489 ,csa_tree_add_51_79_groupi_n_8990);
  xnor csa_tree_add_51_79_groupi_g36651(csa_tree_add_51_79_groupi_n_9471 ,csa_tree_add_51_79_groupi_n_8759 ,csa_tree_add_51_79_groupi_n_8989);
  xnor csa_tree_add_51_79_groupi_g36652(csa_tree_add_51_79_groupi_n_9470 ,csa_tree_add_51_79_groupi_n_8496 ,csa_tree_add_51_79_groupi_n_8988);
  xnor csa_tree_add_51_79_groupi_g36653(csa_tree_add_51_79_groupi_n_9469 ,csa_tree_add_51_79_groupi_n_8465 ,csa_tree_add_51_79_groupi_n_9030);
  xnor csa_tree_add_51_79_groupi_g36654(csa_tree_add_51_79_groupi_n_9466 ,csa_tree_add_51_79_groupi_n_8637 ,csa_tree_add_51_79_groupi_n_9016);
  xnor csa_tree_add_51_79_groupi_g36655(csa_tree_add_51_79_groupi_n_9465 ,csa_tree_add_51_79_groupi_n_8441 ,csa_tree_add_51_79_groupi_n_8971);
  xnor csa_tree_add_51_79_groupi_g36656(csa_tree_add_51_79_groupi_n_9464 ,csa_tree_add_51_79_groupi_n_8639 ,csa_tree_add_51_79_groupi_n_8987);
  xnor csa_tree_add_51_79_groupi_g36657(csa_tree_add_51_79_groupi_n_9463 ,csa_tree_add_51_79_groupi_n_8629 ,csa_tree_add_51_79_groupi_n_8986);
  xnor csa_tree_add_51_79_groupi_g36658(csa_tree_add_51_79_groupi_n_9462 ,csa_tree_add_51_79_groupi_n_8622 ,csa_tree_add_51_79_groupi_n_9015);
  xnor csa_tree_add_51_79_groupi_g36659(csa_tree_add_51_79_groupi_n_9461 ,csa_tree_add_51_79_groupi_n_8336 ,csa_tree_add_51_79_groupi_n_8982);
  xnor csa_tree_add_51_79_groupi_g36660(csa_tree_add_51_79_groupi_n_9460 ,csa_tree_add_51_79_groupi_n_8656 ,csa_tree_add_51_79_groupi_n_8995);
  xnor csa_tree_add_51_79_groupi_g36661(csa_tree_add_51_79_groupi_n_9459 ,csa_tree_add_51_79_groupi_n_8505 ,csa_tree_add_51_79_groupi_n_8981);
  xnor csa_tree_add_51_79_groupi_g36662(csa_tree_add_51_79_groupi_n_9458 ,csa_tree_add_51_79_groupi_n_8375 ,csa_tree_add_51_79_groupi_n_9014);
  xnor csa_tree_add_51_79_groupi_g36663(csa_tree_add_51_79_groupi_n_9457 ,csa_tree_add_51_79_groupi_n_8654 ,csa_tree_add_51_79_groupi_n_8992);
  xnor csa_tree_add_51_79_groupi_g36664(csa_tree_add_51_79_groupi_n_9456 ,csa_tree_add_51_79_groupi_n_8815 ,csa_tree_add_51_79_groupi_n_8979);
  xnor csa_tree_add_51_79_groupi_g36665(csa_tree_add_51_79_groupi_n_9455 ,csa_tree_add_51_79_groupi_n_8453 ,csa_tree_add_51_79_groupi_n_8984);
  xnor csa_tree_add_51_79_groupi_g36666(csa_tree_add_51_79_groupi_n_9454 ,csa_tree_add_51_79_groupi_n_8630 ,csa_tree_add_51_79_groupi_n_8983);
  xnor csa_tree_add_51_79_groupi_g36667(csa_tree_add_51_79_groupi_n_9452 ,csa_tree_add_51_79_groupi_n_9078 ,csa_tree_add_51_79_groupi_n_9013);
  xnor csa_tree_add_51_79_groupi_g36668(csa_tree_add_51_79_groupi_n_9451 ,csa_tree_add_51_79_groupi_n_8442 ,csa_tree_add_51_79_groupi_n_8973);
  xnor csa_tree_add_51_79_groupi_g36669(csa_tree_add_51_79_groupi_n_9450 ,csa_tree_add_51_79_groupi_n_8400 ,csa_tree_add_51_79_groupi_n_8978);
  xnor csa_tree_add_51_79_groupi_g36670(csa_tree_add_51_79_groupi_n_9449 ,csa_tree_add_51_79_groupi_n_8801 ,csa_tree_add_51_79_groupi_n_9023);
  xnor csa_tree_add_51_79_groupi_g36671(csa_tree_add_51_79_groupi_n_9447 ,csa_tree_add_51_79_groupi_n_8431 ,csa_tree_add_51_79_groupi_n_8977);
  xnor csa_tree_add_51_79_groupi_g36672(csa_tree_add_51_79_groupi_n_9445 ,csa_tree_add_51_79_groupi_n_8412 ,csa_tree_add_51_79_groupi_n_30);
  xnor csa_tree_add_51_79_groupi_g36673(csa_tree_add_51_79_groupi_n_9444 ,csa_tree_add_51_79_groupi_n_8821 ,csa_tree_add_51_79_groupi_n_9021);
  xnor csa_tree_add_51_79_groupi_g36674(csa_tree_add_51_79_groupi_n_9442 ,csa_tree_add_51_79_groupi_n_8649 ,csa_tree_add_51_79_groupi_n_9026);
  xnor csa_tree_add_51_79_groupi_g36675(csa_tree_add_51_79_groupi_n_9441 ,csa_tree_add_51_79_groupi_n_8487 ,csa_tree_add_51_79_groupi_n_9017);
  xnor csa_tree_add_51_79_groupi_g36676(csa_tree_add_51_79_groupi_n_9440 ,csa_tree_add_51_79_groupi_n_8646 ,csa_tree_add_51_79_groupi_n_9027);
  xnor csa_tree_add_51_79_groupi_g36677(csa_tree_add_51_79_groupi_n_9439 ,csa_tree_add_51_79_groupi_n_8576 ,csa_tree_add_51_79_groupi_n_9025);
  xnor csa_tree_add_51_79_groupi_g36678(csa_tree_add_51_79_groupi_n_9438 ,csa_tree_add_51_79_groupi_n_8371 ,csa_tree_add_51_79_groupi_n_9028);
  not csa_tree_add_51_79_groupi_g36679(csa_tree_add_51_79_groupi_n_9371 ,csa_tree_add_51_79_groupi_n_9372);
  not csa_tree_add_51_79_groupi_g36680(csa_tree_add_51_79_groupi_n_9364 ,csa_tree_add_51_79_groupi_n_9365);
  not csa_tree_add_51_79_groupi_g36681(csa_tree_add_51_79_groupi_n_9355 ,csa_tree_add_51_79_groupi_n_9356);
  or csa_tree_add_51_79_groupi_g36682(csa_tree_add_51_79_groupi_n_9354 ,csa_tree_add_51_79_groupi_n_8814 ,csa_tree_add_51_79_groupi_n_9117);
  nor csa_tree_add_51_79_groupi_g36683(csa_tree_add_51_79_groupi_n_9353 ,csa_tree_add_51_79_groupi_n_8961 ,csa_tree_add_51_79_groupi_n_9175);
  or csa_tree_add_51_79_groupi_g36684(csa_tree_add_51_79_groupi_n_9352 ,csa_tree_add_51_79_groupi_n_8809 ,csa_tree_add_51_79_groupi_n_9155);
  or csa_tree_add_51_79_groupi_g36685(csa_tree_add_51_79_groupi_n_9351 ,csa_tree_add_51_79_groupi_n_8808 ,csa_tree_add_51_79_groupi_n_9169);
  or csa_tree_add_51_79_groupi_g36686(csa_tree_add_51_79_groupi_n_9350 ,csa_tree_add_51_79_groupi_n_9179 ,csa_tree_add_51_79_groupi_n_9180);
  or csa_tree_add_51_79_groupi_g36687(csa_tree_add_51_79_groupi_n_9349 ,csa_tree_add_51_79_groupi_n_8824 ,csa_tree_add_51_79_groupi_n_9055);
  or csa_tree_add_51_79_groupi_g36688(csa_tree_add_51_79_groupi_n_9348 ,csa_tree_add_51_79_groupi_n_8962 ,csa_tree_add_51_79_groupi_n_9174);
  and csa_tree_add_51_79_groupi_g36689(csa_tree_add_51_79_groupi_n_9347 ,csa_tree_add_51_79_groupi_n_9073 ,csa_tree_add_51_79_groupi_n_8791);
  and csa_tree_add_51_79_groupi_g36690(csa_tree_add_51_79_groupi_n_9346 ,csa_tree_add_51_79_groupi_n_8798 ,csa_tree_add_51_79_groupi_n_9164);
  and csa_tree_add_51_79_groupi_g36691(csa_tree_add_51_79_groupi_n_9345 ,csa_tree_add_51_79_groupi_n_9179 ,csa_tree_add_51_79_groupi_n_9180);
  or csa_tree_add_51_79_groupi_g36692(csa_tree_add_51_79_groupi_n_9344 ,csa_tree_add_51_79_groupi_n_9073 ,csa_tree_add_51_79_groupi_n_8791);
  or csa_tree_add_51_79_groupi_g36693(csa_tree_add_51_79_groupi_n_9343 ,csa_tree_add_51_79_groupi_n_8797 ,csa_tree_add_51_79_groupi_n_9161);
  and csa_tree_add_51_79_groupi_g36694(csa_tree_add_51_79_groupi_n_9342 ,csa_tree_add_51_79_groupi_n_9072 ,csa_tree_add_51_79_groupi_n_9189);
  or csa_tree_add_51_79_groupi_g36695(csa_tree_add_51_79_groupi_n_9341 ,csa_tree_add_51_79_groupi_n_9198 ,csa_tree_add_51_79_groupi_n_9153);
  or csa_tree_add_51_79_groupi_g36696(csa_tree_add_51_79_groupi_n_9340 ,csa_tree_add_51_79_groupi_n_9072 ,csa_tree_add_51_79_groupi_n_9189);
  or csa_tree_add_51_79_groupi_g36697(csa_tree_add_51_79_groupi_n_9339 ,csa_tree_add_51_79_groupi_n_8803 ,csa_tree_add_51_79_groupi_n_9061);
  or csa_tree_add_51_79_groupi_g36698(csa_tree_add_51_79_groupi_n_9338 ,csa_tree_add_51_79_groupi_n_8964 ,csa_tree_add_51_79_groupi_n_9063);
  or csa_tree_add_51_79_groupi_g36699(csa_tree_add_51_79_groupi_n_9337 ,csa_tree_add_51_79_groupi_n_8818 ,csa_tree_add_51_79_groupi_n_9065);
  or csa_tree_add_51_79_groupi_g36700(csa_tree_add_51_79_groupi_n_9336 ,csa_tree_add_51_79_groupi_n_8631 ,csa_tree_add_51_79_groupi_n_9068);
  or csa_tree_add_51_79_groupi_g36701(csa_tree_add_51_79_groupi_n_9335 ,csa_tree_add_51_79_groupi_n_8807 ,csa_tree_add_51_79_groupi_n_9167);
  or csa_tree_add_51_79_groupi_g36702(csa_tree_add_51_79_groupi_n_9334 ,csa_tree_add_51_79_groupi_n_8800 ,csa_tree_add_51_79_groupi_n_9138);
  and csa_tree_add_51_79_groupi_g36703(csa_tree_add_51_79_groupi_n_9333 ,csa_tree_add_51_79_groupi_n_8744 ,csa_tree_add_51_79_groupi_n_9081);
  or csa_tree_add_51_79_groupi_g36704(csa_tree_add_51_79_groupi_n_9332 ,csa_tree_add_51_79_groupi_n_8744 ,csa_tree_add_51_79_groupi_n_9081);
  and csa_tree_add_51_79_groupi_g36705(csa_tree_add_51_79_groupi_n_9331 ,csa_tree_add_51_79_groupi_n_8817 ,csa_tree_add_51_79_groupi_n_9143);
  or csa_tree_add_51_79_groupi_g36706(csa_tree_add_51_79_groupi_n_9330 ,csa_tree_add_51_79_groupi_n_8623 ,csa_tree_add_51_79_groupi_n_9172);
  and csa_tree_add_51_79_groupi_g36707(csa_tree_add_51_79_groupi_n_9329 ,csa_tree_add_51_79_groupi_n_8614 ,csa_tree_add_51_79_groupi_n_9084);
  or csa_tree_add_51_79_groupi_g36708(csa_tree_add_51_79_groupi_n_9328 ,csa_tree_add_51_79_groupi_n_9086 ,csa_tree_add_51_79_groupi_n_9142);
  nor csa_tree_add_51_79_groupi_g36709(csa_tree_add_51_79_groupi_n_9327 ,csa_tree_add_51_79_groupi_n_8813 ,csa_tree_add_51_79_groupi_n_9098);
  nor csa_tree_add_51_79_groupi_g36710(csa_tree_add_51_79_groupi_n_9326 ,csa_tree_add_51_79_groupi_n_8614 ,csa_tree_add_51_79_groupi_n_9084);
  or csa_tree_add_51_79_groupi_g36711(csa_tree_add_51_79_groupi_n_9325 ,csa_tree_add_51_79_groupi_n_8823 ,csa_tree_add_51_79_groupi_n_9135);
  or csa_tree_add_51_79_groupi_g36712(csa_tree_add_51_79_groupi_n_9324 ,csa_tree_add_51_79_groupi_n_9201 ,csa_tree_add_51_79_groupi_n_9101);
  nor csa_tree_add_51_79_groupi_g36713(csa_tree_add_51_79_groupi_n_9323 ,csa_tree_add_51_79_groupi_n_8811 ,csa_tree_add_51_79_groupi_n_9094);
  or csa_tree_add_51_79_groupi_g36714(csa_tree_add_51_79_groupi_n_9322 ,csa_tree_add_51_79_groupi_n_8742 ,csa_tree_add_51_79_groupi_n_9194);
  or csa_tree_add_51_79_groupi_g36715(csa_tree_add_51_79_groupi_n_9321 ,csa_tree_add_51_79_groupi_n_8799 ,csa_tree_add_51_79_groupi_n_9089);
  nor csa_tree_add_51_79_groupi_g36716(csa_tree_add_51_79_groupi_n_9320 ,csa_tree_add_51_79_groupi_n_7818 ,csa_tree_add_51_79_groupi_n_9178);
  and csa_tree_add_51_79_groupi_g36717(csa_tree_add_51_79_groupi_n_9319 ,csa_tree_add_51_79_groupi_n_8812 ,csa_tree_add_51_79_groupi_n_9096);
  or csa_tree_add_51_79_groupi_g36718(csa_tree_add_51_79_groupi_n_9318 ,csa_tree_add_51_79_groupi_n_9204 ,csa_tree_add_51_79_groupi_n_9042);
  and csa_tree_add_51_79_groupi_g36719(csa_tree_add_51_79_groupi_n_9317 ,csa_tree_add_51_79_groupi_n_8742 ,csa_tree_add_51_79_groupi_n_9194);
  or csa_tree_add_51_79_groupi_g36720(csa_tree_add_51_79_groupi_n_9316 ,csa_tree_add_51_79_groupi_n_8802 ,csa_tree_add_51_79_groupi_n_9104);
  or csa_tree_add_51_79_groupi_g36721(csa_tree_add_51_79_groupi_n_9315 ,csa_tree_add_51_79_groupi_n_8804 ,csa_tree_add_51_79_groupi_n_9106);
  or csa_tree_add_51_79_groupi_g36722(csa_tree_add_51_79_groupi_n_9314 ,csa_tree_add_51_79_groupi_n_9176 ,csa_tree_add_51_79_groupi_n_9080);
  and csa_tree_add_51_79_groupi_g36723(csa_tree_add_51_79_groupi_n_9313 ,csa_tree_add_51_79_groupi_n_8816 ,csa_tree_add_51_79_groupi_n_9123);
  and csa_tree_add_51_79_groupi_g36724(csa_tree_add_51_79_groupi_n_9312 ,csa_tree_add_51_79_groupi_n_9176 ,csa_tree_add_51_79_groupi_n_9080);
  or csa_tree_add_51_79_groupi_g36725(csa_tree_add_51_79_groupi_n_9311 ,csa_tree_add_51_79_groupi_n_7819 ,csa_tree_add_51_79_groupi_n_9177);
  or csa_tree_add_51_79_groupi_g36726(csa_tree_add_51_79_groupi_n_9310 ,csa_tree_add_51_79_groupi_n_8642 ,csa_tree_add_51_79_groupi_n_9114);
  or csa_tree_add_51_79_groupi_g36727(csa_tree_add_51_79_groupi_n_9309 ,csa_tree_add_51_79_groupi_n_9196 ,csa_tree_add_51_79_groupi_n_8953);
  and csa_tree_add_51_79_groupi_g36728(csa_tree_add_51_79_groupi_n_9403 ,csa_tree_add_51_79_groupi_n_8904 ,csa_tree_add_51_79_groupi_n_9133);
  and csa_tree_add_51_79_groupi_g36729(csa_tree_add_51_79_groupi_n_9402 ,csa_tree_add_51_79_groupi_n_8843 ,csa_tree_add_51_79_groupi_n_9052);
  and csa_tree_add_51_79_groupi_g36730(csa_tree_add_51_79_groupi_n_9401 ,csa_tree_add_51_79_groupi_n_8941 ,csa_tree_add_51_79_groupi_n_9162);
  and csa_tree_add_51_79_groupi_g36731(csa_tree_add_51_79_groupi_n_9400 ,csa_tree_add_51_79_groupi_n_8874 ,csa_tree_add_51_79_groupi_n_9110);
  and csa_tree_add_51_79_groupi_g36732(csa_tree_add_51_79_groupi_n_9399 ,csa_tree_add_51_79_groupi_n_8708 ,csa_tree_add_51_79_groupi_n_9111);
  and csa_tree_add_51_79_groupi_g36733(csa_tree_add_51_79_groupi_n_9398 ,csa_tree_add_51_79_groupi_n_8938 ,csa_tree_add_51_79_groupi_n_9157);
  and csa_tree_add_51_79_groupi_g36734(csa_tree_add_51_79_groupi_n_9397 ,csa_tree_add_51_79_groupi_n_8832 ,csa_tree_add_51_79_groupi_n_9067);
  and csa_tree_add_51_79_groupi_g36735(csa_tree_add_51_79_groupi_n_9396 ,csa_tree_add_51_79_groupi_n_8870 ,csa_tree_add_51_79_groupi_n_9103);
  and csa_tree_add_51_79_groupi_g36736(csa_tree_add_51_79_groupi_n_9395 ,csa_tree_add_51_79_groupi_n_8697 ,csa_tree_add_51_79_groupi_n_9150);
  or csa_tree_add_51_79_groupi_g36737(csa_tree_add_51_79_groupi_n_9394 ,csa_tree_add_51_79_groupi_n_8957 ,csa_tree_add_51_79_groupi_n_9112);
  and csa_tree_add_51_79_groupi_g36738(csa_tree_add_51_79_groupi_n_9393 ,csa_tree_add_51_79_groupi_n_8889 ,csa_tree_add_51_79_groupi_n_9122);
  and csa_tree_add_51_79_groupi_g36739(csa_tree_add_51_79_groupi_n_9392 ,csa_tree_add_51_79_groupi_n_8834 ,csa_tree_add_51_79_groupi_n_9168);
  or csa_tree_add_51_79_groupi_g36740(csa_tree_add_51_79_groupi_n_9391 ,csa_tree_add_51_79_groupi_n_8921 ,csa_tree_add_51_79_groupi_n_9146);
  and csa_tree_add_51_79_groupi_g36741(csa_tree_add_51_79_groupi_n_9390 ,csa_tree_add_51_79_groupi_n_8897 ,csa_tree_add_51_79_groupi_n_9127);
  and csa_tree_add_51_79_groupi_g36742(csa_tree_add_51_79_groupi_n_9389 ,csa_tree_add_51_79_groupi_n_8924 ,csa_tree_add_51_79_groupi_n_9147);
  and csa_tree_add_51_79_groupi_g36743(csa_tree_add_51_79_groupi_n_9388 ,csa_tree_add_51_79_groupi_n_8250 ,csa_tree_add_51_79_groupi_n_9093);
  and csa_tree_add_51_79_groupi_g36744(csa_tree_add_51_79_groupi_n_9387 ,csa_tree_add_51_79_groupi_n_8696 ,csa_tree_add_51_79_groupi_n_9131);
  and csa_tree_add_51_79_groupi_g36745(csa_tree_add_51_79_groupi_n_9386 ,csa_tree_add_51_79_groupi_n_8899 ,csa_tree_add_51_79_groupi_n_9129);
  and csa_tree_add_51_79_groupi_g36746(csa_tree_add_51_79_groupi_n_9385 ,csa_tree_add_51_79_groupi_n_8881 ,csa_tree_add_51_79_groupi_n_9115);
  and csa_tree_add_51_79_groupi_g36747(csa_tree_add_51_79_groupi_n_9384 ,csa_tree_add_51_79_groupi_n_8846 ,csa_tree_add_51_79_groupi_n_9130);
  and csa_tree_add_51_79_groupi_g36748(csa_tree_add_51_79_groupi_n_9383 ,csa_tree_add_51_79_groupi_n_8849 ,csa_tree_add_51_79_groupi_n_9125);
  and csa_tree_add_51_79_groupi_g36749(csa_tree_add_51_79_groupi_n_9382 ,csa_tree_add_51_79_groupi_n_8928 ,csa_tree_add_51_79_groupi_n_9151);
  and csa_tree_add_51_79_groupi_g36750(csa_tree_add_51_79_groupi_n_9381 ,csa_tree_add_51_79_groupi_n_8852 ,csa_tree_add_51_79_groupi_n_9102);
  and csa_tree_add_51_79_groupi_g36751(csa_tree_add_51_79_groupi_n_9380 ,csa_tree_add_51_79_groupi_n_8903 ,csa_tree_add_51_79_groupi_n_9134);
  and csa_tree_add_51_79_groupi_g36752(csa_tree_add_51_79_groupi_n_9379 ,csa_tree_add_51_79_groupi_n_8911 ,csa_tree_add_51_79_groupi_n_9137);
  and csa_tree_add_51_79_groupi_g36753(csa_tree_add_51_79_groupi_n_9378 ,csa_tree_add_51_79_groupi_n_8830 ,csa_tree_add_51_79_groupi_n_9128);
  and csa_tree_add_51_79_groupi_g36754(csa_tree_add_51_79_groupi_n_9377 ,csa_tree_add_51_79_groupi_n_8845 ,csa_tree_add_51_79_groupi_n_9095);
  and csa_tree_add_51_79_groupi_g36755(csa_tree_add_51_79_groupi_n_9376 ,csa_tree_add_51_79_groupi_n_8842 ,csa_tree_add_51_79_groupi_n_9139);
  and csa_tree_add_51_79_groupi_g36756(csa_tree_add_51_79_groupi_n_9375 ,csa_tree_add_51_79_groupi_n_8840 ,csa_tree_add_51_79_groupi_n_9140);
  and csa_tree_add_51_79_groupi_g36757(csa_tree_add_51_79_groupi_n_9374 ,csa_tree_add_51_79_groupi_n_8926 ,csa_tree_add_51_79_groupi_n_9148);
  and csa_tree_add_51_79_groupi_g36758(csa_tree_add_51_79_groupi_n_9373 ,csa_tree_add_51_79_groupi_n_8894 ,csa_tree_add_51_79_groupi_n_9126);
  and csa_tree_add_51_79_groupi_g36759(csa_tree_add_51_79_groupi_n_9372 ,csa_tree_add_51_79_groupi_n_8862 ,csa_tree_add_51_79_groupi_n_9091);
  and csa_tree_add_51_79_groupi_g36760(csa_tree_add_51_79_groupi_n_9370 ,csa_tree_add_51_79_groupi_n_8872 ,csa_tree_add_51_79_groupi_n_9105);
  and csa_tree_add_51_79_groupi_g36761(csa_tree_add_51_79_groupi_n_9369 ,csa_tree_add_51_79_groupi_n_8851 ,csa_tree_add_51_79_groupi_n_9109);
  or csa_tree_add_51_79_groupi_g36762(csa_tree_add_51_79_groupi_n_9368 ,csa_tree_add_51_79_groupi_n_8930 ,csa_tree_add_51_79_groupi_n_9149);
  and csa_tree_add_51_79_groupi_g36763(csa_tree_add_51_79_groupi_n_9367 ,csa_tree_add_51_79_groupi_n_8933 ,csa_tree_add_51_79_groupi_n_9154);
  and csa_tree_add_51_79_groupi_g36764(csa_tree_add_51_79_groupi_n_9366 ,csa_tree_add_51_79_groupi_n_8936 ,csa_tree_add_51_79_groupi_n_9156);
  or csa_tree_add_51_79_groupi_g36765(csa_tree_add_51_79_groupi_n_9365 ,csa_tree_add_51_79_groupi_n_8888 ,csa_tree_add_51_79_groupi_n_9121);
  and csa_tree_add_51_79_groupi_g36766(csa_tree_add_51_79_groupi_n_9363 ,csa_tree_add_51_79_groupi_n_8828 ,csa_tree_add_51_79_groupi_n_9058);
  and csa_tree_add_51_79_groupi_g36767(csa_tree_add_51_79_groupi_n_9362 ,csa_tree_add_51_79_groupi_n_8826 ,csa_tree_add_51_79_groupi_n_9057);
  and csa_tree_add_51_79_groupi_g36768(csa_tree_add_51_79_groupi_n_9361 ,csa_tree_add_51_79_groupi_n_8836 ,csa_tree_add_51_79_groupi_n_9160);
  and csa_tree_add_51_79_groupi_g36769(csa_tree_add_51_79_groupi_n_9360 ,csa_tree_add_51_79_groupi_n_8693 ,csa_tree_add_51_79_groupi_n_9118);
  and csa_tree_add_51_79_groupi_g36770(csa_tree_add_51_79_groupi_n_9359 ,csa_tree_add_51_79_groupi_n_8946 ,csa_tree_add_51_79_groupi_n_9165);
  and csa_tree_add_51_79_groupi_g36771(csa_tree_add_51_79_groupi_n_9358 ,csa_tree_add_51_79_groupi_n_8880 ,csa_tree_add_51_79_groupi_n_9113);
  or csa_tree_add_51_79_groupi_g36772(csa_tree_add_51_79_groupi_n_9357 ,csa_tree_add_51_79_groupi_n_8940 ,csa_tree_add_51_79_groupi_n_9152);
  and csa_tree_add_51_79_groupi_g36773(csa_tree_add_51_79_groupi_n_9356 ,csa_tree_add_51_79_groupi_n_8883 ,csa_tree_add_51_79_groupi_n_9120);
  not csa_tree_add_51_79_groupi_g36774(csa_tree_add_51_79_groupi_n_9301 ,csa_tree_add_51_79_groupi_n_9300);
  not csa_tree_add_51_79_groupi_g36775(csa_tree_add_51_79_groupi_n_9296 ,csa_tree_add_51_79_groupi_n_9295);
  not csa_tree_add_51_79_groupi_g36776(csa_tree_add_51_79_groupi_n_9293 ,csa_tree_add_51_79_groupi_n_9292);
  not csa_tree_add_51_79_groupi_g36777(csa_tree_add_51_79_groupi_n_9281 ,csa_tree_add_51_79_groupi_n_9280);
  not csa_tree_add_51_79_groupi_g36778(csa_tree_add_51_79_groupi_n_9277 ,csa_tree_add_51_79_groupi_n_9278);
  not csa_tree_add_51_79_groupi_g36779(csa_tree_add_51_79_groupi_n_9275 ,csa_tree_add_51_79_groupi_n_9274);
  not csa_tree_add_51_79_groupi_g36780(csa_tree_add_51_79_groupi_n_9273 ,csa_tree_add_51_79_groupi_n_9272);
  not csa_tree_add_51_79_groupi_g36781(csa_tree_add_51_79_groupi_n_9270 ,csa_tree_add_51_79_groupi_n_9269);
  not csa_tree_add_51_79_groupi_g36782(csa_tree_add_51_79_groupi_n_9260 ,csa_tree_add_51_79_groupi_n_9261);
  not csa_tree_add_51_79_groupi_g36783(csa_tree_add_51_79_groupi_n_9253 ,csa_tree_add_51_79_groupi_n_9254);
  and csa_tree_add_51_79_groupi_g36784(csa_tree_add_51_79_groupi_n_9248 ,csa_tree_add_51_79_groupi_n_9070 ,csa_tree_add_51_79_groupi_n_8750);
  and csa_tree_add_51_79_groupi_g36785(csa_tree_add_51_79_groupi_n_9247 ,csa_tree_add_51_79_groupi_n_8418 ,csa_tree_add_51_79_groupi_n_9078);
  nor csa_tree_add_51_79_groupi_g36786(csa_tree_add_51_79_groupi_n_9246 ,csa_tree_add_51_79_groupi_n_8418 ,csa_tree_add_51_79_groupi_n_9078);
  nor csa_tree_add_51_79_groupi_g36787(csa_tree_add_51_79_groupi_n_9245 ,csa_tree_add_51_79_groupi_n_8770 ,csa_tree_add_51_79_groupi_n_9071);
  and csa_tree_add_51_79_groupi_g36788(csa_tree_add_51_79_groupi_n_9244 ,csa_tree_add_51_79_groupi_n_8770 ,csa_tree_add_51_79_groupi_n_9071);
  or csa_tree_add_51_79_groupi_g36789(csa_tree_add_51_79_groupi_n_9243 ,csa_tree_add_51_79_groupi_n_9070 ,csa_tree_add_51_79_groupi_n_8750);
  or csa_tree_add_51_79_groupi_g36790(csa_tree_add_51_79_groupi_n_9242 ,csa_tree_add_51_79_groupi_n_8819 ,csa_tree_add_51_79_groupi_n_9047);
  nor csa_tree_add_51_79_groupi_g36791(csa_tree_add_51_79_groupi_n_9241 ,csa_tree_add_51_79_groupi_n_9077 ,csa_tree_add_51_79_groupi_n_8787);
  or csa_tree_add_51_79_groupi_g36792(csa_tree_add_51_79_groupi_n_9240 ,csa_tree_add_51_79_groupi_n_9076 ,csa_tree_add_51_79_groupi_n_8788);
  nor csa_tree_add_51_79_groupi_g36793(csa_tree_add_51_79_groupi_n_9239 ,csa_tree_add_51_79_groupi_n_9187 ,csa_tree_add_51_79_groupi_n_9074);
  or csa_tree_add_51_79_groupi_g36794(csa_tree_add_51_79_groupi_n_9238 ,csa_tree_add_51_79_groupi_n_9186 ,csa_tree_add_51_79_groupi_n_9075);
  or csa_tree_add_51_79_groupi_g36795(csa_tree_add_51_79_groupi_n_9237 ,csa_tree_add_51_79_groupi_n_8822 ,csa_tree_add_51_79_groupi_n_9053);
  xnor csa_tree_add_51_79_groupi_g36796(csa_tree_add_51_79_groupi_n_9236 ,csa_tree_add_51_79_groupi_n_8606 ,csa_tree_add_51_79_groupi_n_8790);
  xnor csa_tree_add_51_79_groupi_g36797(csa_tree_add_51_79_groupi_n_9235 ,csa_tree_add_51_79_groupi_n_8760 ,csa_tree_add_51_79_groupi_n_8799);
  xnor csa_tree_add_51_79_groupi_g36798(csa_tree_add_51_79_groupi_n_9234 ,csa_tree_add_51_79_groupi_n_8824 ,csa_tree_add_51_79_groupi_n_8786);
  xnor csa_tree_add_51_79_groupi_g36799(csa_tree_add_51_79_groupi_n_9233 ,csa_tree_add_51_79_groupi_n_8172 ,csa_tree_add_51_79_groupi_n_8719);
  xnor csa_tree_add_51_79_groupi_g36800(csa_tree_add_51_79_groupi_n_9232 ,csa_tree_add_51_79_groupi_n_8794 ,csa_tree_add_51_79_groupi_n_8778);
  xnor csa_tree_add_51_79_groupi_g36801(csa_tree_add_51_79_groupi_n_9231 ,csa_tree_add_51_79_groupi_n_8603 ,csa_tree_add_51_79_groupi_n_8746);
  xnor csa_tree_add_51_79_groupi_g36802(csa_tree_add_51_79_groupi_n_9230 ,csa_tree_add_51_79_groupi_n_8812 ,csa_tree_add_51_79_groupi_n_8732);
  xnor csa_tree_add_51_79_groupi_g36803(csa_tree_add_51_79_groupi_n_9229 ,csa_tree_add_51_79_groupi_n_8800 ,csa_tree_add_51_79_groupi_n_8480);
  xnor csa_tree_add_51_79_groupi_g36804(csa_tree_add_51_79_groupi_n_9228 ,csa_tree_add_51_79_groupi_n_8752 ,csa_tree_add_51_79_groupi_n_8774);
  xnor csa_tree_add_51_79_groupi_g36805(csa_tree_add_51_79_groupi_n_9227 ,csa_tree_add_51_79_groupi_n_8763 ,csa_tree_add_51_79_groupi_n_8754);
  xnor csa_tree_add_51_79_groupi_g36806(csa_tree_add_51_79_groupi_n_9226 ,csa_tree_add_51_79_groupi_n_8749 ,csa_tree_add_51_79_groupi_n_8725);
  xnor csa_tree_add_51_79_groupi_g36807(csa_tree_add_51_79_groupi_n_9225 ,csa_tree_add_51_79_groupi_n_8740 ,csa_tree_add_51_79_groupi_n_8816);
  xor csa_tree_add_51_79_groupi_g36808(csa_tree_add_51_79_groupi_n_9224 ,csa_tree_add_51_79_groupi_n_8737 ,csa_tree_add_51_79_groupi_n_8814);
  xnor csa_tree_add_51_79_groupi_g36809(csa_tree_add_51_79_groupi_n_9223 ,csa_tree_add_51_79_groupi_n_8782 ,csa_tree_add_51_79_groupi_n_8809);
  xnor csa_tree_add_51_79_groupi_g36810(csa_tree_add_51_79_groupi_n_9222 ,csa_tree_add_51_79_groupi_n_8589 ,csa_tree_add_51_79_groupi_n_8717);
  xnor csa_tree_add_51_79_groupi_g36811(csa_tree_add_51_79_groupi_n_9221 ,csa_tree_add_51_79_groupi_n_8735 ,csa_tree_add_51_79_groupi_n_8720);
  xnor csa_tree_add_51_79_groupi_g36812(csa_tree_add_51_79_groupi_n_9220 ,csa_tree_add_51_79_groupi_n_8813 ,csa_tree_add_51_79_groupi_n_8958);
  xnor csa_tree_add_51_79_groupi_g36813(csa_tree_add_51_79_groupi_n_9219 ,csa_tree_add_51_79_groupi_n_8811 ,csa_tree_add_51_79_groupi_n_8452);
  xnor csa_tree_add_51_79_groupi_g36814(csa_tree_add_51_79_groupi_n_9218 ,csa_tree_add_51_79_groupi_n_8818 ,csa_tree_add_51_79_groupi_n_8741);
  xnor csa_tree_add_51_79_groupi_g36815(csa_tree_add_51_79_groupi_n_9217 ,csa_tree_add_51_79_groupi_n_8721 ,csa_tree_add_51_79_groupi_n_8722);
  xnor csa_tree_add_51_79_groupi_g36816(csa_tree_add_51_79_groupi_n_9216 ,csa_tree_add_51_79_groupi_n_8574 ,csa_tree_add_51_79_groupi_n_8768);
  xnor csa_tree_add_51_79_groupi_g36817(csa_tree_add_51_79_groupi_n_9215 ,csa_tree_add_51_79_groupi_n_8592 ,csa_tree_add_51_79_groupi_n_8965);
  xnor csa_tree_add_51_79_groupi_g36818(csa_tree_add_51_79_groupi_n_9214 ,csa_tree_add_51_79_groupi_n_8969 ,csa_tree_add_51_79_groupi_n_8152);
  xnor csa_tree_add_51_79_groupi_g36819(csa_tree_add_51_79_groupi_n_9213 ,csa_tree_add_51_79_groupi_n_8771 ,csa_tree_add_51_79_groupi_n_8819);
  xnor csa_tree_add_51_79_groupi_g36820(csa_tree_add_51_79_groupi_n_9212 ,csa_tree_add_51_79_groupi_n_8807 ,csa_tree_add_51_79_groupi_n_8766);
  xnor csa_tree_add_51_79_groupi_g36821(csa_tree_add_51_79_groupi_n_9211 ,csa_tree_add_51_79_groupi_n_8769 ,csa_tree_add_51_79_groupi_n_8808);
  xnor csa_tree_add_51_79_groupi_g36822(csa_tree_add_51_79_groupi_n_9210 ,csa_tree_add_51_79_groupi_n_8959 ,csa_tree_add_51_79_groupi_n_8631);
  xnor csa_tree_add_51_79_groupi_g36823(csa_tree_add_51_79_groupi_n_9209 ,csa_tree_add_51_79_groupi_n_8734 ,csa_tree_add_51_79_groupi_n_8736);
  xnor csa_tree_add_51_79_groupi_g36824(csa_tree_add_51_79_groupi_n_9208 ,csa_tree_add_51_79_groupi_n_8729 ,csa_tree_add_51_79_groupi_n_8730);
  xnor csa_tree_add_51_79_groupi_g36825(csa_tree_add_51_79_groupi_n_9207 ,csa_tree_add_51_79_groupi_n_8779 ,csa_tree_add_51_79_groupi_n_8822);
  and csa_tree_add_51_79_groupi_g36826(csa_tree_add_51_79_groupi_n_9308 ,csa_tree_add_51_79_groupi_n_8702 ,csa_tree_add_51_79_groupi_n_9032);
  and csa_tree_add_51_79_groupi_g36827(csa_tree_add_51_79_groupi_n_9307 ,csa_tree_add_51_79_groupi_n_8895 ,csa_tree_add_51_79_groupi_n_9049);
  and csa_tree_add_51_79_groupi_g36828(csa_tree_add_51_79_groupi_n_9306 ,csa_tree_add_51_79_groupi_n_8856 ,csa_tree_add_51_79_groupi_n_9041);
  and csa_tree_add_51_79_groupi_g36829(csa_tree_add_51_79_groupi_n_9305 ,csa_tree_add_51_79_groupi_n_8945 ,csa_tree_add_51_79_groupi_n_9031);
  xnor csa_tree_add_51_79_groupi_g36830(csa_tree_add_51_79_groupi_n_9304 ,csa_tree_add_51_79_groupi_n_8820 ,csa_tree_add_51_79_groupi_n_8344);
  xnor csa_tree_add_51_79_groupi_g36831(csa_tree_add_51_79_groupi_n_9303 ,csa_tree_add_51_79_groupi_n_8182 ,csa_tree_add_51_79_groupi_n_8675);
  and csa_tree_add_51_79_groupi_g36832(csa_tree_add_51_79_groupi_n_9302 ,csa_tree_add_51_79_groupi_n_8705 ,csa_tree_add_51_79_groupi_n_9033);
  or csa_tree_add_51_79_groupi_g36833(csa_tree_add_51_79_groupi_n_9300 ,csa_tree_add_51_79_groupi_n_8699 ,csa_tree_add_51_79_groupi_n_9034);
  and csa_tree_add_51_79_groupi_g36834(csa_tree_add_51_79_groupi_n_9299 ,csa_tree_add_51_79_groupi_n_8710 ,csa_tree_add_51_79_groupi_n_9036);
  and csa_tree_add_51_79_groupi_g36835(csa_tree_add_51_79_groupi_n_9298 ,csa_tree_add_51_79_groupi_n_8714 ,csa_tree_add_51_79_groupi_n_9039);
  and csa_tree_add_51_79_groupi_g36836(csa_tree_add_51_79_groupi_n_9297 ,csa_tree_add_51_79_groupi_n_8951 ,csa_tree_add_51_79_groupi_n_9044);
  xnor csa_tree_add_51_79_groupi_g36837(csa_tree_add_51_79_groupi_n_9295 ,csa_tree_add_51_79_groupi_n_8409 ,csa_tree_add_51_79_groupi_n_8684);
  xnor csa_tree_add_51_79_groupi_g36838(csa_tree_add_51_79_groupi_n_9294 ,csa_tree_add_51_79_groupi_n_7825 ,csa_tree_add_51_79_groupi_n_8661);
  xnor csa_tree_add_51_79_groupi_g36839(csa_tree_add_51_79_groupi_n_9292 ,csa_tree_add_51_79_groupi_n_8339 ,csa_tree_add_51_79_groupi_n_8683);
  and csa_tree_add_51_79_groupi_g36840(csa_tree_add_51_79_groupi_n_9291 ,csa_tree_add_51_79_groupi_n_8861 ,csa_tree_add_51_79_groupi_n_9051);
  xnor csa_tree_add_51_79_groupi_g36841(csa_tree_add_51_79_groupi_n_9290 ,csa_tree_add_51_79_groupi_n_8173 ,csa_tree_add_51_79_groupi_n_8682);
  xnor csa_tree_add_51_79_groupi_g36842(csa_tree_add_51_79_groupi_n_9289 ,csa_tree_add_51_79_groupi_n_8293 ,csa_tree_add_51_79_groupi_n_8681);
  or csa_tree_add_51_79_groupi_g36843(csa_tree_add_51_79_groupi_n_9288 ,csa_tree_add_51_79_groupi_n_8923 ,csa_tree_add_51_79_groupi_n_9035);
  xnor csa_tree_add_51_79_groupi_g36844(csa_tree_add_51_79_groupi_n_9287 ,csa_tree_add_51_79_groupi_n_7803 ,csa_tree_add_51_79_groupi_n_8677);
  and csa_tree_add_51_79_groupi_g36845(csa_tree_add_51_79_groupi_n_9286 ,csa_tree_add_51_79_groupi_n_8866 ,csa_tree_add_51_79_groupi_n_9050);
  and csa_tree_add_51_79_groupi_g36846(csa_tree_add_51_79_groupi_n_9285 ,csa_tree_add_51_79_groupi_n_8906 ,csa_tree_add_51_79_groupi_n_9040);
  and csa_tree_add_51_79_groupi_g36847(csa_tree_add_51_79_groupi_n_9284 ,csa_tree_add_51_79_groupi_n_8712 ,csa_tree_add_51_79_groupi_n_9038);
  and csa_tree_add_51_79_groupi_g36848(csa_tree_add_51_79_groupi_n_9283 ,csa_tree_add_51_79_groupi_n_8691 ,csa_tree_add_51_79_groupi_n_9037);
  xnor csa_tree_add_51_79_groupi_g36849(csa_tree_add_51_79_groupi_n_9282 ,csa_tree_add_51_79_groupi_n_8331 ,csa_tree_add_51_79_groupi_n_8676);
  xnor csa_tree_add_51_79_groupi_g36850(csa_tree_add_51_79_groupi_n_9280 ,csa_tree_add_51_79_groupi_n_8485 ,csa_tree_add_51_79_groupi_n_8689);
  xnor csa_tree_add_51_79_groupi_g36851(csa_tree_add_51_79_groupi_n_9279 ,csa_tree_add_51_79_groupi_n_8343 ,csa_tree_add_51_79_groupi_n_8688);
  xnor csa_tree_add_51_79_groupi_g36852(csa_tree_add_51_79_groupi_n_9278 ,csa_tree_add_51_79_groupi_n_8337 ,csa_tree_add_51_79_groupi_n_8679);
  xnor csa_tree_add_51_79_groupi_g36853(csa_tree_add_51_79_groupi_n_9276 ,csa_tree_add_51_79_groupi_n_8154 ,csa_tree_add_51_79_groupi_n_8690);
  xnor csa_tree_add_51_79_groupi_g36854(csa_tree_add_51_79_groupi_n_9274 ,csa_tree_add_51_79_groupi_n_8388 ,csa_tree_add_51_79_groupi_n_8665);
  xnor csa_tree_add_51_79_groupi_g36855(csa_tree_add_51_79_groupi_n_9272 ,csa_tree_add_51_79_groupi_n_8473 ,csa_tree_add_51_79_groupi_n_8662);
  xnor csa_tree_add_51_79_groupi_g36856(csa_tree_add_51_79_groupi_n_9271 ,csa_tree_add_51_79_groupi_n_8275 ,csa_tree_add_51_79_groupi_n_8674);
  and csa_tree_add_51_79_groupi_g36857(csa_tree_add_51_79_groupi_n_9269 ,csa_tree_add_51_79_groupi_n_8878 ,csa_tree_add_51_79_groupi_n_9046);
  xnor csa_tree_add_51_79_groupi_g36858(csa_tree_add_51_79_groupi_n_9268 ,csa_tree_add_51_79_groupi_n_8315 ,csa_tree_add_51_79_groupi_n_8687);
  xnor csa_tree_add_51_79_groupi_g36859(csa_tree_add_51_79_groupi_n_9267 ,csa_tree_add_51_79_groupi_n_8310 ,csa_tree_add_51_79_groupi_n_8666);
  xnor csa_tree_add_51_79_groupi_g36860(csa_tree_add_51_79_groupi_n_9266 ,csa_tree_add_51_79_groupi_n_8318 ,csa_tree_add_51_79_groupi_n_8673);
  xnor csa_tree_add_51_79_groupi_g36861(csa_tree_add_51_79_groupi_n_9265 ,csa_tree_add_51_79_groupi_n_8181 ,csa_tree_add_51_79_groupi_n_8663);
  xnor csa_tree_add_51_79_groupi_g36862(csa_tree_add_51_79_groupi_n_9264 ,csa_tree_add_51_79_groupi_n_8314 ,csa_tree_add_51_79_groupi_n_8672);
  xnor csa_tree_add_51_79_groupi_g36863(csa_tree_add_51_79_groupi_n_9263 ,csa_tree_add_51_79_groupi_n_8023 ,csa_tree_add_51_79_groupi_n_8671);
  xnor csa_tree_add_51_79_groupi_g36864(csa_tree_add_51_79_groupi_n_9262 ,csa_tree_add_51_79_groupi_n_8330 ,csa_tree_add_51_79_groupi_n_8680);
  xnor csa_tree_add_51_79_groupi_g36865(csa_tree_add_51_79_groupi_n_9261 ,csa_tree_add_51_79_groupi_n_8288 ,csa_tree_add_51_79_groupi_n_8670);
  xnor csa_tree_add_51_79_groupi_g36866(csa_tree_add_51_79_groupi_n_9259 ,csa_tree_add_51_79_groupi_n_8658 ,csa_tree_add_51_79_groupi_n_8669);
  xnor csa_tree_add_51_79_groupi_g36867(csa_tree_add_51_79_groupi_n_9258 ,csa_tree_add_51_79_groupi_n_8338 ,csa_tree_add_51_79_groupi_n_8686);
  xnor csa_tree_add_51_79_groupi_g36868(csa_tree_add_51_79_groupi_n_9257 ,csa_tree_add_51_79_groupi_n_8300 ,csa_tree_add_51_79_groupi_n_8668);
  xnor csa_tree_add_51_79_groupi_g36869(csa_tree_add_51_79_groupi_n_9256 ,csa_tree_add_51_79_groupi_n_8320 ,csa_tree_add_51_79_groupi_n_8667);
  xnor csa_tree_add_51_79_groupi_g36870(csa_tree_add_51_79_groupi_n_9255 ,csa_tree_add_51_79_groupi_n_8174 ,csa_tree_add_51_79_groupi_n_8678);
  xnor csa_tree_add_51_79_groupi_g36871(csa_tree_add_51_79_groupi_n_9254 ,csa_tree_add_51_79_groupi_n_8280 ,csa_tree_add_51_79_groupi_n_8664);
  xnor csa_tree_add_51_79_groupi_g36872(csa_tree_add_51_79_groupi_n_9252 ,csa_tree_add_51_79_groupi_n_8175 ,csa_tree_add_51_79_groupi_n_8685);
  and csa_tree_add_51_79_groupi_g36873(csa_tree_add_51_79_groupi_n_9251 ,csa_tree_add_51_79_groupi_n_8908 ,csa_tree_add_51_79_groupi_n_9045);
  xnor csa_tree_add_51_79_groupi_g36874(csa_tree_add_51_79_groupi_n_9250 ,csa_tree_add_51_79_groupi_n_8309 ,csa_tree_add_51_79_groupi_n_8660);
  xnor csa_tree_add_51_79_groupi_g36875(csa_tree_add_51_79_groupi_n_9249 ,csa_tree_add_51_79_groupi_n_8342 ,csa_tree_add_51_79_groupi_n_8659);
  not csa_tree_add_51_79_groupi_g36877(csa_tree_add_51_79_groupi_n_9192 ,csa_tree_add_51_79_groupi_n_9193);
  not csa_tree_add_51_79_groupi_g36878(csa_tree_add_51_79_groupi_n_9187 ,csa_tree_add_51_79_groupi_n_9186);
  not csa_tree_add_51_79_groupi_g36879(csa_tree_add_51_79_groupi_n_9184 ,csa_tree_add_51_79_groupi_n_9185);
  not csa_tree_add_51_79_groupi_g36880(csa_tree_add_51_79_groupi_n_9183 ,csa_tree_add_51_79_groupi_n_9182);
  not csa_tree_add_51_79_groupi_g36881(csa_tree_add_51_79_groupi_n_9177 ,csa_tree_add_51_79_groupi_n_9178);
  not csa_tree_add_51_79_groupi_g36882(csa_tree_add_51_79_groupi_n_9174 ,csa_tree_add_51_79_groupi_n_9175);
  or csa_tree_add_51_79_groupi_g36883(csa_tree_add_51_79_groupi_n_9173 ,csa_tree_add_51_79_groupi_n_8959 ,csa_tree_add_51_79_groupi_n_8423);
  and csa_tree_add_51_79_groupi_g36884(csa_tree_add_51_79_groupi_n_9172 ,csa_tree_add_51_79_groupi_n_8594 ,csa_tree_add_51_79_groupi_n_8759);
  or csa_tree_add_51_79_groupi_g36885(csa_tree_add_51_79_groupi_n_9171 ,csa_tree_add_51_79_groupi_n_8594 ,csa_tree_add_51_79_groupi_n_8759);
  or csa_tree_add_51_79_groupi_g36886(csa_tree_add_51_79_groupi_n_9170 ,csa_tree_add_51_79_groupi_n_8756 ,csa_tree_add_51_79_groupi_n_8769);
  and csa_tree_add_51_79_groupi_g36887(csa_tree_add_51_79_groupi_n_9169 ,csa_tree_add_51_79_groupi_n_8756 ,csa_tree_add_51_79_groupi_n_8769);
  or csa_tree_add_51_79_groupi_g36888(csa_tree_add_51_79_groupi_n_9168 ,csa_tree_add_51_79_groupi_n_8652 ,csa_tree_add_51_79_groupi_n_8833);
  and csa_tree_add_51_79_groupi_g36889(csa_tree_add_51_79_groupi_n_9167 ,csa_tree_add_51_79_groupi_n_8766 ,csa_tree_add_51_79_groupi_n_8764);
  nor csa_tree_add_51_79_groupi_g36890(csa_tree_add_51_79_groupi_n_9166 ,csa_tree_add_51_79_groupi_n_8573 ,csa_tree_add_51_79_groupi_n_8768);
  or csa_tree_add_51_79_groupi_g36891(csa_tree_add_51_79_groupi_n_9165 ,csa_tree_add_51_79_groupi_n_8321 ,csa_tree_add_51_79_groupi_n_8934);
  or csa_tree_add_51_79_groupi_g36892(csa_tree_add_51_79_groupi_n_9164 ,csa_tree_add_51_79_groupi_n_8574 ,csa_tree_add_51_79_groupi_n_8767);
  or csa_tree_add_51_79_groupi_g36893(csa_tree_add_51_79_groupi_n_9163 ,csa_tree_add_51_79_groupi_n_8762 ,csa_tree_add_51_79_groupi_n_8754);
  or csa_tree_add_51_79_groupi_g36894(csa_tree_add_51_79_groupi_n_9162 ,csa_tree_add_51_79_groupi_n_8654 ,csa_tree_add_51_79_groupi_n_8939);
  nor csa_tree_add_51_79_groupi_g36895(csa_tree_add_51_79_groupi_n_9161 ,csa_tree_add_51_79_groupi_n_8763 ,csa_tree_add_51_79_groupi_n_8753);
  or csa_tree_add_51_79_groupi_g36896(csa_tree_add_51_79_groupi_n_9160 ,csa_tree_add_51_79_groupi_n_8653 ,csa_tree_add_51_79_groupi_n_8835);
  or csa_tree_add_51_79_groupi_g36897(csa_tree_add_51_79_groupi_n_9159 ,csa_tree_add_51_79_groupi_n_8752 ,csa_tree_add_51_79_groupi_n_8773);
  or csa_tree_add_51_79_groupi_g36898(csa_tree_add_51_79_groupi_n_9158 ,csa_tree_add_51_79_groupi_n_8766 ,csa_tree_add_51_79_groupi_n_8764);
  or csa_tree_add_51_79_groupi_g36899(csa_tree_add_51_79_groupi_n_9157 ,csa_tree_add_51_79_groupi_n_8506 ,csa_tree_add_51_79_groupi_n_8937);
  or csa_tree_add_51_79_groupi_g36900(csa_tree_add_51_79_groupi_n_9156 ,csa_tree_add_51_79_groupi_n_8324 ,csa_tree_add_51_79_groupi_n_8935);
  nor csa_tree_add_51_79_groupi_g36901(csa_tree_add_51_79_groupi_n_9155 ,csa_tree_add_51_79_groupi_n_8784 ,csa_tree_add_51_79_groupi_n_8782);
  or csa_tree_add_51_79_groupi_g36902(csa_tree_add_51_79_groupi_n_9154 ,csa_tree_add_51_79_groupi_n_8640 ,csa_tree_add_51_79_groupi_n_8929);
  nor csa_tree_add_51_79_groupi_g36903(csa_tree_add_51_79_groupi_n_9153 ,csa_tree_add_51_79_groupi_n_8751 ,csa_tree_add_51_79_groupi_n_8774);
  and csa_tree_add_51_79_groupi_g36904(csa_tree_add_51_79_groupi_n_9152 ,csa_tree_add_51_79_groupi_n_8323 ,csa_tree_add_51_79_groupi_n_8918);
  or csa_tree_add_51_79_groupi_g36905(csa_tree_add_51_79_groupi_n_9151 ,csa_tree_add_51_79_groupi_n_8634 ,csa_tree_add_51_79_groupi_n_8927);
  or csa_tree_add_51_79_groupi_g36906(csa_tree_add_51_79_groupi_n_9150 ,csa_tree_add_51_79_groupi_n_8628 ,csa_tree_add_51_79_groupi_n_8695);
  and csa_tree_add_51_79_groupi_g36907(csa_tree_add_51_79_groupi_n_9149 ,csa_tree_add_51_79_groupi_n_8633 ,csa_tree_add_51_79_groupi_n_8922);
  or csa_tree_add_51_79_groupi_g36908(csa_tree_add_51_79_groupi_n_9148 ,csa_tree_add_51_79_groupi_n_8489 ,csa_tree_add_51_79_groupi_n_8925);
  or csa_tree_add_51_79_groupi_g36909(csa_tree_add_51_79_groupi_n_9147 ,csa_tree_add_51_79_groupi_n_8496 ,csa_tree_add_51_79_groupi_n_8919);
  nor csa_tree_add_51_79_groupi_g36910(csa_tree_add_51_79_groupi_n_9146 ,csa_tree_add_51_79_groupi_n_8625 ,csa_tree_add_51_79_groupi_n_8917);
  nor csa_tree_add_51_79_groupi_g36911(csa_tree_add_51_79_groupi_n_9145 ,csa_tree_add_51_79_groupi_n_8749 ,csa_tree_add_51_79_groupi_n_8724);
  or csa_tree_add_51_79_groupi_g36912(csa_tree_add_51_79_groupi_n_9144 ,csa_tree_add_51_79_groupi_n_8755 ,csa_tree_add_51_79_groupi_n_8747);
  or csa_tree_add_51_79_groupi_g36913(csa_tree_add_51_79_groupi_n_9143 ,csa_tree_add_51_79_groupi_n_8748 ,csa_tree_add_51_79_groupi_n_8725);
  and csa_tree_add_51_79_groupi_g36914(csa_tree_add_51_79_groupi_n_9142 ,csa_tree_add_51_79_groupi_n_8755 ,csa_tree_add_51_79_groupi_n_8747);
  or csa_tree_add_51_79_groupi_g36915(csa_tree_add_51_79_groupi_n_9141 ,csa_tree_add_51_79_groupi_n_8783 ,csa_tree_add_51_79_groupi_n_8781);
  or csa_tree_add_51_79_groupi_g36916(csa_tree_add_51_79_groupi_n_9140 ,csa_tree_add_51_79_groupi_n_8495 ,csa_tree_add_51_79_groupi_n_8839);
  or csa_tree_add_51_79_groupi_g36917(csa_tree_add_51_79_groupi_n_9139 ,csa_tree_add_51_79_groupi_n_8630 ,csa_tree_add_51_79_groupi_n_8841);
  and csa_tree_add_51_79_groupi_g36918(csa_tree_add_51_79_groupi_n_9138 ,csa_tree_add_51_79_groupi_n_8480 ,csa_tree_add_51_79_groupi_n_8723);
  or csa_tree_add_51_79_groupi_g36919(csa_tree_add_51_79_groupi_n_9137 ,csa_tree_add_51_79_groupi_n_8629 ,csa_tree_add_51_79_groupi_n_8910);
  or csa_tree_add_51_79_groupi_g36920(csa_tree_add_51_79_groupi_n_9136 ,csa_tree_add_51_79_groupi_n_8171 ,csa_tree_add_51_79_groupi_n_8718);
  nor csa_tree_add_51_79_groupi_g36921(csa_tree_add_51_79_groupi_n_9135 ,csa_tree_add_51_79_groupi_n_8172 ,csa_tree_add_51_79_groupi_n_8719);
  or csa_tree_add_51_79_groupi_g36922(csa_tree_add_51_79_groupi_n_9134 ,csa_tree_add_51_79_groupi_n_8334 ,csa_tree_add_51_79_groupi_n_8902);
  or csa_tree_add_51_79_groupi_g36923(csa_tree_add_51_79_groupi_n_9133 ,csa_tree_add_51_79_groupi_n_8655 ,csa_tree_add_51_79_groupi_n_8901);
  or csa_tree_add_51_79_groupi_g36924(csa_tree_add_51_79_groupi_n_9132 ,csa_tree_add_51_79_groupi_n_8480 ,csa_tree_add_51_79_groupi_n_8723);
  or csa_tree_add_51_79_groupi_g36925(csa_tree_add_51_79_groupi_n_9131 ,csa_tree_add_51_79_groupi_n_8651 ,csa_tree_add_51_79_groupi_n_8694);
  or csa_tree_add_51_79_groupi_g36926(csa_tree_add_51_79_groupi_n_9130 ,csa_tree_add_51_79_groupi_n_8650 ,csa_tree_add_51_79_groupi_n_8885);
  or csa_tree_add_51_79_groupi_g36927(csa_tree_add_51_79_groupi_n_9129 ,csa_tree_add_51_79_groupi_n_8336 ,csa_tree_add_51_79_groupi_n_8898);
  or csa_tree_add_51_79_groupi_g36928(csa_tree_add_51_79_groupi_n_9128 ,csa_tree_add_51_79_groupi_n_8656 ,csa_tree_add_51_79_groupi_n_8829);
  or csa_tree_add_51_79_groupi_g36929(csa_tree_add_51_79_groupi_n_9127 ,csa_tree_add_51_79_groupi_n_8505 ,csa_tree_add_51_79_groupi_n_8896);
  or csa_tree_add_51_79_groupi_g36930(csa_tree_add_51_79_groupi_n_9126 ,csa_tree_add_51_79_groupi_n_8341 ,csa_tree_add_51_79_groupi_n_8893);
  or csa_tree_add_51_79_groupi_g36931(csa_tree_add_51_79_groupi_n_9125 ,csa_tree_add_51_79_groupi_n_8648 ,csa_tree_add_51_79_groupi_n_8847);
  nor csa_tree_add_51_79_groupi_g36932(csa_tree_add_51_79_groupi_n_9124 ,csa_tree_add_51_79_groupi_n_8740 ,csa_tree_add_51_79_groupi_n_8758);
  or csa_tree_add_51_79_groupi_g36933(csa_tree_add_51_79_groupi_n_9123 ,csa_tree_add_51_79_groupi_n_8739 ,csa_tree_add_51_79_groupi_n_8757);
  or csa_tree_add_51_79_groupi_g36934(csa_tree_add_51_79_groupi_n_9122 ,csa_tree_add_51_79_groupi_n_8647 ,csa_tree_add_51_79_groupi_n_8887);
  and csa_tree_add_51_79_groupi_g36935(csa_tree_add_51_79_groupi_n_9121 ,csa_tree_add_51_79_groupi_n_8649 ,csa_tree_add_51_79_groupi_n_8884);
  or csa_tree_add_51_79_groupi_g36936(csa_tree_add_51_79_groupi_n_9120 ,csa_tree_add_51_79_groupi_n_8487 ,csa_tree_add_51_79_groupi_n_8882);
  or csa_tree_add_51_79_groupi_g36937(csa_tree_add_51_79_groupi_n_9119 ,csa_tree_add_51_79_groupi_n_8738 ,csa_tree_add_51_79_groupi_n_8737);
  or csa_tree_add_51_79_groupi_g36938(csa_tree_add_51_79_groupi_n_9118 ,csa_tree_add_51_79_groupi_n_8645 ,csa_tree_add_51_79_groupi_n_8692);
  and csa_tree_add_51_79_groupi_g36939(csa_tree_add_51_79_groupi_n_9117 ,csa_tree_add_51_79_groupi_n_8738 ,csa_tree_add_51_79_groupi_n_8737);
  or csa_tree_add_51_79_groupi_g36940(csa_tree_add_51_79_groupi_n_9116 ,csa_tree_add_51_79_groupi_n_8717 ,csa_tree_add_51_79_groupi_n_8589);
  or csa_tree_add_51_79_groupi_g36941(csa_tree_add_51_79_groupi_n_9115 ,csa_tree_add_51_79_groupi_n_8641 ,csa_tree_add_51_79_groupi_n_8879);
  and csa_tree_add_51_79_groupi_g36942(csa_tree_add_51_79_groupi_n_9114 ,csa_tree_add_51_79_groupi_n_8717 ,csa_tree_add_51_79_groupi_n_8589);
  or csa_tree_add_51_79_groupi_g36943(csa_tree_add_51_79_groupi_n_9113 ,csa_tree_add_51_79_groupi_n_8497 ,csa_tree_add_51_79_groupi_n_8877);
  nor csa_tree_add_51_79_groupi_g36944(csa_tree_add_51_79_groupi_n_9112 ,csa_tree_add_51_79_groupi_n_8644 ,csa_tree_add_51_79_groupi_n_8873);
  or csa_tree_add_51_79_groupi_g36945(csa_tree_add_51_79_groupi_n_9111 ,csa_tree_add_51_79_groupi_n_8031 ,csa_tree_add_51_79_groupi_n_8707);
  or csa_tree_add_51_79_groupi_g36946(csa_tree_add_51_79_groupi_n_9110 ,csa_tree_add_51_79_groupi_n_8637 ,csa_tree_add_51_79_groupi_n_8868);
  or csa_tree_add_51_79_groupi_g36947(csa_tree_add_51_79_groupi_n_9109 ,csa_tree_add_51_79_groupi_n_8643 ,csa_tree_add_51_79_groupi_n_8848);
  or csa_tree_add_51_79_groupi_g36948(csa_tree_add_51_79_groupi_n_9108 ,csa_tree_add_51_79_groupi_n_8720 ,csa_tree_add_51_79_groupi_n_8735);
  or csa_tree_add_51_79_groupi_g36949(csa_tree_add_51_79_groupi_n_9107 ,csa_tree_add_51_79_groupi_n_8602 ,csa_tree_add_51_79_groupi_n_8745);
  and csa_tree_add_51_79_groupi_g36950(csa_tree_add_51_79_groupi_n_9106 ,csa_tree_add_51_79_groupi_n_8720 ,csa_tree_add_51_79_groupi_n_8735);
  or csa_tree_add_51_79_groupi_g36951(csa_tree_add_51_79_groupi_n_9105 ,csa_tree_add_51_79_groupi_n_8486 ,csa_tree_add_51_79_groupi_n_8871);
  nor csa_tree_add_51_79_groupi_g36952(csa_tree_add_51_79_groupi_n_9104 ,csa_tree_add_51_79_groupi_n_8603 ,csa_tree_add_51_79_groupi_n_8746);
  or csa_tree_add_51_79_groupi_g36953(csa_tree_add_51_79_groupi_n_9103 ,csa_tree_add_51_79_groupi_n_8869 ,csa_tree_add_51_79_groupi_n_8801);
  or csa_tree_add_51_79_groupi_g36954(csa_tree_add_51_79_groupi_n_9102 ,csa_tree_add_51_79_groupi_n_8490 ,csa_tree_add_51_79_groupi_n_8850);
  and csa_tree_add_51_79_groupi_g36955(csa_tree_add_51_79_groupi_n_9101 ,csa_tree_add_51_79_groupi_n_8722 ,csa_tree_add_51_79_groupi_n_8721);
  or csa_tree_add_51_79_groupi_g36956(csa_tree_add_51_79_groupi_n_9100 ,csa_tree_add_51_79_groupi_n_8722 ,csa_tree_add_51_79_groupi_n_8721);
  nor csa_tree_add_51_79_groupi_g36957(csa_tree_add_51_79_groupi_n_9099 ,csa_tree_add_51_79_groupi_n_7591 ,csa_tree_add_51_79_groupi_n_8777);
  and csa_tree_add_51_79_groupi_g36958(csa_tree_add_51_79_groupi_n_9098 ,csa_tree_add_51_79_groupi_n_8958 ,csa_tree_add_51_79_groupi_n_8960);
  nor csa_tree_add_51_79_groupi_g36959(csa_tree_add_51_79_groupi_n_9097 ,csa_tree_add_51_79_groupi_n_8728 ,csa_tree_add_51_79_groupi_n_8731);
  or csa_tree_add_51_79_groupi_g36960(csa_tree_add_51_79_groupi_n_9096 ,csa_tree_add_51_79_groupi_n_8727 ,csa_tree_add_51_79_groupi_n_8732);
  or csa_tree_add_51_79_groupi_g36961(csa_tree_add_51_79_groupi_n_9095 ,csa_tree_add_51_79_groupi_n_8335 ,csa_tree_add_51_79_groupi_n_8844);
  and csa_tree_add_51_79_groupi_g36962(csa_tree_add_51_79_groupi_n_9094 ,csa_tree_add_51_79_groupi_n_8452 ,csa_tree_add_51_79_groupi_n_8793);
  or csa_tree_add_51_79_groupi_g36963(csa_tree_add_51_79_groupi_n_9093 ,csa_tree_add_51_79_groupi_n_8252 ,csa_tree_add_51_79_groupi_n_8820);
  or csa_tree_add_51_79_groupi_g36964(csa_tree_add_51_79_groupi_n_9092 ,csa_tree_add_51_79_groupi_n_7592 ,csa_tree_add_51_79_groupi_n_8776);
  or csa_tree_add_51_79_groupi_g36965(csa_tree_add_51_79_groupi_n_9091 ,csa_tree_add_51_79_groupi_n_8624 ,csa_tree_add_51_79_groupi_n_8860);
  or csa_tree_add_51_79_groupi_g36966(csa_tree_add_51_79_groupi_n_9090 ,csa_tree_add_51_79_groupi_n_8726 ,csa_tree_add_51_79_groupi_n_8760);
  and csa_tree_add_51_79_groupi_g36967(csa_tree_add_51_79_groupi_n_9089 ,csa_tree_add_51_79_groupi_n_8726 ,csa_tree_add_51_79_groupi_n_8760);
  nor csa_tree_add_51_79_groupi_g36968(csa_tree_add_51_79_groupi_n_9088 ,csa_tree_add_51_79_groupi_n_8958 ,csa_tree_add_51_79_groupi_n_8960);
  nor csa_tree_add_51_79_groupi_g36969(csa_tree_add_51_79_groupi_n_9087 ,csa_tree_add_51_79_groupi_n_8452 ,csa_tree_add_51_79_groupi_n_8793);
  and csa_tree_add_51_79_groupi_g36970(csa_tree_add_51_79_groupi_n_9206 ,csa_tree_add_51_79_groupi_n_8555 ,csa_tree_add_51_79_groupi_n_8837);
  and csa_tree_add_51_79_groupi_g36971(csa_tree_add_51_79_groupi_n_9205 ,csa_tree_add_51_79_groupi_n_8538 ,csa_tree_add_51_79_groupi_n_8854);
  and csa_tree_add_51_79_groupi_g36972(csa_tree_add_51_79_groupi_n_9204 ,csa_tree_add_51_79_groupi_n_8516 ,csa_tree_add_51_79_groupi_n_8867);
  and csa_tree_add_51_79_groupi_g36973(csa_tree_add_51_79_groupi_n_9203 ,csa_tree_add_51_79_groupi_n_8548 ,csa_tree_add_51_79_groupi_n_8915);
  and csa_tree_add_51_79_groupi_g36974(csa_tree_add_51_79_groupi_n_9202 ,csa_tree_add_51_79_groupi_n_8521 ,csa_tree_add_51_79_groupi_n_8912);
  and csa_tree_add_51_79_groupi_g36975(csa_tree_add_51_79_groupi_n_9201 ,csa_tree_add_51_79_groupi_n_8540 ,csa_tree_add_51_79_groupi_n_8853);
  and csa_tree_add_51_79_groupi_g36976(csa_tree_add_51_79_groupi_n_9200 ,csa_tree_add_51_79_groupi_n_8522 ,csa_tree_add_51_79_groupi_n_8913);
  and csa_tree_add_51_79_groupi_g36977(csa_tree_add_51_79_groupi_n_9199 ,csa_tree_add_51_79_groupi_n_8542 ,csa_tree_add_51_79_groupi_n_8931);
  and csa_tree_add_51_79_groupi_g36978(csa_tree_add_51_79_groupi_n_9198 ,csa_tree_add_51_79_groupi_n_8546 ,csa_tree_add_51_79_groupi_n_8932);
  and csa_tree_add_51_79_groupi_g36979(csa_tree_add_51_79_groupi_n_9197 ,csa_tree_add_51_79_groupi_n_8563 ,csa_tree_add_51_79_groupi_n_8950);
  and csa_tree_add_51_79_groupi_g36980(csa_tree_add_51_79_groupi_n_9196 ,csa_tree_add_51_79_groupi_n_8357 ,csa_tree_add_51_79_groupi_n_8952);
  and csa_tree_add_51_79_groupi_g36981(csa_tree_add_51_79_groupi_n_9195 ,csa_tree_add_51_79_groupi_n_8509 ,csa_tree_add_51_79_groupi_n_8890);
  and csa_tree_add_51_79_groupi_g36982(csa_tree_add_51_79_groupi_n_9194 ,csa_tree_add_51_79_groupi_n_8507 ,csa_tree_add_51_79_groupi_n_8900);
  and csa_tree_add_51_79_groupi_g36983(csa_tree_add_51_79_groupi_n_9193 ,csa_tree_add_51_79_groupi_n_8508 ,csa_tree_add_51_79_groupi_n_8892);
  and csa_tree_add_51_79_groupi_g36984(csa_tree_add_51_79_groupi_n_9191 ,csa_tree_add_51_79_groupi_n_8524 ,csa_tree_add_51_79_groupi_n_8914);
  and csa_tree_add_51_79_groupi_g36985(csa_tree_add_51_79_groupi_n_9190 ,csa_tree_add_51_79_groupi_n_8530 ,csa_tree_add_51_79_groupi_n_8858);
  and csa_tree_add_51_79_groupi_g36986(csa_tree_add_51_79_groupi_n_9189 ,csa_tree_add_51_79_groupi_n_8554 ,csa_tree_add_51_79_groupi_n_8838);
  and csa_tree_add_51_79_groupi_g36987(csa_tree_add_51_79_groupi_n_9188 ,csa_tree_add_51_79_groupi_n_8533 ,csa_tree_add_51_79_groupi_n_8857);
  or csa_tree_add_51_79_groupi_g36988(csa_tree_add_51_79_groupi_n_9186 ,csa_tree_add_51_79_groupi_n_8520 ,csa_tree_add_51_79_groupi_n_8886);
  and csa_tree_add_51_79_groupi_g36989(csa_tree_add_51_79_groupi_n_9185 ,csa_tree_add_51_79_groupi_n_8237 ,csa_tree_add_51_79_groupi_n_8864);
  and csa_tree_add_51_79_groupi_g36990(csa_tree_add_51_79_groupi_n_9182 ,csa_tree_add_51_79_groupi_n_8534 ,csa_tree_add_51_79_groupi_n_8956);
  and csa_tree_add_51_79_groupi_g36991(csa_tree_add_51_79_groupi_n_9181 ,csa_tree_add_51_79_groupi_n_8515 ,csa_tree_add_51_79_groupi_n_8865);
  and csa_tree_add_51_79_groupi_g36992(csa_tree_add_51_79_groupi_n_9180 ,csa_tree_add_51_79_groupi_n_8552 ,csa_tree_add_51_79_groupi_n_8942);
  and csa_tree_add_51_79_groupi_g36993(csa_tree_add_51_79_groupi_n_9179 ,csa_tree_add_51_79_groupi_n_8558 ,csa_tree_add_51_79_groupi_n_8944);
  or csa_tree_add_51_79_groupi_g36994(csa_tree_add_51_79_groupi_n_9178 ,csa_tree_add_51_79_groupi_n_8519 ,csa_tree_add_51_79_groupi_n_8916);
  and csa_tree_add_51_79_groupi_g36995(csa_tree_add_51_79_groupi_n_9176 ,csa_tree_add_51_79_groupi_n_8366 ,csa_tree_add_51_79_groupi_n_8891);
  and csa_tree_add_51_79_groupi_g36996(csa_tree_add_51_79_groupi_n_9175 ,csa_tree_add_51_79_groupi_n_8562 ,csa_tree_add_51_79_groupi_n_8947);
  not csa_tree_add_51_79_groupi_g36997(csa_tree_add_51_79_groupi_n_9077 ,csa_tree_add_51_79_groupi_n_9076);
  not csa_tree_add_51_79_groupi_g36998(csa_tree_add_51_79_groupi_n_9075 ,csa_tree_add_51_79_groupi_n_9074);
  and csa_tree_add_51_79_groupi_g36999(csa_tree_add_51_79_groupi_n_9068 ,csa_tree_add_51_79_groupi_n_8959 ,csa_tree_add_51_79_groupi_n_8423);
  or csa_tree_add_51_79_groupi_g37000(csa_tree_add_51_79_groupi_n_9067 ,csa_tree_add_51_79_groupi_n_8639 ,csa_tree_add_51_79_groupi_n_8831);
  or csa_tree_add_51_79_groupi_g37001(csa_tree_add_51_79_groupi_n_9066 ,csa_tree_add_51_79_groupi_n_8743 ,csa_tree_add_51_79_groupi_n_8741);
  and csa_tree_add_51_79_groupi_g37002(csa_tree_add_51_79_groupi_n_9065 ,csa_tree_add_51_79_groupi_n_8743 ,csa_tree_add_51_79_groupi_n_8741);
  or csa_tree_add_51_79_groupi_g37003(csa_tree_add_51_79_groupi_n_9064 ,csa_tree_add_51_79_groupi_n_8736 ,csa_tree_add_51_79_groupi_n_8734);
  and csa_tree_add_51_79_groupi_g37004(csa_tree_add_51_79_groupi_n_9063 ,csa_tree_add_51_79_groupi_n_8736 ,csa_tree_add_51_79_groupi_n_8734);
  or csa_tree_add_51_79_groupi_g37005(csa_tree_add_51_79_groupi_n_9062 ,csa_tree_add_51_79_groupi_n_8730 ,csa_tree_add_51_79_groupi_n_8729);
  and csa_tree_add_51_79_groupi_g37006(csa_tree_add_51_79_groupi_n_9061 ,csa_tree_add_51_79_groupi_n_8730 ,csa_tree_add_51_79_groupi_n_8729);
  or csa_tree_add_51_79_groupi_g37007(csa_tree_add_51_79_groupi_n_9060 ,csa_tree_add_51_79_groupi_n_8778 ,csa_tree_add_51_79_groupi_n_8794);
  and csa_tree_add_51_79_groupi_g37008(csa_tree_add_51_79_groupi_n_9059 ,csa_tree_add_51_79_groupi_n_8778 ,csa_tree_add_51_79_groupi_n_8794);
  or csa_tree_add_51_79_groupi_g37009(csa_tree_add_51_79_groupi_n_9058 ,csa_tree_add_51_79_groupi_n_8501 ,csa_tree_add_51_79_groupi_n_8827);
  or csa_tree_add_51_79_groupi_g37010(csa_tree_add_51_79_groupi_n_9057 ,csa_tree_add_51_79_groupi_n_8825 ,csa_tree_add_51_79_groupi_n_8815);
  or csa_tree_add_51_79_groupi_g37011(csa_tree_add_51_79_groupi_n_9056 ,csa_tree_add_51_79_groupi_n_8786 ,csa_tree_add_51_79_groupi_n_8785);
  and csa_tree_add_51_79_groupi_g37012(csa_tree_add_51_79_groupi_n_9055 ,csa_tree_add_51_79_groupi_n_8786 ,csa_tree_add_51_79_groupi_n_8785);
  or csa_tree_add_51_79_groupi_g37013(csa_tree_add_51_79_groupi_n_9054 ,csa_tree_add_51_79_groupi_n_8780 ,csa_tree_add_51_79_groupi_n_8779);
  and csa_tree_add_51_79_groupi_g37014(csa_tree_add_51_79_groupi_n_9053 ,csa_tree_add_51_79_groupi_n_8780 ,csa_tree_add_51_79_groupi_n_8779);
  or csa_tree_add_51_79_groupi_g37015(csa_tree_add_51_79_groupi_n_9052 ,csa_tree_add_51_79_groupi_n_8498 ,csa_tree_add_51_79_groupi_n_8859);
  or csa_tree_add_51_79_groupi_g37016(csa_tree_add_51_79_groupi_n_9051 ,csa_tree_add_51_79_groupi_n_8488 ,csa_tree_add_51_79_groupi_n_8863);
  or csa_tree_add_51_79_groupi_g37017(csa_tree_add_51_79_groupi_n_9050 ,csa_tree_add_51_79_groupi_n_8638 ,csa_tree_add_51_79_groupi_n_8875);
  or csa_tree_add_51_79_groupi_g37018(csa_tree_add_51_79_groupi_n_9049 ,csa_tree_add_51_79_groupi_n_8494 ,csa_tree_add_51_79_groupi_n_8909);
  or csa_tree_add_51_79_groupi_g37019(csa_tree_add_51_79_groupi_n_9048 ,csa_tree_add_51_79_groupi_n_8772 ,csa_tree_add_51_79_groupi_n_8771);
  and csa_tree_add_51_79_groupi_g37020(csa_tree_add_51_79_groupi_n_9047 ,csa_tree_add_51_79_groupi_n_8772 ,csa_tree_add_51_79_groupi_n_8771);
  or csa_tree_add_51_79_groupi_g37021(csa_tree_add_51_79_groupi_n_9046 ,csa_tree_add_51_79_groupi_n_8500 ,csa_tree_add_51_79_groupi_n_8876);
  or csa_tree_add_51_79_groupi_g37022(csa_tree_add_51_79_groupi_n_9045 ,csa_tree_add_51_79_groupi_n_8632 ,csa_tree_add_51_79_groupi_n_8907);
  or csa_tree_add_51_79_groupi_g37023(csa_tree_add_51_79_groupi_n_9044 ,csa_tree_add_51_79_groupi_n_7832 ,csa_tree_add_51_79_groupi_n_8954);
  or csa_tree_add_51_79_groupi_g37024(csa_tree_add_51_79_groupi_n_9043 ,csa_tree_add_51_79_groupi_n_8605 ,csa_tree_add_51_79_groupi_n_8789);
  nor csa_tree_add_51_79_groupi_g37025(csa_tree_add_51_79_groupi_n_9042 ,csa_tree_add_51_79_groupi_n_8606 ,csa_tree_add_51_79_groupi_n_8790);
  or csa_tree_add_51_79_groupi_g37026(csa_tree_add_51_79_groupi_n_9041 ,csa_tree_add_51_79_groupi_n_8636 ,csa_tree_add_51_79_groupi_n_8855);
  or csa_tree_add_51_79_groupi_g37027(csa_tree_add_51_79_groupi_n_9040 ,csa_tree_add_51_79_groupi_n_8504 ,csa_tree_add_51_79_groupi_n_8905);
  or csa_tree_add_51_79_groupi_g37028(csa_tree_add_51_79_groupi_n_9039 ,csa_tree_add_51_79_groupi_n_8502 ,csa_tree_add_51_79_groupi_n_8713);
  or csa_tree_add_51_79_groupi_g37029(csa_tree_add_51_79_groupi_n_9038 ,csa_tree_add_51_79_groupi_n_8185 ,csa_tree_add_51_79_groupi_n_8711);
  or csa_tree_add_51_79_groupi_g37030(csa_tree_add_51_79_groupi_n_9037 ,csa_tree_add_51_79_groupi_n_8030 ,csa_tree_add_51_79_groupi_n_8703);
  or csa_tree_add_51_79_groupi_g37031(csa_tree_add_51_79_groupi_n_9036 ,csa_tree_add_51_79_groupi_n_8178 ,csa_tree_add_51_79_groupi_n_8709);
  nor csa_tree_add_51_79_groupi_g37032(csa_tree_add_51_79_groupi_n_9035 ,csa_tree_add_51_79_groupi_n_8491 ,csa_tree_add_51_79_groupi_n_8920);
  and csa_tree_add_51_79_groupi_g37033(csa_tree_add_51_79_groupi_n_9034 ,csa_tree_add_51_79_groupi_n_8965 ,csa_tree_add_51_79_groupi_n_8704);
  or csa_tree_add_51_79_groupi_g37034(csa_tree_add_51_79_groupi_n_9033 ,csa_tree_add_51_79_groupi_n_8701 ,csa_tree_add_51_79_groupi_n_8821);
  or csa_tree_add_51_79_groupi_g37035(csa_tree_add_51_79_groupi_n_9032 ,csa_tree_add_51_79_groupi_n_8627 ,csa_tree_add_51_79_groupi_n_8700);
  or csa_tree_add_51_79_groupi_g37036(csa_tree_add_51_79_groupi_n_9031 ,csa_tree_add_51_79_groupi_n_8657 ,csa_tree_add_51_79_groupi_n_8943);
  xor csa_tree_add_51_79_groupi_g37037(csa_tree_add_51_79_groupi_n_9030 ,csa_tree_add_51_79_groupi_n_8625 ,csa_tree_add_51_79_groupi_n_8615);
  xnor csa_tree_add_51_79_groupi_g37038(csa_tree_add_51_79_groupi_n_9029 ,csa_tree_add_51_79_groupi_n_8596 ,csa_tree_add_51_79_groupi_n_8640);
  xnor csa_tree_add_51_79_groupi_g37039(csa_tree_add_51_79_groupi_n_9028 ,csa_tree_add_51_79_groupi_n_8650 ,csa_tree_add_51_79_groupi_n_8588);
  xnor csa_tree_add_51_79_groupi_g37040(csa_tree_add_51_79_groupi_n_9027 ,csa_tree_add_51_79_groupi_n_8459 ,csa_tree_add_51_79_groupi_n_8391);
  xnor csa_tree_add_51_79_groupi_g37041(csa_tree_add_51_79_groupi_n_9026 ,csa_tree_add_51_79_groupi_n_8578 ,csa_tree_add_51_79_groupi_n_8584);
  xnor csa_tree_add_51_79_groupi_g37042(csa_tree_add_51_79_groupi_n_9025 ,csa_tree_add_51_79_groupi_n_8581 ,csa_tree_add_51_79_groupi_n_8655);
  xnor csa_tree_add_51_79_groupi_g37043(csa_tree_add_51_79_groupi_n_9024 ,csa_tree_add_51_79_groupi_n_8464 ,csa_tree_add_51_79_groupi_n_8396);
  xnor csa_tree_add_51_79_groupi_g37044(csa_tree_add_51_79_groupi_n_9023 ,csa_tree_add_51_79_groupi_n_8613 ,csa_tree_add_51_79_groupi_n_8477);
  xnor csa_tree_add_51_79_groupi_g37045(csa_tree_add_51_79_groupi_n_9022 ,csa_tree_add_51_79_groupi_n_8304 ,csa_tree_add_51_79_groupi_n_8632);
  xnor csa_tree_add_51_79_groupi_g37046(csa_tree_add_51_79_groupi_n_9021 ,csa_tree_add_51_79_groupi_n_8165 ,csa_tree_add_51_79_groupi_n_8414);
  xnor csa_tree_add_51_79_groupi_g37047(csa_tree_add_51_79_groupi_n_9020 ,csa_tree_add_51_79_groupi_n_8377 ,csa_tree_add_51_79_groupi_n_8417);
  xnor csa_tree_add_51_79_groupi_g37048(csa_tree_add_51_79_groupi_n_9019 ,csa_tree_add_51_79_groupi_n_8381 ,csa_tree_add_51_79_groupi_n_8460);
  xnor csa_tree_add_51_79_groupi_g37049(csa_tree_add_51_79_groupi_n_9018 ,csa_tree_add_51_79_groupi_n_8620 ,csa_tree_add_51_79_groupi_n_8626);
  xnor csa_tree_add_51_79_groupi_g37050(csa_tree_add_51_79_groupi_n_9017 ,csa_tree_add_51_79_groupi_n_8387 ,csa_tree_add_51_79_groupi_n_8389);
  xnor csa_tree_add_51_79_groupi_g37051(csa_tree_add_51_79_groupi_n_9016 ,csa_tree_add_51_79_groupi_n_8598 ,csa_tree_add_51_79_groupi_n_8383);
  xnor csa_tree_add_51_79_groupi_g37052(csa_tree_add_51_79_groupi_n_9015 ,csa_tree_add_51_79_groupi_n_8643 ,csa_tree_add_51_79_groupi_n_8451);
  xnor csa_tree_add_51_79_groupi_g37053(csa_tree_add_51_79_groupi_n_9014 ,csa_tree_add_51_79_groupi_n_8438 ,csa_tree_add_51_79_groupi_n_8636);
  xnor csa_tree_add_51_79_groupi_g37054(csa_tree_add_51_79_groupi_n_9013 ,csa_tree_add_51_79_groupi_n_8418 ,csa_tree_add_51_79_groupi_n_8635);
  xnor csa_tree_add_51_79_groupi_g37056(csa_tree_add_51_79_groupi_n_9012 ,csa_tree_add_51_79_groupi_n_8472 ,csa_tree_add_51_79_groupi_n_8020);
  xnor csa_tree_add_51_79_groupi_g37057(csa_tree_add_51_79_groupi_n_9011 ,csa_tree_add_51_79_groupi_n_8600 ,csa_tree_add_51_79_groupi_n_8609);
  xnor csa_tree_add_51_79_groupi_g37058(csa_tree_add_51_79_groupi_n_9010 ,csa_tree_add_51_79_groupi_n_8482 ,csa_tree_add_51_79_groupi_n_8651);
  xnor csa_tree_add_51_79_groupi_g37059(csa_tree_add_51_79_groupi_n_9009 ,csa_tree_add_51_79_groupi_n_8401 ,csa_tree_add_51_79_groupi_n_8491);
  xnor csa_tree_add_51_79_groupi_g37060(csa_tree_add_51_79_groupi_n_9008 ,csa_tree_add_51_79_groupi_n_8586 ,csa_tree_add_51_79_groupi_n_8645);
  xnor csa_tree_add_51_79_groupi_g37061(csa_tree_add_51_79_groupi_n_9007 ,csa_tree_add_51_79_groupi_n_8159 ,csa_tree_add_51_79_groupi_n_8380);
  xnor csa_tree_add_51_79_groupi_g37062(csa_tree_add_51_79_groupi_n_9006 ,csa_tree_add_51_79_groupi_n_8415 ,csa_tree_add_51_79_groupi_n_8176);
  xnor csa_tree_add_51_79_groupi_g37063(csa_tree_add_51_79_groupi_n_9005 ,csa_tree_add_51_79_groupi_n_8461 ,csa_tree_add_51_79_groupi_n_7806);
  xnor csa_tree_add_51_79_groupi_g37064(csa_tree_add_51_79_groupi_n_9004 ,csa_tree_add_51_79_groupi_n_8462 ,csa_tree_add_51_79_groupi_n_8286);
  xnor csa_tree_add_51_79_groupi_g37065(csa_tree_add_51_79_groupi_n_9003 ,csa_tree_add_51_79_groupi_n_8641 ,csa_tree_add_51_79_groupi_n_8467);
  xnor csa_tree_add_51_79_groupi_g37066(csa_tree_add_51_79_groupi_n_9002 ,csa_tree_add_51_79_groupi_n_8030 ,csa_tree_add_51_79_groupi_n_8455);
  xnor csa_tree_add_51_79_groupi_g37067(csa_tree_add_51_79_groupi_n_9001 ,csa_tree_add_51_79_groupi_n_8324 ,csa_tree_add_51_79_groupi_n_8449);
  xnor csa_tree_add_51_79_groupi_g37068(csa_tree_add_51_79_groupi_n_9000 ,csa_tree_add_51_79_groupi_n_8616 ,csa_tree_add_51_79_groupi_n_26);
  xnor csa_tree_add_51_79_groupi_g37069(csa_tree_add_51_79_groupi_n_8999 ,csa_tree_add_51_79_groupi_n_8428 ,csa_tree_add_51_79_groupi_n_8429);
  xnor csa_tree_add_51_79_groupi_g37070(csa_tree_add_51_79_groupi_n_8998 ,csa_tree_add_51_79_groupi_n_8572 ,csa_tree_add_51_79_groupi_n_8447);
  xnor csa_tree_add_51_79_groupi_g37071(csa_tree_add_51_79_groupi_n_8997 ,csa_tree_add_51_79_groupi_n_8638 ,csa_tree_add_51_79_groupi_n_8607);
  xnor csa_tree_add_51_79_groupi_g37072(csa_tree_add_51_79_groupi_n_8996 ,csa_tree_add_51_79_groupi_n_8648 ,csa_tree_add_51_79_groupi_n_8590);
  xnor csa_tree_add_51_79_groupi_g37073(csa_tree_add_51_79_groupi_n_8995 ,csa_tree_add_51_79_groupi_n_8567 ,csa_tree_add_51_79_groupi_n_8475);
  xnor csa_tree_add_51_79_groupi_g37074(csa_tree_add_51_79_groupi_n_8994 ,csa_tree_add_51_79_groupi_n_8593 ,csa_tree_add_51_79_groupi_n_8506);
  xnor csa_tree_add_51_79_groupi_g37075(csa_tree_add_51_79_groupi_n_8993 ,csa_tree_add_51_79_groupi_n_8427 ,csa_tree_add_51_79_groupi_n_8444);
  xnor csa_tree_add_51_79_groupi_g37076(csa_tree_add_51_79_groupi_n_8992 ,csa_tree_add_51_79_groupi_n_8410 ,csa_tree_add_51_79_groupi_n_8445);
  xnor csa_tree_add_51_79_groupi_g37077(csa_tree_add_51_79_groupi_n_8991 ,csa_tree_add_51_79_groupi_n_8579 ,csa_tree_add_51_79_groupi_n_8426);
  xnor csa_tree_add_51_79_groupi_g37078(csa_tree_add_51_79_groupi_n_8990 ,csa_tree_add_51_79_groupi_n_8425 ,csa_tree_add_51_79_groupi_n_8404);
  xnor csa_tree_add_51_79_groupi_g37079(csa_tree_add_51_79_groupi_n_8989 ,csa_tree_add_51_79_groupi_n_8594 ,csa_tree_add_51_79_groupi_n_8623);
  xnor csa_tree_add_51_79_groupi_g37080(csa_tree_add_51_79_groupi_n_8988 ,csa_tree_add_51_79_groupi_n_8443 ,csa_tree_add_51_79_groupi_n_8270);
  xnor csa_tree_add_51_79_groupi_g37081(csa_tree_add_51_79_groupi_n_8987 ,csa_tree_add_51_79_groupi_n_8611 ,csa_tree_add_51_79_groupi_n_8378);
  xnor csa_tree_add_51_79_groupi_g37082(csa_tree_add_51_79_groupi_n_8986 ,csa_tree_add_51_79_groupi_n_8424 ,csa_tree_add_51_79_groupi_n_8399);
  xnor csa_tree_add_51_79_groupi_g37083(csa_tree_add_51_79_groupi_n_8985 ,csa_tree_add_51_79_groupi_n_8421 ,csa_tree_add_51_79_groupi_n_8498);
  xnor csa_tree_add_51_79_groupi_g37084(csa_tree_add_51_79_groupi_n_8984 ,csa_tree_add_51_79_groupi_n_8501 ,csa_tree_add_51_79_groupi_n_8435);
  xnor csa_tree_add_51_79_groupi_g37085(csa_tree_add_51_79_groupi_n_8983 ,csa_tree_add_51_79_groupi_n_8474 ,csa_tree_add_51_79_groupi_n_8157);
  xnor csa_tree_add_51_79_groupi_g37086(csa_tree_add_51_79_groupi_n_8982 ,csa_tree_add_51_79_groupi_n_8393 ,csa_tree_add_51_79_groupi_n_8440);
  xnor csa_tree_add_51_79_groupi_g37087(csa_tree_add_51_79_groupi_n_8981 ,csa_tree_add_51_79_groupi_n_8439 ,csa_tree_add_51_79_groupi_n_8392);
  xnor csa_tree_add_51_79_groupi_g37088(csa_tree_add_51_79_groupi_n_8980 ,csa_tree_add_51_79_groupi_n_8384 ,csa_tree_add_51_79_groupi_n_8497);
  xnor csa_tree_add_51_79_groupi_g37089(csa_tree_add_51_79_groupi_n_8979 ,csa_tree_add_51_79_groupi_n_8422 ,csa_tree_add_51_79_groupi_n_8582);
  xnor csa_tree_add_51_79_groupi_g37090(csa_tree_add_51_79_groupi_n_8978 ,csa_tree_add_51_79_groupi_n_8430 ,csa_tree_add_51_79_groupi_n_8488);
  xnor csa_tree_add_51_79_groupi_g37091(csa_tree_add_51_79_groupi_n_8977 ,csa_tree_add_51_79_groupi_n_8495 ,csa_tree_add_51_79_groupi_n_8155);
  xnor csa_tree_add_51_79_groupi_g37092(csa_tree_add_51_79_groupi_n_8976 ,csa_tree_add_51_79_groupi_n_8433 ,csa_tree_add_51_79_groupi_n_8335);
  xnor csa_tree_add_51_79_groupi_g37093(csa_tree_add_51_79_groupi_n_8975 ,csa_tree_add_51_79_groupi_n_8373 ,csa_tree_add_51_79_groupi_n_8269);
  xnor csa_tree_add_51_79_groupi_g37094(csa_tree_add_51_79_groupi_n_8974 ,csa_tree_add_51_79_groupi_n_8569 ,csa_tree_add_51_79_groupi_n_8624);
  xor csa_tree_add_51_79_groupi_g37095(csa_tree_add_51_79_groupi_n_8973 ,csa_tree_add_51_79_groupi_n_8644 ,csa_tree_add_51_79_groupi_n_8446);
  xnor csa_tree_add_51_79_groupi_g37096(csa_tree_add_51_79_groupi_n_8972 ,csa_tree_add_51_79_groupi_n_8610 ,csa_tree_add_51_79_groupi_n_8601);
  xnor csa_tree_add_51_79_groupi_g37097(csa_tree_add_51_79_groupi_n_8971 ,csa_tree_add_51_79_groupi_n_8394 ,csa_tree_add_51_79_groupi_n_8334);
  and csa_tree_add_51_79_groupi_g37098(csa_tree_add_51_79_groupi_n_9086 ,csa_tree_add_51_79_groupi_n_8362 ,csa_tree_add_51_79_groupi_n_8706);
  xnor csa_tree_add_51_79_groupi_g37099(csa_tree_add_51_79_groupi_n_9085 ,csa_tree_add_51_79_groupi_n_8272 ,csa_tree_add_51_79_groupi_n_8345);
  xnor csa_tree_add_51_79_groupi_g37100(csa_tree_add_51_79_groupi_n_9084 ,csa_tree_add_51_79_groupi_n_7833 ,csa_tree_add_51_79_groupi_n_8353);
  xnor csa_tree_add_51_79_groupi_g37101(csa_tree_add_51_79_groupi_n_9083 ,csa_tree_add_51_79_groupi_n_8448 ,csa_tree_add_51_79_groupi_n_8347);
  xnor csa_tree_add_51_79_groupi_g37102(csa_tree_add_51_79_groupi_n_9082 ,csa_tree_add_51_79_groupi_n_8492 ,csa_tree_add_51_79_groupi_n_8355);
  and csa_tree_add_51_79_groupi_g37103(csa_tree_add_51_79_groupi_n_9081 ,csa_tree_add_51_79_groupi_n_8368 ,csa_tree_add_51_79_groupi_n_8716);
  xnor csa_tree_add_51_79_groupi_g37104(csa_tree_add_51_79_groupi_n_9080 ,csa_tree_add_51_79_groupi_n_7204 ,csa_tree_add_51_79_groupi_n_8352);
  xnor csa_tree_add_51_79_groupi_g37105(csa_tree_add_51_79_groupi_n_9079 ,csa_tree_add_51_79_groupi_n_8179 ,csa_tree_add_51_79_groupi_n_8346);
  xnor csa_tree_add_51_79_groupi_g37106(csa_tree_add_51_79_groupi_n_9078 ,csa_tree_add_51_79_groupi_n_8322 ,csa_tree_add_51_79_groupi_n_8350);
  xnor csa_tree_add_51_79_groupi_g37107(csa_tree_add_51_79_groupi_n_9076 ,csa_tree_add_51_79_groupi_n_7372 ,csa_tree_add_51_79_groupi_n_8349);
  xnor csa_tree_add_51_79_groupi_g37108(csa_tree_add_51_79_groupi_n_9074 ,csa_tree_add_51_79_groupi_n_7822 ,csa_tree_add_51_79_groupi_n_8351);
  and csa_tree_add_51_79_groupi_g37109(csa_tree_add_51_79_groupi_n_9073 ,csa_tree_add_51_79_groupi_n_8364 ,csa_tree_add_51_79_groupi_n_8715);
  xnor csa_tree_add_51_79_groupi_g37110(csa_tree_add_51_79_groupi_n_9072 ,csa_tree_add_51_79_groupi_n_7826 ,csa_tree_add_51_79_groupi_n_8348);
  xnor csa_tree_add_51_79_groupi_g37111(csa_tree_add_51_79_groupi_n_9071 ,csa_tree_add_51_79_groupi_n_7170 ,csa_tree_add_51_79_groupi_n_8356);
  xnor csa_tree_add_51_79_groupi_g37112(csa_tree_add_51_79_groupi_n_9070 ,csa_tree_add_51_79_groupi_n_7230 ,csa_tree_add_51_79_groupi_n_8354);
  or csa_tree_add_51_79_groupi_g37113(csa_tree_add_51_79_groupi_n_9069 ,csa_tree_add_51_79_groupi_n_8358 ,csa_tree_add_51_79_groupi_n_8698);
  not csa_tree_add_51_79_groupi_g37115(csa_tree_add_51_79_groupi_n_8962 ,csa_tree_add_51_79_groupi_n_8961);
  and csa_tree_add_51_79_groupi_g37116(csa_tree_add_51_79_groupi_n_8957 ,csa_tree_add_51_79_groupi_n_8446 ,csa_tree_add_51_79_groupi_n_8442);
  or csa_tree_add_51_79_groupi_g37117(csa_tree_add_51_79_groupi_n_8956 ,csa_tree_add_51_79_groupi_n_8312 ,csa_tree_add_51_79_groupi_n_8561);
  or csa_tree_add_51_79_groupi_g37118(csa_tree_add_51_79_groupi_n_8955 ,csa_tree_add_51_79_groupi_n_8447 ,csa_tree_add_51_79_groupi_n_8572);
  and csa_tree_add_51_79_groupi_g37119(csa_tree_add_51_79_groupi_n_8954 ,csa_tree_add_51_79_groupi_n_7810 ,csa_tree_add_51_79_groupi_n_8448);
  and csa_tree_add_51_79_groupi_g37120(csa_tree_add_51_79_groupi_n_8953 ,csa_tree_add_51_79_groupi_n_8447 ,csa_tree_add_51_79_groupi_n_8572);
  or csa_tree_add_51_79_groupi_g37121(csa_tree_add_51_79_groupi_n_8952 ,csa_tree_add_51_79_groupi_n_7340 ,csa_tree_add_51_79_groupi_n_8369);
  or csa_tree_add_51_79_groupi_g37122(csa_tree_add_51_79_groupi_n_8951 ,csa_tree_add_51_79_groupi_n_7810 ,csa_tree_add_51_79_groupi_n_8448);
  or csa_tree_add_51_79_groupi_g37123(csa_tree_add_51_79_groupi_n_8950 ,csa_tree_add_51_79_groupi_n_8560 ,csa_tree_add_51_79_groupi_n_8658);
  and csa_tree_add_51_79_groupi_g37124(csa_tree_add_51_79_groupi_n_8949 ,csa_tree_add_51_79_groupi_n_26 ,csa_tree_add_51_79_groupi_n_8616);
  or csa_tree_add_51_79_groupi_g37125(csa_tree_add_51_79_groupi_n_8948 ,csa_tree_add_51_79_groupi_n_26 ,csa_tree_add_51_79_groupi_n_8616);
  or csa_tree_add_51_79_groupi_g37126(csa_tree_add_51_79_groupi_n_8947 ,csa_tree_add_51_79_groupi_n_8318 ,csa_tree_add_51_79_groupi_n_8557);
  or csa_tree_add_51_79_groupi_g37127(csa_tree_add_51_79_groupi_n_8946 ,csa_tree_add_51_79_groupi_n_8291 ,csa_tree_add_51_79_groupi_n_8388);
  or csa_tree_add_51_79_groupi_g37128(csa_tree_add_51_79_groupi_n_8945 ,csa_tree_add_51_79_groupi_n_8570 ,csa_tree_add_51_79_groupi_n_8412);
  or csa_tree_add_51_79_groupi_g37129(csa_tree_add_51_79_groupi_n_8944 ,csa_tree_add_51_79_groupi_n_8320 ,csa_tree_add_51_79_groupi_n_8553);
  nor csa_tree_add_51_79_groupi_g37130(csa_tree_add_51_79_groupi_n_8943 ,csa_tree_add_51_79_groupi_n_8571 ,csa_tree_add_51_79_groupi_n_8411);
  or csa_tree_add_51_79_groupi_g37131(csa_tree_add_51_79_groupi_n_8942 ,csa_tree_add_51_79_groupi_n_8177 ,csa_tree_add_51_79_groupi_n_8550);
  or csa_tree_add_51_79_groupi_g37132(csa_tree_add_51_79_groupi_n_8941 ,csa_tree_add_51_79_groupi_n_8445 ,csa_tree_add_51_79_groupi_n_8410);
  nor csa_tree_add_51_79_groupi_g37133(csa_tree_add_51_79_groupi_n_8940 ,csa_tree_add_51_79_groupi_n_7824 ,csa_tree_add_51_79_groupi_n_8409);
  and csa_tree_add_51_79_groupi_g37134(csa_tree_add_51_79_groupi_n_8939 ,csa_tree_add_51_79_groupi_n_8445 ,csa_tree_add_51_79_groupi_n_8410);
  or csa_tree_add_51_79_groupi_g37135(csa_tree_add_51_79_groupi_n_8938 ,csa_tree_add_51_79_groupi_n_8593 ,csa_tree_add_51_79_groupi_n_8407);
  and csa_tree_add_51_79_groupi_g37136(csa_tree_add_51_79_groupi_n_8937 ,csa_tree_add_51_79_groupi_n_8593 ,csa_tree_add_51_79_groupi_n_8407);
  or csa_tree_add_51_79_groupi_g37137(csa_tree_add_51_79_groupi_n_8936 ,csa_tree_add_51_79_groupi_n_8016 ,csa_tree_add_51_79_groupi_n_8449);
  and csa_tree_add_51_79_groupi_g37138(csa_tree_add_51_79_groupi_n_8935 ,csa_tree_add_51_79_groupi_n_8016 ,csa_tree_add_51_79_groupi_n_8449);
  and csa_tree_add_51_79_groupi_g37139(csa_tree_add_51_79_groupi_n_8934 ,csa_tree_add_51_79_groupi_n_8291 ,csa_tree_add_51_79_groupi_n_8388);
  or csa_tree_add_51_79_groupi_g37140(csa_tree_add_51_79_groupi_n_8933 ,csa_tree_add_51_79_groupi_n_8595 ,csa_tree_add_51_79_groupi_n_8406);
  or csa_tree_add_51_79_groupi_g37141(csa_tree_add_51_79_groupi_n_8932 ,csa_tree_add_51_79_groupi_n_8325 ,csa_tree_add_51_79_groupi_n_8539);
  or csa_tree_add_51_79_groupi_g37142(csa_tree_add_51_79_groupi_n_8931 ,csa_tree_add_51_79_groupi_n_8327 ,csa_tree_add_51_79_groupi_n_8537);
  nor csa_tree_add_51_79_groupi_g37143(csa_tree_add_51_79_groupi_n_8930 ,csa_tree_add_51_79_groupi_n_8599 ,csa_tree_add_51_79_groupi_n_8609);
  nor csa_tree_add_51_79_groupi_g37144(csa_tree_add_51_79_groupi_n_8929 ,csa_tree_add_51_79_groupi_n_8596 ,csa_tree_add_51_79_groupi_n_8405);
  or csa_tree_add_51_79_groupi_g37145(csa_tree_add_51_79_groupi_n_8928 ,csa_tree_add_51_79_groupi_n_8601 ,csa_tree_add_51_79_groupi_n_8610);
  and csa_tree_add_51_79_groupi_g37146(csa_tree_add_51_79_groupi_n_8927 ,csa_tree_add_51_79_groupi_n_8601 ,csa_tree_add_51_79_groupi_n_8610);
  or csa_tree_add_51_79_groupi_g37147(csa_tree_add_51_79_groupi_n_8926 ,csa_tree_add_51_79_groupi_n_8404 ,csa_tree_add_51_79_groupi_n_8425);
  and csa_tree_add_51_79_groupi_g37148(csa_tree_add_51_79_groupi_n_8925 ,csa_tree_add_51_79_groupi_n_8404 ,csa_tree_add_51_79_groupi_n_8425);
  or csa_tree_add_51_79_groupi_g37149(csa_tree_add_51_79_groupi_n_8924 ,csa_tree_add_51_79_groupi_n_8270 ,csa_tree_add_51_79_groupi_n_8443);
  nor csa_tree_add_51_79_groupi_g37150(csa_tree_add_51_79_groupi_n_8923 ,csa_tree_add_51_79_groupi_n_8401 ,csa_tree_add_51_79_groupi_n_8471);
  or csa_tree_add_51_79_groupi_g37151(csa_tree_add_51_79_groupi_n_8922 ,csa_tree_add_51_79_groupi_n_8600 ,csa_tree_add_51_79_groupi_n_8608);
  and csa_tree_add_51_79_groupi_g37152(csa_tree_add_51_79_groupi_n_8921 ,csa_tree_add_51_79_groupi_n_8615 ,csa_tree_add_51_79_groupi_n_8465);
  and csa_tree_add_51_79_groupi_g37153(csa_tree_add_51_79_groupi_n_8920 ,csa_tree_add_51_79_groupi_n_8401 ,csa_tree_add_51_79_groupi_n_8471);
  and csa_tree_add_51_79_groupi_g37154(csa_tree_add_51_79_groupi_n_8919 ,csa_tree_add_51_79_groupi_n_8270 ,csa_tree_add_51_79_groupi_n_8443);
  or csa_tree_add_51_79_groupi_g37155(csa_tree_add_51_79_groupi_n_8918 ,csa_tree_add_51_79_groupi_n_7823 ,csa_tree_add_51_79_groupi_n_8408);
  nor csa_tree_add_51_79_groupi_g37156(csa_tree_add_51_79_groupi_n_8917 ,csa_tree_add_51_79_groupi_n_8615 ,csa_tree_add_51_79_groupi_n_8465);
  and csa_tree_add_51_79_groupi_g37157(csa_tree_add_51_79_groupi_n_8916 ,csa_tree_add_51_79_groupi_n_8330 ,csa_tree_add_51_79_groupi_n_8528);
  or csa_tree_add_51_79_groupi_g37158(csa_tree_add_51_79_groupi_n_8915 ,csa_tree_add_51_79_groupi_n_8331 ,csa_tree_add_51_79_groupi_n_8549);
  or csa_tree_add_51_79_groupi_g37159(csa_tree_add_51_79_groupi_n_8914 ,csa_tree_add_51_79_groupi_n_8339 ,csa_tree_add_51_79_groupi_n_8565);
  or csa_tree_add_51_79_groupi_g37160(csa_tree_add_51_79_groupi_n_8913 ,csa_tree_add_51_79_groupi_n_8332 ,csa_tree_add_51_79_groupi_n_8518);
  or csa_tree_add_51_79_groupi_g37161(csa_tree_add_51_79_groupi_n_8912 ,csa_tree_add_51_79_groupi_n_8333 ,csa_tree_add_51_79_groupi_n_8512);
  or csa_tree_add_51_79_groupi_g37162(csa_tree_add_51_79_groupi_n_8911 ,csa_tree_add_51_79_groupi_n_8399 ,csa_tree_add_51_79_groupi_n_8424);
  and csa_tree_add_51_79_groupi_g37163(csa_tree_add_51_79_groupi_n_8910 ,csa_tree_add_51_79_groupi_n_8399 ,csa_tree_add_51_79_groupi_n_8424);
  and csa_tree_add_51_79_groupi_g37164(csa_tree_add_51_79_groupi_n_8909 ,csa_tree_add_51_79_groupi_n_8429 ,csa_tree_add_51_79_groupi_n_8428);
  or csa_tree_add_51_79_groupi_g37165(csa_tree_add_51_79_groupi_n_8908 ,csa_tree_add_51_79_groupi_n_8303 ,csa_tree_add_51_79_groupi_n_8398);
  nor csa_tree_add_51_79_groupi_g37166(csa_tree_add_51_79_groupi_n_8907 ,csa_tree_add_51_79_groupi_n_8304 ,csa_tree_add_51_79_groupi_n_8397);
  or csa_tree_add_51_79_groupi_g37167(csa_tree_add_51_79_groupi_n_8906 ,csa_tree_add_51_79_groupi_n_8463 ,csa_tree_add_51_79_groupi_n_8396);
  nor csa_tree_add_51_79_groupi_g37168(csa_tree_add_51_79_groupi_n_8905 ,csa_tree_add_51_79_groupi_n_8464 ,csa_tree_add_51_79_groupi_n_8395);
  or csa_tree_add_51_79_groupi_g37169(csa_tree_add_51_79_groupi_n_8904 ,csa_tree_add_51_79_groupi_n_8580 ,csa_tree_add_51_79_groupi_n_8575);
  or csa_tree_add_51_79_groupi_g37170(csa_tree_add_51_79_groupi_n_8903 ,csa_tree_add_51_79_groupi_n_8441 ,csa_tree_add_51_79_groupi_n_8394);
  and csa_tree_add_51_79_groupi_g37171(csa_tree_add_51_79_groupi_n_8902 ,csa_tree_add_51_79_groupi_n_8441 ,csa_tree_add_51_79_groupi_n_8394);
  nor csa_tree_add_51_79_groupi_g37172(csa_tree_add_51_79_groupi_n_8901 ,csa_tree_add_51_79_groupi_n_8581 ,csa_tree_add_51_79_groupi_n_8576);
  or csa_tree_add_51_79_groupi_g37173(csa_tree_add_51_79_groupi_n_8900 ,csa_tree_add_51_79_groupi_n_8181 ,csa_tree_add_51_79_groupi_n_8510);
  or csa_tree_add_51_79_groupi_g37174(csa_tree_add_51_79_groupi_n_8899 ,csa_tree_add_51_79_groupi_n_8440 ,csa_tree_add_51_79_groupi_n_8393);
  and csa_tree_add_51_79_groupi_g37175(csa_tree_add_51_79_groupi_n_8898 ,csa_tree_add_51_79_groupi_n_8440 ,csa_tree_add_51_79_groupi_n_8393);
  or csa_tree_add_51_79_groupi_g37176(csa_tree_add_51_79_groupi_n_8897 ,csa_tree_add_51_79_groupi_n_8392 ,csa_tree_add_51_79_groupi_n_8439);
  and csa_tree_add_51_79_groupi_g37177(csa_tree_add_51_79_groupi_n_8896 ,csa_tree_add_51_79_groupi_n_8392 ,csa_tree_add_51_79_groupi_n_8439);
  or csa_tree_add_51_79_groupi_g37178(csa_tree_add_51_79_groupi_n_8895 ,csa_tree_add_51_79_groupi_n_8429 ,csa_tree_add_51_79_groupi_n_8428);
  or csa_tree_add_51_79_groupi_g37179(csa_tree_add_51_79_groupi_n_8894 ,csa_tree_add_51_79_groupi_n_8305 ,csa_tree_add_51_79_groupi_n_8473);
  and csa_tree_add_51_79_groupi_g37180(csa_tree_add_51_79_groupi_n_8893 ,csa_tree_add_51_79_groupi_n_8305 ,csa_tree_add_51_79_groupi_n_8473);
  or csa_tree_add_51_79_groupi_g37181(csa_tree_add_51_79_groupi_n_8892 ,csa_tree_add_51_79_groupi_n_8342 ,csa_tree_add_51_79_groupi_n_8511);
  or csa_tree_add_51_79_groupi_g37182(csa_tree_add_51_79_groupi_n_8891 ,csa_tree_add_51_79_groupi_n_8338 ,csa_tree_add_51_79_groupi_n_8365);
  or csa_tree_add_51_79_groupi_g37183(csa_tree_add_51_79_groupi_n_8890 ,csa_tree_add_51_79_groupi_n_8337 ,csa_tree_add_51_79_groupi_n_8514);
  or csa_tree_add_51_79_groupi_g37184(csa_tree_add_51_79_groupi_n_8889 ,csa_tree_add_51_79_groupi_n_8458 ,csa_tree_add_51_79_groupi_n_8391);
  nor csa_tree_add_51_79_groupi_g37185(csa_tree_add_51_79_groupi_n_8888 ,csa_tree_add_51_79_groupi_n_8578 ,csa_tree_add_51_79_groupi_n_8583);
  nor csa_tree_add_51_79_groupi_g37186(csa_tree_add_51_79_groupi_n_8887 ,csa_tree_add_51_79_groupi_n_8459 ,csa_tree_add_51_79_groupi_n_8390);
  and csa_tree_add_51_79_groupi_g37187(csa_tree_add_51_79_groupi_n_8886 ,csa_tree_add_51_79_groupi_n_8343 ,csa_tree_add_51_79_groupi_n_8513);
  nor csa_tree_add_51_79_groupi_g37188(csa_tree_add_51_79_groupi_n_8885 ,csa_tree_add_51_79_groupi_n_8370 ,csa_tree_add_51_79_groupi_n_8588);
  or csa_tree_add_51_79_groupi_g37189(csa_tree_add_51_79_groupi_n_8884 ,csa_tree_add_51_79_groupi_n_8577 ,csa_tree_add_51_79_groupi_n_8584);
  or csa_tree_add_51_79_groupi_g37190(csa_tree_add_51_79_groupi_n_8883 ,csa_tree_add_51_79_groupi_n_8389 ,csa_tree_add_51_79_groupi_n_8387);
  and csa_tree_add_51_79_groupi_g37191(csa_tree_add_51_79_groupi_n_8882 ,csa_tree_add_51_79_groupi_n_8389 ,csa_tree_add_51_79_groupi_n_8387);
  or csa_tree_add_51_79_groupi_g37192(csa_tree_add_51_79_groupi_n_8881 ,csa_tree_add_51_79_groupi_n_8466 ,csa_tree_add_51_79_groupi_n_8386);
  or csa_tree_add_51_79_groupi_g37193(csa_tree_add_51_79_groupi_n_8880 ,csa_tree_add_51_79_groupi_n_8436 ,csa_tree_add_51_79_groupi_n_8384);
  nor csa_tree_add_51_79_groupi_g37194(csa_tree_add_51_79_groupi_n_8879 ,csa_tree_add_51_79_groupi_n_8467 ,csa_tree_add_51_79_groupi_n_8385);
  or csa_tree_add_51_79_groupi_g37195(csa_tree_add_51_79_groupi_n_8878 ,csa_tree_add_51_79_groupi_n_8377 ,csa_tree_add_51_79_groupi_n_8416);
  and csa_tree_add_51_79_groupi_g37196(csa_tree_add_51_79_groupi_n_8877 ,csa_tree_add_51_79_groupi_n_8436 ,csa_tree_add_51_79_groupi_n_8384);
  nor csa_tree_add_51_79_groupi_g37197(csa_tree_add_51_79_groupi_n_8876 ,csa_tree_add_51_79_groupi_n_8376 ,csa_tree_add_51_79_groupi_n_8417);
  and csa_tree_add_51_79_groupi_g37198(csa_tree_add_51_79_groupi_n_8875 ,csa_tree_add_51_79_groupi_n_8607 ,csa_tree_add_51_79_groupi_n_8604);
  or csa_tree_add_51_79_groupi_g37199(csa_tree_add_51_79_groupi_n_8874 ,csa_tree_add_51_79_groupi_n_8597 ,csa_tree_add_51_79_groupi_n_8383);
  nor csa_tree_add_51_79_groupi_g37200(csa_tree_add_51_79_groupi_n_8873 ,csa_tree_add_51_79_groupi_n_8446 ,csa_tree_add_51_79_groupi_n_8442);
  or csa_tree_add_51_79_groupi_g37201(csa_tree_add_51_79_groupi_n_8872 ,csa_tree_add_51_79_groupi_n_8460 ,csa_tree_add_51_79_groupi_n_8381);
  and csa_tree_add_51_79_groupi_g37202(csa_tree_add_51_79_groupi_n_8871 ,csa_tree_add_51_79_groupi_n_8460 ,csa_tree_add_51_79_groupi_n_8381);
  or csa_tree_add_51_79_groupi_g37203(csa_tree_add_51_79_groupi_n_8870 ,csa_tree_add_51_79_groupi_n_8613 ,csa_tree_add_51_79_groupi_n_8476);
  nor csa_tree_add_51_79_groupi_g37204(csa_tree_add_51_79_groupi_n_8869 ,csa_tree_add_51_79_groupi_n_8612 ,csa_tree_add_51_79_groupi_n_8477);
  nor csa_tree_add_51_79_groupi_g37205(csa_tree_add_51_79_groupi_n_8868 ,csa_tree_add_51_79_groupi_n_8598 ,csa_tree_add_51_79_groupi_n_8382);
  or csa_tree_add_51_79_groupi_g37206(csa_tree_add_51_79_groupi_n_8867 ,csa_tree_add_51_79_groupi_n_8326 ,csa_tree_add_51_79_groupi_n_8523);
  or csa_tree_add_51_79_groupi_g37207(csa_tree_add_51_79_groupi_n_8866 ,csa_tree_add_51_79_groupi_n_8607 ,csa_tree_add_51_79_groupi_n_8604);
  or csa_tree_add_51_79_groupi_g37208(csa_tree_add_51_79_groupi_n_8865 ,csa_tree_add_51_79_groupi_n_8485 ,csa_tree_add_51_79_groupi_n_8527);
  or csa_tree_add_51_79_groupi_g37209(csa_tree_add_51_79_groupi_n_8864 ,csa_tree_add_51_79_groupi_n_8493 ,csa_tree_add_51_79_groupi_n_8236);
  and csa_tree_add_51_79_groupi_g37210(csa_tree_add_51_79_groupi_n_8863 ,csa_tree_add_51_79_groupi_n_8430 ,csa_tree_add_51_79_groupi_n_8400);
  or csa_tree_add_51_79_groupi_g37211(csa_tree_add_51_79_groupi_n_8862 ,csa_tree_add_51_79_groupi_n_8402 ,csa_tree_add_51_79_groupi_n_8569);
  or csa_tree_add_51_79_groupi_g37212(csa_tree_add_51_79_groupi_n_8861 ,csa_tree_add_51_79_groupi_n_8430 ,csa_tree_add_51_79_groupi_n_8400);
  nor csa_tree_add_51_79_groupi_g37213(csa_tree_add_51_79_groupi_n_8860 ,csa_tree_add_51_79_groupi_n_8403 ,csa_tree_add_51_79_groupi_n_8568);
  and csa_tree_add_51_79_groupi_g37214(csa_tree_add_51_79_groupi_n_8859 ,csa_tree_add_51_79_groupi_n_8434 ,csa_tree_add_51_79_groupi_n_8421);
  or csa_tree_add_51_79_groupi_g37215(csa_tree_add_51_79_groupi_n_8858 ,csa_tree_add_51_79_groupi_n_8317 ,csa_tree_add_51_79_groupi_n_8535);
  or csa_tree_add_51_79_groupi_g37216(csa_tree_add_51_79_groupi_n_8857 ,csa_tree_add_51_79_groupi_n_8316 ,csa_tree_add_51_79_groupi_n_8536);
  or csa_tree_add_51_79_groupi_g37217(csa_tree_add_51_79_groupi_n_8856 ,csa_tree_add_51_79_groupi_n_8437 ,csa_tree_add_51_79_groupi_n_8375);
  nor csa_tree_add_51_79_groupi_g37218(csa_tree_add_51_79_groupi_n_8855 ,csa_tree_add_51_79_groupi_n_8438 ,csa_tree_add_51_79_groupi_n_8374);
  or csa_tree_add_51_79_groupi_g37219(csa_tree_add_51_79_groupi_n_8854 ,csa_tree_add_51_79_groupi_n_8314 ,csa_tree_add_51_79_groupi_n_8541);
  or csa_tree_add_51_79_groupi_g37220(csa_tree_add_51_79_groupi_n_8853 ,csa_tree_add_51_79_groupi_n_7830 ,csa_tree_add_51_79_groupi_n_8543);
  or csa_tree_add_51_79_groupi_g37221(csa_tree_add_51_79_groupi_n_8852 ,csa_tree_add_51_79_groupi_n_8269 ,csa_tree_add_51_79_groupi_n_8373);
  or csa_tree_add_51_79_groupi_g37222(csa_tree_add_51_79_groupi_n_8851 ,csa_tree_add_51_79_groupi_n_8450 ,csa_tree_add_51_79_groupi_n_8622);
  and csa_tree_add_51_79_groupi_g37223(csa_tree_add_51_79_groupi_n_8850 ,csa_tree_add_51_79_groupi_n_8269 ,csa_tree_add_51_79_groupi_n_8373);
  or csa_tree_add_51_79_groupi_g37224(csa_tree_add_51_79_groupi_n_8849 ,csa_tree_add_51_79_groupi_n_8590 ,csa_tree_add_51_79_groupi_n_8372);
  nor csa_tree_add_51_79_groupi_g37225(csa_tree_add_51_79_groupi_n_8848 ,csa_tree_add_51_79_groupi_n_8451 ,csa_tree_add_51_79_groupi_n_8621);
  and csa_tree_add_51_79_groupi_g37226(csa_tree_add_51_79_groupi_n_8847 ,csa_tree_add_51_79_groupi_n_8590 ,csa_tree_add_51_79_groupi_n_8372);
  or csa_tree_add_51_79_groupi_g37227(csa_tree_add_51_79_groupi_n_8846 ,csa_tree_add_51_79_groupi_n_8371 ,csa_tree_add_51_79_groupi_n_8587);
  or csa_tree_add_51_79_groupi_g37228(csa_tree_add_51_79_groupi_n_8845 ,csa_tree_add_51_79_groupi_n_8419 ,csa_tree_add_51_79_groupi_n_8433);
  nor csa_tree_add_51_79_groupi_g37229(csa_tree_add_51_79_groupi_n_8844 ,csa_tree_add_51_79_groupi_n_8420 ,csa_tree_add_51_79_groupi_n_8432);
  or csa_tree_add_51_79_groupi_g37230(csa_tree_add_51_79_groupi_n_8843 ,csa_tree_add_51_79_groupi_n_8434 ,csa_tree_add_51_79_groupi_n_8421);
  or csa_tree_add_51_79_groupi_g37231(csa_tree_add_51_79_groupi_n_8842 ,csa_tree_add_51_79_groupi_n_8157 ,csa_tree_add_51_79_groupi_n_8474);
  and csa_tree_add_51_79_groupi_g37232(csa_tree_add_51_79_groupi_n_8841 ,csa_tree_add_51_79_groupi_n_8157 ,csa_tree_add_51_79_groupi_n_8474);
  or csa_tree_add_51_79_groupi_g37233(csa_tree_add_51_79_groupi_n_8840 ,csa_tree_add_51_79_groupi_n_8155 ,csa_tree_add_51_79_groupi_n_8431);
  and csa_tree_add_51_79_groupi_g37234(csa_tree_add_51_79_groupi_n_8839 ,csa_tree_add_51_79_groupi_n_8155 ,csa_tree_add_51_79_groupi_n_8431);
  or csa_tree_add_51_79_groupi_g37235(csa_tree_add_51_79_groupi_n_8838 ,csa_tree_add_51_79_groupi_n_8182 ,csa_tree_add_51_79_groupi_n_8551);
  or csa_tree_add_51_79_groupi_g37236(csa_tree_add_51_79_groupi_n_8837 ,csa_tree_add_51_79_groupi_n_8180 ,csa_tree_add_51_79_groupi_n_8559);
  or csa_tree_add_51_79_groupi_g37237(csa_tree_add_51_79_groupi_n_8836 ,csa_tree_add_51_79_groupi_n_8444 ,csa_tree_add_51_79_groupi_n_8427);
  and csa_tree_add_51_79_groupi_g37238(csa_tree_add_51_79_groupi_n_8835 ,csa_tree_add_51_79_groupi_n_8444 ,csa_tree_add_51_79_groupi_n_8427);
  or csa_tree_add_51_79_groupi_g37239(csa_tree_add_51_79_groupi_n_8834 ,csa_tree_add_51_79_groupi_n_8426 ,csa_tree_add_51_79_groupi_n_8579);
  and csa_tree_add_51_79_groupi_g37240(csa_tree_add_51_79_groupi_n_8833 ,csa_tree_add_51_79_groupi_n_8426 ,csa_tree_add_51_79_groupi_n_8579);
  or csa_tree_add_51_79_groupi_g37241(csa_tree_add_51_79_groupi_n_8832 ,csa_tree_add_51_79_groupi_n_8378 ,csa_tree_add_51_79_groupi_n_8611);
  and csa_tree_add_51_79_groupi_g37242(csa_tree_add_51_79_groupi_n_8831 ,csa_tree_add_51_79_groupi_n_8378 ,csa_tree_add_51_79_groupi_n_8611);
  or csa_tree_add_51_79_groupi_g37243(csa_tree_add_51_79_groupi_n_8830 ,csa_tree_add_51_79_groupi_n_8475 ,csa_tree_add_51_79_groupi_n_8567);
  and csa_tree_add_51_79_groupi_g37244(csa_tree_add_51_79_groupi_n_8829 ,csa_tree_add_51_79_groupi_n_8475 ,csa_tree_add_51_79_groupi_n_8567);
  or csa_tree_add_51_79_groupi_g37245(csa_tree_add_51_79_groupi_n_8828 ,csa_tree_add_51_79_groupi_n_8453 ,csa_tree_add_51_79_groupi_n_8435);
  and csa_tree_add_51_79_groupi_g37246(csa_tree_add_51_79_groupi_n_8827 ,csa_tree_add_51_79_groupi_n_8453 ,csa_tree_add_51_79_groupi_n_8435);
  or csa_tree_add_51_79_groupi_g37247(csa_tree_add_51_79_groupi_n_8826 ,csa_tree_add_51_79_groupi_n_8582 ,csa_tree_add_51_79_groupi_n_8422);
  and csa_tree_add_51_79_groupi_g37248(csa_tree_add_51_79_groupi_n_8825 ,csa_tree_add_51_79_groupi_n_8582 ,csa_tree_add_51_79_groupi_n_8422);
  and csa_tree_add_51_79_groupi_g37249(csa_tree_add_51_79_groupi_n_8970 ,csa_tree_add_51_79_groupi_n_7902 ,csa_tree_add_51_79_groupi_n_8566);
  and csa_tree_add_51_79_groupi_g37250(csa_tree_add_51_79_groupi_n_8969 ,csa_tree_add_51_79_groupi_n_8122 ,csa_tree_add_51_79_groupi_n_8544);
  and csa_tree_add_51_79_groupi_g37251(csa_tree_add_51_79_groupi_n_8968 ,csa_tree_add_51_79_groupi_n_7845 ,csa_tree_add_51_79_groupi_n_8529);
  and csa_tree_add_51_79_groupi_g37252(csa_tree_add_51_79_groupi_n_8967 ,csa_tree_add_51_79_groupi_n_8240 ,csa_tree_add_51_79_groupi_n_8545);
  and csa_tree_add_51_79_groupi_g37253(csa_tree_add_51_79_groupi_n_8966 ,csa_tree_add_51_79_groupi_n_8234 ,csa_tree_add_51_79_groupi_n_8526);
  or csa_tree_add_51_79_groupi_g37254(csa_tree_add_51_79_groupi_n_8965 ,csa_tree_add_51_79_groupi_n_8210 ,csa_tree_add_51_79_groupi_n_8525);
  and csa_tree_add_51_79_groupi_g37255(csa_tree_add_51_79_groupi_n_8964 ,csa_tree_add_51_79_groupi_n_8141 ,csa_tree_add_51_79_groupi_n_8547);
  and csa_tree_add_51_79_groupi_g37256(csa_tree_add_51_79_groupi_n_8963 ,csa_tree_add_51_79_groupi_n_8255 ,csa_tree_add_51_79_groupi_n_8556);
  and csa_tree_add_51_79_groupi_g37257(csa_tree_add_51_79_groupi_n_8961 ,csa_tree_add_51_79_groupi_n_8012 ,csa_tree_add_51_79_groupi_n_8564);
  and csa_tree_add_51_79_groupi_g37258(csa_tree_add_51_79_groupi_n_8960 ,csa_tree_add_51_79_groupi_n_8254 ,csa_tree_add_51_79_groupi_n_8532);
  and csa_tree_add_51_79_groupi_g37259(csa_tree_add_51_79_groupi_n_8959 ,csa_tree_add_51_79_groupi_n_8202 ,csa_tree_add_51_79_groupi_n_8517);
  and csa_tree_add_51_79_groupi_g37260(csa_tree_add_51_79_groupi_n_8958 ,csa_tree_add_51_79_groupi_n_8145 ,csa_tree_add_51_79_groupi_n_8531);
  not csa_tree_add_51_79_groupi_g37261(csa_tree_add_51_79_groupi_n_8797 ,csa_tree_add_51_79_groupi_n_8796);
  not csa_tree_add_51_79_groupi_g37262(csa_tree_add_51_79_groupi_n_8793 ,csa_tree_add_51_79_groupi_n_8792);
  not csa_tree_add_51_79_groupi_g37263(csa_tree_add_51_79_groupi_n_8789 ,csa_tree_add_51_79_groupi_n_8790);
  not csa_tree_add_51_79_groupi_g37264(csa_tree_add_51_79_groupi_n_8787 ,csa_tree_add_51_79_groupi_n_8788);
  not csa_tree_add_51_79_groupi_g37265(csa_tree_add_51_79_groupi_n_8783 ,csa_tree_add_51_79_groupi_n_8784);
  not csa_tree_add_51_79_groupi_g37266(csa_tree_add_51_79_groupi_n_8781 ,csa_tree_add_51_79_groupi_n_8782);
  not csa_tree_add_51_79_groupi_g37267(csa_tree_add_51_79_groupi_n_8776 ,csa_tree_add_51_79_groupi_n_8777);
  not csa_tree_add_51_79_groupi_g37268(csa_tree_add_51_79_groupi_n_8773 ,csa_tree_add_51_79_groupi_n_8774);
  not csa_tree_add_51_79_groupi_g37269(csa_tree_add_51_79_groupi_n_8768 ,csa_tree_add_51_79_groupi_n_8767);
  not csa_tree_add_51_79_groupi_g37270(csa_tree_add_51_79_groupi_n_8762 ,csa_tree_add_51_79_groupi_n_8763);
  not csa_tree_add_51_79_groupi_g37271(csa_tree_add_51_79_groupi_n_8757 ,csa_tree_add_51_79_groupi_n_8758);
  not csa_tree_add_51_79_groupi_g37272(csa_tree_add_51_79_groupi_n_8753 ,csa_tree_add_51_79_groupi_n_8754);
  not csa_tree_add_51_79_groupi_g37273(csa_tree_add_51_79_groupi_n_8751 ,csa_tree_add_51_79_groupi_n_8752);
  not csa_tree_add_51_79_groupi_g37274(csa_tree_add_51_79_groupi_n_8748 ,csa_tree_add_51_79_groupi_n_8749);
  not csa_tree_add_51_79_groupi_g37275(csa_tree_add_51_79_groupi_n_8745 ,csa_tree_add_51_79_groupi_n_8746);
  not csa_tree_add_51_79_groupi_g37276(csa_tree_add_51_79_groupi_n_8739 ,csa_tree_add_51_79_groupi_n_8740);
  not csa_tree_add_51_79_groupi_g37277(csa_tree_add_51_79_groupi_n_8731 ,csa_tree_add_51_79_groupi_n_8732);
  not csa_tree_add_51_79_groupi_g37278(csa_tree_add_51_79_groupi_n_8727 ,csa_tree_add_51_79_groupi_n_8728);
  not csa_tree_add_51_79_groupi_g37279(csa_tree_add_51_79_groupi_n_8724 ,csa_tree_add_51_79_groupi_n_8725);
  not csa_tree_add_51_79_groupi_g37280(csa_tree_add_51_79_groupi_n_8718 ,csa_tree_add_51_79_groupi_n_8719);
  or csa_tree_add_51_79_groupi_g37281(csa_tree_add_51_79_groupi_n_8716 ,csa_tree_add_51_79_groupi_n_8183 ,csa_tree_add_51_79_groupi_n_8367);
  or csa_tree_add_51_79_groupi_g37282(csa_tree_add_51_79_groupi_n_8715 ,csa_tree_add_51_79_groupi_n_7370 ,csa_tree_add_51_79_groupi_n_8363);
  or csa_tree_add_51_79_groupi_g37283(csa_tree_add_51_79_groupi_n_8714 ,csa_tree_add_51_79_groupi_n_8176 ,csa_tree_add_51_79_groupi_n_8415);
  and csa_tree_add_51_79_groupi_g37284(csa_tree_add_51_79_groupi_n_8713 ,csa_tree_add_51_79_groupi_n_8176 ,csa_tree_add_51_79_groupi_n_8415);
  or csa_tree_add_51_79_groupi_g37285(csa_tree_add_51_79_groupi_n_8712 ,csa_tree_add_51_79_groupi_n_7806 ,csa_tree_add_51_79_groupi_n_8461);
  and csa_tree_add_51_79_groupi_g37286(csa_tree_add_51_79_groupi_n_8711 ,csa_tree_add_51_79_groupi_n_7806 ,csa_tree_add_51_79_groupi_n_8461);
  or csa_tree_add_51_79_groupi_g37287(csa_tree_add_51_79_groupi_n_8710 ,csa_tree_add_51_79_groupi_n_8020 ,csa_tree_add_51_79_groupi_n_8472);
  and csa_tree_add_51_79_groupi_g37288(csa_tree_add_51_79_groupi_n_8709 ,csa_tree_add_51_79_groupi_n_8020 ,csa_tree_add_51_79_groupi_n_8472);
  or csa_tree_add_51_79_groupi_g37289(csa_tree_add_51_79_groupi_n_8708 ,csa_tree_add_51_79_groupi_n_8286 ,csa_tree_add_51_79_groupi_n_8462);
  and csa_tree_add_51_79_groupi_g37290(csa_tree_add_51_79_groupi_n_8707 ,csa_tree_add_51_79_groupi_n_8286 ,csa_tree_add_51_79_groupi_n_8462);
  or csa_tree_add_51_79_groupi_g37291(csa_tree_add_51_79_groupi_n_8706 ,csa_tree_add_51_79_groupi_n_7356 ,csa_tree_add_51_79_groupi_n_8361);
  or csa_tree_add_51_79_groupi_g37292(csa_tree_add_51_79_groupi_n_8705 ,csa_tree_add_51_79_groupi_n_8165 ,csa_tree_add_51_79_groupi_n_8413);
  or csa_tree_add_51_79_groupi_g37293(csa_tree_add_51_79_groupi_n_8704 ,csa_tree_add_51_79_groupi_n_8592 ,csa_tree_add_51_79_groupi_n_8478);
  nor csa_tree_add_51_79_groupi_g37294(csa_tree_add_51_79_groupi_n_8703 ,csa_tree_add_51_79_groupi_n_8457 ,csa_tree_add_51_79_groupi_n_8455);
  or csa_tree_add_51_79_groupi_g37295(csa_tree_add_51_79_groupi_n_8702 ,csa_tree_add_51_79_groupi_n_8619 ,csa_tree_add_51_79_groupi_n_8617);
  nor csa_tree_add_51_79_groupi_g37296(csa_tree_add_51_79_groupi_n_8701 ,csa_tree_add_51_79_groupi_n_8164 ,csa_tree_add_51_79_groupi_n_8414);
  nor csa_tree_add_51_79_groupi_g37297(csa_tree_add_51_79_groupi_n_8700 ,csa_tree_add_51_79_groupi_n_8620 ,csa_tree_add_51_79_groupi_n_8618);
  nor csa_tree_add_51_79_groupi_g37298(csa_tree_add_51_79_groupi_n_8699 ,csa_tree_add_51_79_groupi_n_8591 ,csa_tree_add_51_79_groupi_n_8479);
  and csa_tree_add_51_79_groupi_g37299(csa_tree_add_51_79_groupi_n_8698 ,csa_tree_add_51_79_groupi_n_8315 ,csa_tree_add_51_79_groupi_n_8359);
  or csa_tree_add_51_79_groupi_g37300(csa_tree_add_51_79_groupi_n_8697 ,csa_tree_add_51_79_groupi_n_8158 ,csa_tree_add_51_79_groupi_n_8379);
  or csa_tree_add_51_79_groupi_g37301(csa_tree_add_51_79_groupi_n_8696 ,csa_tree_add_51_79_groupi_n_8483 ,csa_tree_add_51_79_groupi_n_8481);
  nor csa_tree_add_51_79_groupi_g37302(csa_tree_add_51_79_groupi_n_8695 ,csa_tree_add_51_79_groupi_n_8159 ,csa_tree_add_51_79_groupi_n_8380);
  nor csa_tree_add_51_79_groupi_g37303(csa_tree_add_51_79_groupi_n_8694 ,csa_tree_add_51_79_groupi_n_8484 ,csa_tree_add_51_79_groupi_n_8482);
  or csa_tree_add_51_79_groupi_g37304(csa_tree_add_51_79_groupi_n_8693 ,csa_tree_add_51_79_groupi_n_8585 ,csa_tree_add_51_79_groupi_n_8468);
  nor csa_tree_add_51_79_groupi_g37305(csa_tree_add_51_79_groupi_n_8692 ,csa_tree_add_51_79_groupi_n_8586 ,csa_tree_add_51_79_groupi_n_8469);
  or csa_tree_add_51_79_groupi_g37306(csa_tree_add_51_79_groupi_n_8691 ,csa_tree_add_51_79_groupi_n_8456 ,csa_tree_add_51_79_groupi_n_8454);
  xnor csa_tree_add_51_79_groupi_g37307(csa_tree_add_51_79_groupi_n_8690 ,csa_tree_add_51_79_groupi_n_8183 ,csa_tree_add_51_79_groupi_n_8168);
  xnor csa_tree_add_51_79_groupi_g37308(csa_tree_add_51_79_groupi_n_8689 ,csa_tree_add_51_79_groupi_n_8298 ,csa_tree_add_51_79_groupi_n_8265);
  xnor csa_tree_add_51_79_groupi_g37309(csa_tree_add_51_79_groupi_n_8688 ,csa_tree_add_51_79_groupi_n_8295 ,csa_tree_add_51_79_groupi_n_7301);
  xnor csa_tree_add_51_79_groupi_g37310(csa_tree_add_51_79_groupi_n_8687 ,csa_tree_add_51_79_groupi_n_8019 ,csa_tree_add_51_79_groupi_n_8163);
  xnor csa_tree_add_51_79_groupi_g37311(csa_tree_add_51_79_groupi_n_8686 ,csa_tree_add_51_79_groupi_n_8153 ,csa_tree_add_51_79_groupi_n_8166);
  xnor csa_tree_add_51_79_groupi_g37312(csa_tree_add_51_79_groupi_n_8685 ,csa_tree_add_51_79_groupi_n_8180 ,csa_tree_add_51_79_groupi_n_8151);
  xnor csa_tree_add_51_79_groupi_g37313(csa_tree_add_51_79_groupi_n_8684 ,csa_tree_add_51_79_groupi_n_7824 ,csa_tree_add_51_79_groupi_n_8323);
  xnor csa_tree_add_51_79_groupi_g37314(csa_tree_add_51_79_groupi_n_8683 ,csa_tree_add_51_79_groupi_n_8302 ,csa_tree_add_51_79_groupi_n_8017);
  xnor csa_tree_add_51_79_groupi_g37315(csa_tree_add_51_79_groupi_n_8682 ,csa_tree_add_51_79_groupi_n_8170 ,csa_tree_add_51_79_groupi_n_7340);
  xnor csa_tree_add_51_79_groupi_g37316(csa_tree_add_51_79_groupi_n_8681 ,csa_tree_add_51_79_groupi_n_8177 ,csa_tree_add_51_79_groupi_n_8169);
  xnor csa_tree_add_51_79_groupi_g37317(csa_tree_add_51_79_groupi_n_8680 ,csa_tree_add_51_79_groupi_n_6855 ,csa_tree_add_51_79_groupi_n_8267);
  xnor csa_tree_add_51_79_groupi_g37318(csa_tree_add_51_79_groupi_n_8679 ,csa_tree_add_51_79_groupi_n_7607 ,csa_tree_add_51_79_groupi_n_8307);
  xnor csa_tree_add_51_79_groupi_g37319(csa_tree_add_51_79_groupi_n_8678 ,csa_tree_add_51_79_groupi_n_8167 ,csa_tree_add_51_79_groupi_n_7370);
  xnor csa_tree_add_51_79_groupi_g37320(csa_tree_add_51_79_groupi_n_8677 ,csa_tree_add_51_79_groupi_n_8283 ,csa_tree_add_51_79_groupi_n_8316);
  xnor csa_tree_add_51_79_groupi_g37321(csa_tree_add_51_79_groupi_n_8676 ,csa_tree_add_51_79_groupi_n_8292 ,csa_tree_add_51_79_groupi_n_8161);
  xnor csa_tree_add_51_79_groupi_g37322(csa_tree_add_51_79_groupi_n_8675 ,csa_tree_add_51_79_groupi_n_8276 ,csa_tree_add_51_79_groupi_n_8160);
  xnor csa_tree_add_51_79_groupi_g37323(csa_tree_add_51_79_groupi_n_8674 ,csa_tree_add_51_79_groupi_n_8282 ,csa_tree_add_51_79_groupi_n_8312);
  xnor csa_tree_add_51_79_groupi_g37324(csa_tree_add_51_79_groupi_n_8673 ,csa_tree_add_51_79_groupi_n_8278 ,csa_tree_add_51_79_groupi_n_7249);
  xnor csa_tree_add_51_79_groupi_g37325(csa_tree_add_51_79_groupi_n_8672 ,csa_tree_add_51_79_groupi_n_8273 ,csa_tree_add_51_79_groupi_n_7804);
  xnor csa_tree_add_51_79_groupi_g37326(csa_tree_add_51_79_groupi_n_8671 ,csa_tree_add_51_79_groupi_n_8319 ,csa_tree_add_51_79_groupi_n_7820);
  xnor csa_tree_add_51_79_groupi_g37327(csa_tree_add_51_79_groupi_n_8670 ,csa_tree_add_51_79_groupi_n_8296 ,csa_tree_add_51_79_groupi_n_8317);
  xnor csa_tree_add_51_79_groupi_g37328(csa_tree_add_51_79_groupi_n_8669 ,csa_tree_add_51_79_groupi_n_8279 ,csa_tree_add_51_79_groupi_n_8277);
  xnor csa_tree_add_51_79_groupi_g37329(csa_tree_add_51_79_groupi_n_8668 ,csa_tree_add_51_79_groupi_n_8325 ,csa_tree_add_51_79_groupi_n_8297);
  xnor csa_tree_add_51_79_groupi_g37330(csa_tree_add_51_79_groupi_n_8667 ,csa_tree_add_51_79_groupi_n_8290 ,csa_tree_add_51_79_groupi_n_8289);
  xnor csa_tree_add_51_79_groupi_g37331(csa_tree_add_51_79_groupi_n_8666 ,csa_tree_add_51_79_groupi_n_8308 ,csa_tree_add_51_79_groupi_n_8327);
  xnor csa_tree_add_51_79_groupi_g37332(csa_tree_add_51_79_groupi_n_8665 ,csa_tree_add_51_79_groupi_n_8321 ,csa_tree_add_51_79_groupi_n_8291);
  xnor csa_tree_add_51_79_groupi_g37333(csa_tree_add_51_79_groupi_n_8664 ,csa_tree_add_51_79_groupi_n_8287 ,csa_tree_add_51_79_groupi_n_8332);
  xnor csa_tree_add_51_79_groupi_g37334(csa_tree_add_51_79_groupi_n_8663 ,csa_tree_add_51_79_groupi_n_8299 ,csa_tree_add_51_79_groupi_n_8284);
  xnor csa_tree_add_51_79_groupi_g37335(csa_tree_add_51_79_groupi_n_8662 ,csa_tree_add_51_79_groupi_n_8305 ,csa_tree_add_51_79_groupi_n_8341);
  xnor csa_tree_add_51_79_groupi_g37336(csa_tree_add_51_79_groupi_n_8661 ,csa_tree_add_51_79_groupi_n_8333 ,csa_tree_add_51_79_groupi_n_8285);
  xnor csa_tree_add_51_79_groupi_g37337(csa_tree_add_51_79_groupi_n_8660 ,csa_tree_add_51_79_groupi_n_8311 ,csa_tree_add_51_79_groupi_n_8326);
  xnor csa_tree_add_51_79_groupi_g37338(csa_tree_add_51_79_groupi_n_8659 ,csa_tree_add_51_79_groupi_n_8301 ,csa_tree_add_51_79_groupi_n_8268);
  xnor csa_tree_add_51_79_groupi_g37339(csa_tree_add_51_79_groupi_n_8824 ,csa_tree_add_51_79_groupi_n_7363 ,csa_tree_add_51_79_groupi_n_8060);
  xnor csa_tree_add_51_79_groupi_g37340(csa_tree_add_51_79_groupi_n_8823 ,csa_tree_add_51_79_groupi_n_7827 ,csa_tree_add_51_79_groupi_n_8036);
  xnor csa_tree_add_51_79_groupi_g37341(csa_tree_add_51_79_groupi_n_8822 ,csa_tree_add_51_79_groupi_n_7368 ,csa_tree_add_51_79_groupi_n_8058);
  xnor csa_tree_add_51_79_groupi_g37342(csa_tree_add_51_79_groupi_n_8821 ,csa_tree_add_51_79_groupi_n_7241 ,csa_tree_add_51_79_groupi_n_8054);
  xnor csa_tree_add_51_79_groupi_g37343(csa_tree_add_51_79_groupi_n_8820 ,csa_tree_add_51_79_groupi_n_7295 ,csa_tree_add_51_79_groupi_n_8056);
  xnor csa_tree_add_51_79_groupi_g37344(csa_tree_add_51_79_groupi_n_8819 ,csa_tree_add_51_79_groupi_n_7175 ,csa_tree_add_51_79_groupi_n_8102);
  xnor csa_tree_add_51_79_groupi_g37345(csa_tree_add_51_79_groupi_n_8818 ,csa_tree_add_51_79_groupi_n_8156 ,csa_tree_add_51_79_groupi_n_8075);
  xnor csa_tree_add_51_79_groupi_g37346(csa_tree_add_51_79_groupi_n_8817 ,csa_tree_add_51_79_groupi_n_7324 ,csa_tree_add_51_79_groupi_n_8112);
  xnor csa_tree_add_51_79_groupi_g37347(csa_tree_add_51_79_groupi_n_8816 ,csa_tree_add_51_79_groupi_n_7600 ,csa_tree_add_51_79_groupi_n_8033);
  xnor csa_tree_add_51_79_groupi_g37348(csa_tree_add_51_79_groupi_n_8815 ,csa_tree_add_51_79_groupi_n_7374 ,csa_tree_add_51_79_groupi_n_8064);
  xor csa_tree_add_51_79_groupi_g37349(csa_tree_add_51_79_groupi_n_8814 ,csa_tree_add_51_79_groupi_n_6404 ,csa_tree_add_51_79_groupi_n_8048);
  xnor csa_tree_add_51_79_groupi_g37350(csa_tree_add_51_79_groupi_n_8813 ,csa_tree_add_51_79_groupi_n_7215 ,csa_tree_add_51_79_groupi_n_8092);
  xnor csa_tree_add_51_79_groupi_g37351(csa_tree_add_51_79_groupi_n_8812 ,csa_tree_add_51_79_groupi_n_7345 ,csa_tree_add_51_79_groupi_n_8047);
  xor csa_tree_add_51_79_groupi_g37352(csa_tree_add_51_79_groupi_n_8811 ,csa_tree_add_51_79_groupi_n_7593 ,csa_tree_add_51_79_groupi_n_8116);
  xnor csa_tree_add_51_79_groupi_g37353(csa_tree_add_51_79_groupi_n_8810 ,csa_tree_add_51_79_groupi_n_7805 ,csa_tree_add_51_79_groupi_n_8098);
  xnor csa_tree_add_51_79_groupi_g37354(csa_tree_add_51_79_groupi_n_8809 ,csa_tree_add_51_79_groupi_n_7290 ,csa_tree_add_51_79_groupi_n_8100);
  xnor csa_tree_add_51_79_groupi_g37355(csa_tree_add_51_79_groupi_n_8808 ,csa_tree_add_51_79_groupi_n_7148 ,csa_tree_add_51_79_groupi_n_8088);
  xnor csa_tree_add_51_79_groupi_g37356(csa_tree_add_51_79_groupi_n_8807 ,csa_tree_add_51_79_groupi_n_7341 ,csa_tree_add_51_79_groupi_n_8085);
  xnor csa_tree_add_51_79_groupi_g37357(csa_tree_add_51_79_groupi_n_8806 ,csa_tree_add_51_79_groupi_n_7339 ,csa_tree_add_51_79_groupi_n_8079);
  xnor csa_tree_add_51_79_groupi_g37358(csa_tree_add_51_79_groupi_n_8805 ,csa_tree_add_51_79_groupi_n_7201 ,csa_tree_add_51_79_groupi_n_8071);
  xnor csa_tree_add_51_79_groupi_g37359(csa_tree_add_51_79_groupi_n_8804 ,csa_tree_add_51_79_groupi_n_7293 ,csa_tree_add_51_79_groupi_n_8107);
  xnor csa_tree_add_51_79_groupi_g37360(csa_tree_add_51_79_groupi_n_8803 ,csa_tree_add_51_79_groupi_n_7381 ,csa_tree_add_51_79_groupi_n_8069);
  xnor csa_tree_add_51_79_groupi_g37361(csa_tree_add_51_79_groupi_n_8802 ,csa_tree_add_51_79_groupi_n_7633 ,csa_tree_add_51_79_groupi_n_8106);
  xnor csa_tree_add_51_79_groupi_g37362(csa_tree_add_51_79_groupi_n_8801 ,csa_tree_add_51_79_groupi_n_7347 ,csa_tree_add_51_79_groupi_n_8103);
  xnor csa_tree_add_51_79_groupi_g37363(csa_tree_add_51_79_groupi_n_8800 ,csa_tree_add_51_79_groupi_n_7182 ,csa_tree_add_51_79_groupi_n_8067);
  xnor csa_tree_add_51_79_groupi_g37364(csa_tree_add_51_79_groupi_n_8799 ,csa_tree_add_51_79_groupi_n_7328 ,csa_tree_add_51_79_groupi_n_8070);
  xnor csa_tree_add_51_79_groupi_g37365(csa_tree_add_51_79_groupi_n_8798 ,csa_tree_add_51_79_groupi_n_7318 ,csa_tree_add_51_79_groupi_n_8115);
  xnor csa_tree_add_51_79_groupi_g37366(csa_tree_add_51_79_groupi_n_8796 ,csa_tree_add_51_79_groupi_n_7152 ,csa_tree_add_51_79_groupi_n_8114);
  xnor csa_tree_add_51_79_groupi_g37367(csa_tree_add_51_79_groupi_n_8795 ,csa_tree_add_51_79_groupi_n_7829 ,csa_tree_add_51_79_groupi_n_8053);
  xnor csa_tree_add_51_79_groupi_g37368(csa_tree_add_51_79_groupi_n_8794 ,csa_tree_add_51_79_groupi_n_7327 ,csa_tree_add_51_79_groupi_n_8065);
  xnor csa_tree_add_51_79_groupi_g37369(csa_tree_add_51_79_groupi_n_8792 ,csa_tree_add_51_79_groupi_n_7621 ,csa_tree_add_51_79_groupi_n_8093);
  xnor csa_tree_add_51_79_groupi_g37370(csa_tree_add_51_79_groupi_n_8791 ,csa_tree_add_51_79_groupi_n_7314 ,csa_tree_add_51_79_groupi_n_8050);
  xnor csa_tree_add_51_79_groupi_g37371(csa_tree_add_51_79_groupi_n_8790 ,csa_tree_add_51_79_groupi_n_8340 ,csa_tree_add_51_79_groupi_n_8101);
  xnor csa_tree_add_51_79_groupi_g37372(csa_tree_add_51_79_groupi_n_8788 ,csa_tree_add_51_79_groupi_n_7276 ,csa_tree_add_51_79_groupi_n_8063);
  xnor csa_tree_add_51_79_groupi_g37373(csa_tree_add_51_79_groupi_n_8786 ,csa_tree_add_51_79_groupi_n_7311 ,csa_tree_add_51_79_groupi_n_8062);
  xnor csa_tree_add_51_79_groupi_g37374(csa_tree_add_51_79_groupi_n_8785 ,csa_tree_add_51_79_groupi_n_7309 ,csa_tree_add_51_79_groupi_n_8061);
  xnor csa_tree_add_51_79_groupi_g37375(csa_tree_add_51_79_groupi_n_8784 ,csa_tree_add_51_79_groupi_n_7316 ,csa_tree_add_51_79_groupi_n_8091);
  xnor csa_tree_add_51_79_groupi_g37376(csa_tree_add_51_79_groupi_n_8782 ,csa_tree_add_51_79_groupi_n_7145 ,csa_tree_add_51_79_groupi_n_8090);
  xnor csa_tree_add_51_79_groupi_g37377(csa_tree_add_51_79_groupi_n_8780 ,csa_tree_add_51_79_groupi_n_7367 ,csa_tree_add_51_79_groupi_n_8055);
  xnor csa_tree_add_51_79_groupi_g37378(csa_tree_add_51_79_groupi_n_8779 ,csa_tree_add_51_79_groupi_n_7259 ,csa_tree_add_51_79_groupi_n_8059);
  xnor csa_tree_add_51_79_groupi_g37379(csa_tree_add_51_79_groupi_n_8778 ,csa_tree_add_51_79_groupi_n_7166 ,csa_tree_add_51_79_groupi_n_8066);
  xnor csa_tree_add_51_79_groupi_g37380(csa_tree_add_51_79_groupi_n_8777 ,csa_tree_add_51_79_groupi_n_6720 ,csa_tree_add_51_79_groupi_n_8097);
  xnor csa_tree_add_51_79_groupi_g37381(csa_tree_add_51_79_groupi_n_8775 ,csa_tree_add_51_79_groupi_n_8184 ,csa_tree_add_51_79_groupi_n_8057);
  xnor csa_tree_add_51_79_groupi_g37382(csa_tree_add_51_79_groupi_n_8774 ,csa_tree_add_51_79_groupi_n_7344 ,csa_tree_add_51_79_groupi_n_8041);
  xnor csa_tree_add_51_79_groupi_g37383(csa_tree_add_51_79_groupi_n_8772 ,csa_tree_add_51_79_groupi_n_7161 ,csa_tree_add_51_79_groupi_n_8052);
  xnor csa_tree_add_51_79_groupi_g37384(csa_tree_add_51_79_groupi_n_8771 ,csa_tree_add_51_79_groupi_n_7343 ,csa_tree_add_51_79_groupi_n_8096);
  xnor csa_tree_add_51_79_groupi_g37385(csa_tree_add_51_79_groupi_n_8770 ,csa_tree_add_51_79_groupi_n_7307 ,csa_tree_add_51_79_groupi_n_8099);
  xnor csa_tree_add_51_79_groupi_g37386(csa_tree_add_51_79_groupi_n_8769 ,csa_tree_add_51_79_groupi_n_7141 ,csa_tree_add_51_79_groupi_n_8089);
  xnor csa_tree_add_51_79_groupi_g37387(csa_tree_add_51_79_groupi_n_8767 ,csa_tree_add_51_79_groupi_n_6428 ,csa_tree_add_51_79_groupi_n_8095);
  xnor csa_tree_add_51_79_groupi_g37388(csa_tree_add_51_79_groupi_n_8766 ,csa_tree_add_51_79_groupi_n_7596 ,csa_tree_add_51_79_groupi_n_8087);
  xnor csa_tree_add_51_79_groupi_g37389(csa_tree_add_51_79_groupi_n_8765 ,csa_tree_add_51_79_groupi_n_8027 ,csa_tree_add_51_79_groupi_n_8049);
  xnor csa_tree_add_51_79_groupi_g37390(csa_tree_add_51_79_groupi_n_8764 ,csa_tree_add_51_79_groupi_n_7149 ,csa_tree_add_51_79_groupi_n_8086);
  xnor csa_tree_add_51_79_groupi_g37391(csa_tree_add_51_79_groupi_n_8763 ,csa_tree_add_51_79_groupi_n_7219 ,csa_tree_add_51_79_groupi_n_8043);
  xnor csa_tree_add_51_79_groupi_g37392(csa_tree_add_51_79_groupi_n_8761 ,csa_tree_add_51_79_groupi_n_7281 ,csa_tree_add_51_79_groupi_n_8083);
  xnor csa_tree_add_51_79_groupi_g37393(csa_tree_add_51_79_groupi_n_8760 ,csa_tree_add_51_79_groupi_n_7165 ,csa_tree_add_51_79_groupi_n_8045);
  xnor csa_tree_add_51_79_groupi_g37394(csa_tree_add_51_79_groupi_n_8759 ,csa_tree_add_51_79_groupi_n_7257 ,csa_tree_add_51_79_groupi_n_8082);
  xnor csa_tree_add_51_79_groupi_g37395(csa_tree_add_51_79_groupi_n_8758 ,csa_tree_add_51_79_groupi_n_7102 ,csa_tree_add_51_79_groupi_n_8111);
  xnor csa_tree_add_51_79_groupi_g37396(csa_tree_add_51_79_groupi_n_8756 ,csa_tree_add_51_79_groupi_n_7142 ,csa_tree_add_51_79_groupi_n_8044);
  xnor csa_tree_add_51_79_groupi_g37397(csa_tree_add_51_79_groupi_n_8755 ,csa_tree_add_51_79_groupi_n_7263 ,csa_tree_add_51_79_groupi_n_8081);
  xnor csa_tree_add_51_79_groupi_g37398(csa_tree_add_51_79_groupi_n_8754 ,csa_tree_add_51_79_groupi_n_7139 ,csa_tree_add_51_79_groupi_n_8042);
  xnor csa_tree_add_51_79_groupi_g37399(csa_tree_add_51_79_groupi_n_8752 ,csa_tree_add_51_79_groupi_n_7631 ,csa_tree_add_51_79_groupi_n_8113);
  xnor csa_tree_add_51_79_groupi_g37400(csa_tree_add_51_79_groupi_n_8750 ,csa_tree_add_51_79_groupi_n_7385 ,csa_tree_add_51_79_groupi_n_8080);
  xnor csa_tree_add_51_79_groupi_g37401(csa_tree_add_51_79_groupi_n_8749 ,csa_tree_add_51_79_groupi_n_7329 ,csa_tree_add_51_79_groupi_n_8040);
  xnor csa_tree_add_51_79_groupi_g37402(csa_tree_add_51_79_groupi_n_8747 ,csa_tree_add_51_79_groupi_n_7228 ,csa_tree_add_51_79_groupi_n_8038);
  xnor csa_tree_add_51_79_groupi_g37403(csa_tree_add_51_79_groupi_n_8746 ,csa_tree_add_51_79_groupi_n_7211 ,csa_tree_add_51_79_groupi_n_8105);
  xnor csa_tree_add_51_79_groupi_g37404(csa_tree_add_51_79_groupi_n_8744 ,csa_tree_add_51_79_groupi_n_7226 ,csa_tree_add_51_79_groupi_n_8078);
  xnor csa_tree_add_51_79_groupi_g37405(csa_tree_add_51_79_groupi_n_8743 ,csa_tree_add_51_79_groupi_n_7576 ,csa_tree_add_51_79_groupi_n_8077);
  xnor csa_tree_add_51_79_groupi_g37406(csa_tree_add_51_79_groupi_n_8742 ,csa_tree_add_51_79_groupi_n_8313 ,csa_tree_add_51_79_groupi_n_8035);
  xnor csa_tree_add_51_79_groupi_g37407(csa_tree_add_51_79_groupi_n_8741 ,csa_tree_add_51_79_groupi_n_7212 ,csa_tree_add_51_79_groupi_n_8076);
  xnor csa_tree_add_51_79_groupi_g37408(csa_tree_add_51_79_groupi_n_8740 ,csa_tree_add_51_79_groupi_n_7235 ,csa_tree_add_51_79_groupi_n_8034);
  xnor csa_tree_add_51_79_groupi_g37409(csa_tree_add_51_79_groupi_n_8738 ,csa_tree_add_51_79_groupi_n_7580 ,csa_tree_add_51_79_groupi_n_8110);
  xnor csa_tree_add_51_79_groupi_g37410(csa_tree_add_51_79_groupi_n_8737 ,csa_tree_add_51_79_groupi_n_7614 ,csa_tree_add_51_79_groupi_n_8109);
  xnor csa_tree_add_51_79_groupi_g37411(csa_tree_add_51_79_groupi_n_8736 ,csa_tree_add_51_79_groupi_n_7245 ,csa_tree_add_51_79_groupi_n_8074);
  xnor csa_tree_add_51_79_groupi_g37412(csa_tree_add_51_79_groupi_n_8735 ,csa_tree_add_51_79_groupi_n_7582 ,csa_tree_add_51_79_groupi_n_8108);
  xnor csa_tree_add_51_79_groupi_g37413(csa_tree_add_51_79_groupi_n_8734 ,csa_tree_add_51_79_groupi_n_7334 ,csa_tree_add_51_79_groupi_n_8073);
  xnor csa_tree_add_51_79_groupi_g37414(csa_tree_add_51_79_groupi_n_8733 ,csa_tree_add_51_79_groupi_n_7207 ,csa_tree_add_51_79_groupi_n_8072);
  xnor csa_tree_add_51_79_groupi_g37415(csa_tree_add_51_79_groupi_n_8732 ,csa_tree_add_51_79_groupi_n_7247 ,csa_tree_add_51_79_groupi_n_8046);
  xnor csa_tree_add_51_79_groupi_g37416(csa_tree_add_51_79_groupi_n_8730 ,csa_tree_add_51_79_groupi_n_7379 ,csa_tree_add_51_79_groupi_n_8084);
  xnor csa_tree_add_51_79_groupi_g37417(csa_tree_add_51_79_groupi_n_8729 ,csa_tree_add_51_79_groupi_n_7377 ,csa_tree_add_51_79_groupi_n_8118);
  xnor csa_tree_add_51_79_groupi_g37418(csa_tree_add_51_79_groupi_n_8728 ,csa_tree_add_51_79_groupi_n_7185 ,csa_tree_add_51_79_groupi_n_8032);
  xnor csa_tree_add_51_79_groupi_g37419(csa_tree_add_51_79_groupi_n_8726 ,csa_tree_add_51_79_groupi_n_7196 ,csa_tree_add_51_79_groupi_n_8051);
  xnor csa_tree_add_51_79_groupi_g37420(csa_tree_add_51_79_groupi_n_8725 ,csa_tree_add_51_79_groupi_n_7289 ,csa_tree_add_51_79_groupi_n_8039);
  xnor csa_tree_add_51_79_groupi_g37421(csa_tree_add_51_79_groupi_n_8723 ,csa_tree_add_51_79_groupi_n_7190 ,csa_tree_add_51_79_groupi_n_8068);
  xnor csa_tree_add_51_79_groupi_g37422(csa_tree_add_51_79_groupi_n_8722 ,csa_tree_add_51_79_groupi_n_7605 ,csa_tree_add_51_79_groupi_n_8104);
  xnor csa_tree_add_51_79_groupi_g37423(csa_tree_add_51_79_groupi_n_8721 ,csa_tree_add_51_79_groupi_n_7336 ,csa_tree_add_51_79_groupi_n_8117);
  xnor csa_tree_add_51_79_groupi_g37424(csa_tree_add_51_79_groupi_n_8720 ,csa_tree_add_51_79_groupi_n_7326 ,csa_tree_add_51_79_groupi_n_8094);
  xnor csa_tree_add_51_79_groupi_g37425(csa_tree_add_51_79_groupi_n_8719 ,csa_tree_add_51_79_groupi_n_7619 ,csa_tree_add_51_79_groupi_n_8037);
  and csa_tree_add_51_79_groupi_g37426(csa_tree_add_51_79_groupi_n_8717 ,csa_tree_add_51_79_groupi_n_8138 ,csa_tree_add_51_79_groupi_n_8360);
  not csa_tree_add_51_79_groupi_g37428(csa_tree_add_51_79_groupi_n_8647 ,csa_tree_add_51_79_groupi_n_8646);
  not csa_tree_add_51_79_groupi_g37429(csa_tree_add_51_79_groupi_n_8627 ,csa_tree_add_51_79_groupi_n_8626);
  not csa_tree_add_51_79_groupi_g37430(csa_tree_add_51_79_groupi_n_8621 ,csa_tree_add_51_79_groupi_n_8622);
  not csa_tree_add_51_79_groupi_g37431(csa_tree_add_51_79_groupi_n_8620 ,csa_tree_add_51_79_groupi_n_8619);
  not csa_tree_add_51_79_groupi_g37432(csa_tree_add_51_79_groupi_n_8617 ,csa_tree_add_51_79_groupi_n_8618);
  not csa_tree_add_51_79_groupi_g37433(csa_tree_add_51_79_groupi_n_8612 ,csa_tree_add_51_79_groupi_n_8613);
  not csa_tree_add_51_79_groupi_g37434(csa_tree_add_51_79_groupi_n_8608 ,csa_tree_add_51_79_groupi_n_8609);
  not csa_tree_add_51_79_groupi_g37435(csa_tree_add_51_79_groupi_n_8606 ,csa_tree_add_51_79_groupi_n_8605);
  not csa_tree_add_51_79_groupi_g37436(csa_tree_add_51_79_groupi_n_8602 ,csa_tree_add_51_79_groupi_n_8603);
  not csa_tree_add_51_79_groupi_g37437(csa_tree_add_51_79_groupi_n_8600 ,csa_tree_add_51_79_groupi_n_8599);
  not csa_tree_add_51_79_groupi_g37438(csa_tree_add_51_79_groupi_n_8598 ,csa_tree_add_51_79_groupi_n_8597);
  not csa_tree_add_51_79_groupi_g37439(csa_tree_add_51_79_groupi_n_8595 ,csa_tree_add_51_79_groupi_n_8596);
  not csa_tree_add_51_79_groupi_g37440(csa_tree_add_51_79_groupi_n_8592 ,csa_tree_add_51_79_groupi_n_8591);
  not csa_tree_add_51_79_groupi_g37441(csa_tree_add_51_79_groupi_n_8587 ,csa_tree_add_51_79_groupi_n_8588);
  not csa_tree_add_51_79_groupi_g37442(csa_tree_add_51_79_groupi_n_8586 ,csa_tree_add_51_79_groupi_n_8585);
  not csa_tree_add_51_79_groupi_g37443(csa_tree_add_51_79_groupi_n_8583 ,csa_tree_add_51_79_groupi_n_8584);
  not csa_tree_add_51_79_groupi_g37444(csa_tree_add_51_79_groupi_n_8580 ,csa_tree_add_51_79_groupi_n_8581);
  not csa_tree_add_51_79_groupi_g37445(csa_tree_add_51_79_groupi_n_8577 ,csa_tree_add_51_79_groupi_n_8578);
  not csa_tree_add_51_79_groupi_g37446(csa_tree_add_51_79_groupi_n_8575 ,csa_tree_add_51_79_groupi_n_8576);
  not csa_tree_add_51_79_groupi_g37447(csa_tree_add_51_79_groupi_n_8573 ,csa_tree_add_51_79_groupi_n_8574);
  not csa_tree_add_51_79_groupi_g37448(csa_tree_add_51_79_groupi_n_8570 ,csa_tree_add_51_79_groupi_n_8571);
  not csa_tree_add_51_79_groupi_g37449(csa_tree_add_51_79_groupi_n_8568 ,csa_tree_add_51_79_groupi_n_8569);
  or csa_tree_add_51_79_groupi_g37450(csa_tree_add_51_79_groupi_n_8566 ,csa_tree_add_51_79_groupi_n_7901 ,csa_tree_add_51_79_groupi_n_8340);
  and csa_tree_add_51_79_groupi_g37451(csa_tree_add_51_79_groupi_n_8565 ,csa_tree_add_51_79_groupi_n_8017 ,csa_tree_add_51_79_groupi_n_8302);
  or csa_tree_add_51_79_groupi_g37452(csa_tree_add_51_79_groupi_n_8564 ,csa_tree_add_51_79_groupi_n_8011 ,csa_tree_add_51_79_groupi_n_8313);
  or csa_tree_add_51_79_groupi_g37453(csa_tree_add_51_79_groupi_n_8563 ,csa_tree_add_51_79_groupi_n_8277 ,csa_tree_add_51_79_groupi_n_8279);
  or csa_tree_add_51_79_groupi_g37454(csa_tree_add_51_79_groupi_n_8562 ,csa_tree_add_51_79_groupi_n_7249 ,csa_tree_add_51_79_groupi_n_8278);
  nor csa_tree_add_51_79_groupi_g37455(csa_tree_add_51_79_groupi_n_8561 ,csa_tree_add_51_79_groupi_n_8282 ,csa_tree_add_51_79_groupi_n_8275);
  and csa_tree_add_51_79_groupi_g37456(csa_tree_add_51_79_groupi_n_8560 ,csa_tree_add_51_79_groupi_n_8277 ,csa_tree_add_51_79_groupi_n_8279);
  and csa_tree_add_51_79_groupi_g37457(csa_tree_add_51_79_groupi_n_8559 ,csa_tree_add_51_79_groupi_n_8175 ,csa_tree_add_51_79_groupi_n_8151);
  or csa_tree_add_51_79_groupi_g37458(csa_tree_add_51_79_groupi_n_8558 ,csa_tree_add_51_79_groupi_n_8289 ,csa_tree_add_51_79_groupi_n_8290);
  and csa_tree_add_51_79_groupi_g37459(csa_tree_add_51_79_groupi_n_8557 ,csa_tree_add_51_79_groupi_n_7249 ,csa_tree_add_51_79_groupi_n_8278);
  or csa_tree_add_51_79_groupi_g37460(csa_tree_add_51_79_groupi_n_8556 ,csa_tree_add_51_79_groupi_n_8251 ,csa_tree_add_51_79_groupi_n_7834);
  or csa_tree_add_51_79_groupi_g37461(csa_tree_add_51_79_groupi_n_8555 ,csa_tree_add_51_79_groupi_n_8175 ,csa_tree_add_51_79_groupi_n_8151);
  or csa_tree_add_51_79_groupi_g37462(csa_tree_add_51_79_groupi_n_8554 ,csa_tree_add_51_79_groupi_n_8160 ,csa_tree_add_51_79_groupi_n_8276);
  and csa_tree_add_51_79_groupi_g37463(csa_tree_add_51_79_groupi_n_8553 ,csa_tree_add_51_79_groupi_n_8289 ,csa_tree_add_51_79_groupi_n_8290);
  or csa_tree_add_51_79_groupi_g37464(csa_tree_add_51_79_groupi_n_8552 ,csa_tree_add_51_79_groupi_n_8169 ,csa_tree_add_51_79_groupi_n_8293);
  and csa_tree_add_51_79_groupi_g37465(csa_tree_add_51_79_groupi_n_8551 ,csa_tree_add_51_79_groupi_n_8160 ,csa_tree_add_51_79_groupi_n_8276);
  and csa_tree_add_51_79_groupi_g37466(csa_tree_add_51_79_groupi_n_8550 ,csa_tree_add_51_79_groupi_n_8169 ,csa_tree_add_51_79_groupi_n_8293);
  and csa_tree_add_51_79_groupi_g37467(csa_tree_add_51_79_groupi_n_8549 ,csa_tree_add_51_79_groupi_n_8161 ,csa_tree_add_51_79_groupi_n_8292);
  or csa_tree_add_51_79_groupi_g37468(csa_tree_add_51_79_groupi_n_8548 ,csa_tree_add_51_79_groupi_n_8161 ,csa_tree_add_51_79_groupi_n_8292);
  or csa_tree_add_51_79_groupi_g37469(csa_tree_add_51_79_groupi_n_8547 ,csa_tree_add_51_79_groupi_n_7831 ,csa_tree_add_51_79_groupi_n_8140);
  or csa_tree_add_51_79_groupi_g37470(csa_tree_add_51_79_groupi_n_8546 ,csa_tree_add_51_79_groupi_n_8297 ,csa_tree_add_51_79_groupi_n_8300);
  or csa_tree_add_51_79_groupi_g37471(csa_tree_add_51_79_groupi_n_8545 ,csa_tree_add_51_79_groupi_n_7319 ,csa_tree_add_51_79_groupi_n_8149);
  or csa_tree_add_51_79_groupi_g37472(csa_tree_add_51_79_groupi_n_8544 ,csa_tree_add_51_79_groupi_n_8121 ,csa_tree_add_51_79_groupi_n_8322);
  nor csa_tree_add_51_79_groupi_g37473(csa_tree_add_51_79_groupi_n_8543 ,csa_tree_add_51_79_groupi_n_7597 ,csa_tree_add_51_79_groupi_n_8272);
  or csa_tree_add_51_79_groupi_g37474(csa_tree_add_51_79_groupi_n_8542 ,csa_tree_add_51_79_groupi_n_8308 ,csa_tree_add_51_79_groupi_n_8310);
  and csa_tree_add_51_79_groupi_g37475(csa_tree_add_51_79_groupi_n_8541 ,csa_tree_add_51_79_groupi_n_7804 ,csa_tree_add_51_79_groupi_n_8273);
  or csa_tree_add_51_79_groupi_g37476(csa_tree_add_51_79_groupi_n_8540 ,csa_tree_add_51_79_groupi_n_7598 ,csa_tree_add_51_79_groupi_n_8271);
  and csa_tree_add_51_79_groupi_g37477(csa_tree_add_51_79_groupi_n_8539 ,csa_tree_add_51_79_groupi_n_8297 ,csa_tree_add_51_79_groupi_n_8300);
  or csa_tree_add_51_79_groupi_g37478(csa_tree_add_51_79_groupi_n_8538 ,csa_tree_add_51_79_groupi_n_7804 ,csa_tree_add_51_79_groupi_n_8273);
  and csa_tree_add_51_79_groupi_g37479(csa_tree_add_51_79_groupi_n_8537 ,csa_tree_add_51_79_groupi_n_8308 ,csa_tree_add_51_79_groupi_n_8310);
  and csa_tree_add_51_79_groupi_g37480(csa_tree_add_51_79_groupi_n_8536 ,csa_tree_add_51_79_groupi_n_7803 ,csa_tree_add_51_79_groupi_n_8283);
  and csa_tree_add_51_79_groupi_g37481(csa_tree_add_51_79_groupi_n_8535 ,csa_tree_add_51_79_groupi_n_8296 ,csa_tree_add_51_79_groupi_n_8288);
  or csa_tree_add_51_79_groupi_g37482(csa_tree_add_51_79_groupi_n_8534 ,csa_tree_add_51_79_groupi_n_8281 ,csa_tree_add_51_79_groupi_n_8274);
  or csa_tree_add_51_79_groupi_g37483(csa_tree_add_51_79_groupi_n_8533 ,csa_tree_add_51_79_groupi_n_7803 ,csa_tree_add_51_79_groupi_n_8283);
  or csa_tree_add_51_79_groupi_g37484(csa_tree_add_51_79_groupi_n_8532 ,csa_tree_add_51_79_groupi_n_8319 ,csa_tree_add_51_79_groupi_n_8257);
  or csa_tree_add_51_79_groupi_g37485(csa_tree_add_51_79_groupi_n_8531 ,csa_tree_add_51_79_groupi_n_7627 ,csa_tree_add_51_79_groupi_n_8144);
  or csa_tree_add_51_79_groupi_g37486(csa_tree_add_51_79_groupi_n_8530 ,csa_tree_add_51_79_groupi_n_8296 ,csa_tree_add_51_79_groupi_n_8288);
  or csa_tree_add_51_79_groupi_g37487(csa_tree_add_51_79_groupi_n_8529 ,csa_tree_add_51_79_groupi_n_7844 ,csa_tree_add_51_79_groupi_n_8184);
  or csa_tree_add_51_79_groupi_g37488(csa_tree_add_51_79_groupi_n_8528 ,csa_tree_add_51_79_groupi_n_6854 ,csa_tree_add_51_79_groupi_n_8267);
  and csa_tree_add_51_79_groupi_g37489(csa_tree_add_51_79_groupi_n_8527 ,csa_tree_add_51_79_groupi_n_8265 ,csa_tree_add_51_79_groupi_n_8298);
  or csa_tree_add_51_79_groupi_g37490(csa_tree_add_51_79_groupi_n_8526 ,csa_tree_add_51_79_groupi_n_8179 ,csa_tree_add_51_79_groupi_n_8235);
  and csa_tree_add_51_79_groupi_g37491(csa_tree_add_51_79_groupi_n_8525 ,csa_tree_add_51_79_groupi_n_7628 ,csa_tree_add_51_79_groupi_n_8213);
  or csa_tree_add_51_79_groupi_g37492(csa_tree_add_51_79_groupi_n_8524 ,csa_tree_add_51_79_groupi_n_8017 ,csa_tree_add_51_79_groupi_n_8302);
  and csa_tree_add_51_79_groupi_g37493(csa_tree_add_51_79_groupi_n_8523 ,csa_tree_add_51_79_groupi_n_8311 ,csa_tree_add_51_79_groupi_n_8309);
  or csa_tree_add_51_79_groupi_g37494(csa_tree_add_51_79_groupi_n_8522 ,csa_tree_add_51_79_groupi_n_8280 ,csa_tree_add_51_79_groupi_n_8287);
  or csa_tree_add_51_79_groupi_g37495(csa_tree_add_51_79_groupi_n_8521 ,csa_tree_add_51_79_groupi_n_8285 ,csa_tree_add_51_79_groupi_n_7825);
  nor csa_tree_add_51_79_groupi_g37496(csa_tree_add_51_79_groupi_n_8520 ,csa_tree_add_51_79_groupi_n_7301 ,csa_tree_add_51_79_groupi_n_8295);
  nor csa_tree_add_51_79_groupi_g37497(csa_tree_add_51_79_groupi_n_8519 ,csa_tree_add_51_79_groupi_n_6855 ,csa_tree_add_51_79_groupi_n_8266);
  and csa_tree_add_51_79_groupi_g37498(csa_tree_add_51_79_groupi_n_8518 ,csa_tree_add_51_79_groupi_n_8280 ,csa_tree_add_51_79_groupi_n_8287);
  or csa_tree_add_51_79_groupi_g37499(csa_tree_add_51_79_groupi_n_8517 ,csa_tree_add_51_79_groupi_n_7380 ,csa_tree_add_51_79_groupi_n_8200);
  or csa_tree_add_51_79_groupi_g37500(csa_tree_add_51_79_groupi_n_8516 ,csa_tree_add_51_79_groupi_n_8311 ,csa_tree_add_51_79_groupi_n_8309);
  or csa_tree_add_51_79_groupi_g37501(csa_tree_add_51_79_groupi_n_8515 ,csa_tree_add_51_79_groupi_n_8265 ,csa_tree_add_51_79_groupi_n_8298);
  nor csa_tree_add_51_79_groupi_g37502(csa_tree_add_51_79_groupi_n_8514 ,csa_tree_add_51_79_groupi_n_7607 ,csa_tree_add_51_79_groupi_n_8306);
  or csa_tree_add_51_79_groupi_g37503(csa_tree_add_51_79_groupi_n_8513 ,csa_tree_add_51_79_groupi_n_7300 ,csa_tree_add_51_79_groupi_n_8294);
  and csa_tree_add_51_79_groupi_g37504(csa_tree_add_51_79_groupi_n_8512 ,csa_tree_add_51_79_groupi_n_8285 ,csa_tree_add_51_79_groupi_n_7825);
  and csa_tree_add_51_79_groupi_g37505(csa_tree_add_51_79_groupi_n_8511 ,csa_tree_add_51_79_groupi_n_8268 ,csa_tree_add_51_79_groupi_n_8301);
  and csa_tree_add_51_79_groupi_g37506(csa_tree_add_51_79_groupi_n_8510 ,csa_tree_add_51_79_groupi_n_8284 ,csa_tree_add_51_79_groupi_n_8299);
  or csa_tree_add_51_79_groupi_g37507(csa_tree_add_51_79_groupi_n_8509 ,csa_tree_add_51_79_groupi_n_7606 ,csa_tree_add_51_79_groupi_n_8307);
  or csa_tree_add_51_79_groupi_g37508(csa_tree_add_51_79_groupi_n_8508 ,csa_tree_add_51_79_groupi_n_8268 ,csa_tree_add_51_79_groupi_n_8301);
  or csa_tree_add_51_79_groupi_g37509(csa_tree_add_51_79_groupi_n_8507 ,csa_tree_add_51_79_groupi_n_8284 ,csa_tree_add_51_79_groupi_n_8299);
  and csa_tree_add_51_79_groupi_g37510(csa_tree_add_51_79_groupi_n_8658 ,csa_tree_add_51_79_groupi_n_8005 ,csa_tree_add_51_79_groupi_n_8256);
  and csa_tree_add_51_79_groupi_g37511(csa_tree_add_51_79_groupi_n_8657 ,csa_tree_add_51_79_groupi_n_7996 ,csa_tree_add_51_79_groupi_n_8247);
  and csa_tree_add_51_79_groupi_g37512(csa_tree_add_51_79_groupi_n_8656 ,csa_tree_add_51_79_groupi_n_7756 ,csa_tree_add_51_79_groupi_n_8187);
  and csa_tree_add_51_79_groupi_g37513(csa_tree_add_51_79_groupi_n_8655 ,csa_tree_add_51_79_groupi_n_7912 ,csa_tree_add_51_79_groupi_n_8191);
  and csa_tree_add_51_79_groupi_g37514(csa_tree_add_51_79_groupi_n_8654 ,csa_tree_add_51_79_groupi_n_7989 ,csa_tree_add_51_79_groupi_n_8244);
  and csa_tree_add_51_79_groupi_g37515(csa_tree_add_51_79_groupi_n_8653 ,csa_tree_add_51_79_groupi_n_7987 ,csa_tree_add_51_79_groupi_n_8242);
  and csa_tree_add_51_79_groupi_g37516(csa_tree_add_51_79_groupi_n_8652 ,csa_tree_add_51_79_groupi_n_7982 ,csa_tree_add_51_79_groupi_n_8239);
  and csa_tree_add_51_79_groupi_g37517(csa_tree_add_51_79_groupi_n_8651 ,csa_tree_add_51_79_groupi_n_7950 ,csa_tree_add_51_79_groupi_n_8143);
  and csa_tree_add_51_79_groupi_g37518(csa_tree_add_51_79_groupi_n_8650 ,csa_tree_add_51_79_groupi_n_7785 ,csa_tree_add_51_79_groupi_n_8264);
  or csa_tree_add_51_79_groupi_g37519(csa_tree_add_51_79_groupi_n_8649 ,csa_tree_add_51_79_groupi_n_7887 ,csa_tree_add_51_79_groupi_n_8195);
  and csa_tree_add_51_79_groupi_g37520(csa_tree_add_51_79_groupi_n_8648 ,csa_tree_add_51_79_groupi_n_7791 ,csa_tree_add_51_79_groupi_n_8147);
  or csa_tree_add_51_79_groupi_g37521(csa_tree_add_51_79_groupi_n_8646 ,csa_tree_add_51_79_groupi_n_7947 ,csa_tree_add_51_79_groupi_n_8189);
  and csa_tree_add_51_79_groupi_g37522(csa_tree_add_51_79_groupi_n_8645 ,csa_tree_add_51_79_groupi_n_7882 ,csa_tree_add_51_79_groupi_n_8204);
  and csa_tree_add_51_79_groupi_g37523(csa_tree_add_51_79_groupi_n_8644 ,csa_tree_add_51_79_groupi_n_7880 ,csa_tree_add_51_79_groupi_n_8209);
  and csa_tree_add_51_79_groupi_g37524(csa_tree_add_51_79_groupi_n_8643 ,csa_tree_add_51_79_groupi_n_7794 ,csa_tree_add_51_79_groupi_n_8150);
  and csa_tree_add_51_79_groupi_g37525(csa_tree_add_51_79_groupi_n_8642 ,csa_tree_add_51_79_groupi_n_7878 ,csa_tree_add_51_79_groupi_n_8206);
  and csa_tree_add_51_79_groupi_g37526(csa_tree_add_51_79_groupi_n_8641 ,csa_tree_add_51_79_groupi_n_7877 ,csa_tree_add_51_79_groupi_n_8207);
  and csa_tree_add_51_79_groupi_g37527(csa_tree_add_51_79_groupi_n_8640 ,csa_tree_add_51_79_groupi_n_7965 ,csa_tree_add_51_79_groupi_n_8227);
  and csa_tree_add_51_79_groupi_g37528(csa_tree_add_51_79_groupi_n_8639 ,csa_tree_add_51_79_groupi_n_7921 ,csa_tree_add_51_79_groupi_n_8196);
  and csa_tree_add_51_79_groupi_g37529(csa_tree_add_51_79_groupi_n_8638 ,csa_tree_add_51_79_groupi_n_8002 ,csa_tree_add_51_79_groupi_n_8261);
  and csa_tree_add_51_79_groupi_g37530(csa_tree_add_51_79_groupi_n_8637 ,csa_tree_add_51_79_groupi_n_7865 ,csa_tree_add_51_79_groupi_n_8229);
  and csa_tree_add_51_79_groupi_g37531(csa_tree_add_51_79_groupi_n_8636 ,csa_tree_add_51_79_groupi_n_7899 ,csa_tree_add_51_79_groupi_n_8260);
  and csa_tree_add_51_79_groupi_g37532(csa_tree_add_51_79_groupi_n_8635 ,csa_tree_add_51_79_groupi_n_7862 ,csa_tree_add_51_79_groupi_n_8232);
  and csa_tree_add_51_79_groupi_g37533(csa_tree_add_51_79_groupi_n_8634 ,csa_tree_add_51_79_groupi_n_7959 ,csa_tree_add_51_79_groupi_n_8223);
  or csa_tree_add_51_79_groupi_g37534(csa_tree_add_51_79_groupi_n_8633 ,csa_tree_add_51_79_groupi_n_7957 ,csa_tree_add_51_79_groupi_n_8221);
  and csa_tree_add_51_79_groupi_g37535(csa_tree_add_51_79_groupi_n_8632 ,csa_tree_add_51_79_groupi_n_7924 ,csa_tree_add_51_79_groupi_n_8197);
  and csa_tree_add_51_79_groupi_g37536(csa_tree_add_51_79_groupi_n_8631 ,csa_tree_add_51_79_groupi_n_7929 ,csa_tree_add_51_79_groupi_n_8199);
  and csa_tree_add_51_79_groupi_g37537(csa_tree_add_51_79_groupi_n_8630 ,csa_tree_add_51_79_groupi_n_7857 ,csa_tree_add_51_79_groupi_n_8233);
  and csa_tree_add_51_79_groupi_g37538(csa_tree_add_51_79_groupi_n_8629 ,csa_tree_add_51_79_groupi_n_7931 ,csa_tree_add_51_79_groupi_n_8203);
  and csa_tree_add_51_79_groupi_g37539(csa_tree_add_51_79_groupi_n_8628 ,csa_tree_add_51_79_groupi_n_7955 ,csa_tree_add_51_79_groupi_n_8220);
  or csa_tree_add_51_79_groupi_g37540(csa_tree_add_51_79_groupi_n_8626 ,csa_tree_add_51_79_groupi_n_7838 ,csa_tree_add_51_79_groupi_n_8253);
  and csa_tree_add_51_79_groupi_g37541(csa_tree_add_51_79_groupi_n_8625 ,csa_tree_add_51_79_groupi_n_7943 ,csa_tree_add_51_79_groupi_n_8215);
  and csa_tree_add_51_79_groupi_g37542(csa_tree_add_51_79_groupi_n_8624 ,csa_tree_add_51_79_groupi_n_7840 ,csa_tree_add_51_79_groupi_n_8188);
  and csa_tree_add_51_79_groupi_g37543(csa_tree_add_51_79_groupi_n_8623 ,csa_tree_add_51_79_groupi_n_7802 ,csa_tree_add_51_79_groupi_n_8216);
  and csa_tree_add_51_79_groupi_g37544(csa_tree_add_51_79_groupi_n_8622 ,csa_tree_add_51_79_groupi_n_7797 ,csa_tree_add_51_79_groupi_n_8263);
  and csa_tree_add_51_79_groupi_g37545(csa_tree_add_51_79_groupi_n_8619 ,csa_tree_add_51_79_groupi_n_7841 ,csa_tree_add_51_79_groupi_n_8246);
  or csa_tree_add_51_79_groupi_g37546(csa_tree_add_51_79_groupi_n_8618 ,csa_tree_add_51_79_groupi_n_8013 ,csa_tree_add_51_79_groupi_n_8249);
  and csa_tree_add_51_79_groupi_g37547(csa_tree_add_51_79_groupi_n_8616 ,csa_tree_add_51_79_groupi_n_7778 ,csa_tree_add_51_79_groupi_n_8211);
  or csa_tree_add_51_79_groupi_g37548(csa_tree_add_51_79_groupi_n_8615 ,csa_tree_add_51_79_groupi_n_7951 ,csa_tree_add_51_79_groupi_n_8218);
  or csa_tree_add_51_79_groupi_g37549(csa_tree_add_51_79_groupi_n_8614 ,csa_tree_add_51_79_groupi_n_7942 ,csa_tree_add_51_79_groupi_n_8214);
  and csa_tree_add_51_79_groupi_g37550(csa_tree_add_51_79_groupi_n_8613 ,csa_tree_add_51_79_groupi_n_7728 ,csa_tree_add_51_79_groupi_n_8222);
  and csa_tree_add_51_79_groupi_g37551(csa_tree_add_51_79_groupi_n_8611 ,csa_tree_add_51_79_groupi_n_7923 ,csa_tree_add_51_79_groupi_n_8198);
  and csa_tree_add_51_79_groupi_g37552(csa_tree_add_51_79_groupi_n_8610 ,csa_tree_add_51_79_groupi_n_7765 ,csa_tree_add_51_79_groupi_n_8225);
  and csa_tree_add_51_79_groupi_g37553(csa_tree_add_51_79_groupi_n_8609 ,csa_tree_add_51_79_groupi_n_7961 ,csa_tree_add_51_79_groupi_n_8224);
  and csa_tree_add_51_79_groupi_g37554(csa_tree_add_51_79_groupi_n_8607 ,csa_tree_add_51_79_groupi_n_7896 ,csa_tree_add_51_79_groupi_n_8258);
  and csa_tree_add_51_79_groupi_g37555(csa_tree_add_51_79_groupi_n_8605 ,csa_tree_add_51_79_groupi_n_7784 ,csa_tree_add_51_79_groupi_n_8230);
  and csa_tree_add_51_79_groupi_g37556(csa_tree_add_51_79_groupi_n_8604 ,csa_tree_add_51_79_groupi_n_7934 ,csa_tree_add_51_79_groupi_n_8259);
  or csa_tree_add_51_79_groupi_g37557(csa_tree_add_51_79_groupi_n_8603 ,csa_tree_add_51_79_groupi_n_7866 ,csa_tree_add_51_79_groupi_n_8219);
  and csa_tree_add_51_79_groupi_g37558(csa_tree_add_51_79_groupi_n_8601 ,csa_tree_add_51_79_groupi_n_7782 ,csa_tree_add_51_79_groupi_n_8226);
  and csa_tree_add_51_79_groupi_g37559(csa_tree_add_51_79_groupi_n_8599 ,csa_tree_add_51_79_groupi_n_7966 ,csa_tree_add_51_79_groupi_n_8228);
  and csa_tree_add_51_79_groupi_g37560(csa_tree_add_51_79_groupi_n_8597 ,csa_tree_add_51_79_groupi_n_7873 ,csa_tree_add_51_79_groupi_n_8212);
  or csa_tree_add_51_79_groupi_g37561(csa_tree_add_51_79_groupi_n_8596 ,csa_tree_add_51_79_groupi_n_7971 ,csa_tree_add_51_79_groupi_n_8231);
  and csa_tree_add_51_79_groupi_g37562(csa_tree_add_51_79_groupi_n_8594 ,csa_tree_add_51_79_groupi_n_7946 ,csa_tree_add_51_79_groupi_n_8217);
  and csa_tree_add_51_79_groupi_g37563(csa_tree_add_51_79_groupi_n_8593 ,csa_tree_add_51_79_groupi_n_7979 ,csa_tree_add_51_79_groupi_n_8238);
  and csa_tree_add_51_79_groupi_g37564(csa_tree_add_51_79_groupi_n_8591 ,csa_tree_add_51_79_groupi_n_7875 ,csa_tree_add_51_79_groupi_n_8208);
  and csa_tree_add_51_79_groupi_g37565(csa_tree_add_51_79_groupi_n_8590 ,csa_tree_add_51_79_groupi_n_7793 ,csa_tree_add_51_79_groupi_n_8148);
  and csa_tree_add_51_79_groupi_g37566(csa_tree_add_51_79_groupi_n_8589 ,csa_tree_add_51_79_groupi_n_7751 ,csa_tree_add_51_79_groupi_n_8205);
  or csa_tree_add_51_79_groupi_g37567(csa_tree_add_51_79_groupi_n_8588 ,csa_tree_add_51_79_groupi_n_7788 ,csa_tree_add_51_79_groupi_n_8146);
  and csa_tree_add_51_79_groupi_g37568(csa_tree_add_51_79_groupi_n_8585 ,csa_tree_add_51_79_groupi_n_7886 ,csa_tree_add_51_79_groupi_n_8201);
  or csa_tree_add_51_79_groupi_g37569(csa_tree_add_51_79_groupi_n_8584 ,csa_tree_add_51_79_groupi_n_7889 ,csa_tree_add_51_79_groupi_n_8192);
  and csa_tree_add_51_79_groupi_g37570(csa_tree_add_51_79_groupi_n_8582 ,csa_tree_add_51_79_groupi_n_7780 ,csa_tree_add_51_79_groupi_n_8142);
  or csa_tree_add_51_79_groupi_g37571(csa_tree_add_51_79_groupi_n_8581 ,csa_tree_add_51_79_groupi_n_7917 ,csa_tree_add_51_79_groupi_n_8194);
  and csa_tree_add_51_79_groupi_g37572(csa_tree_add_51_79_groupi_n_8579 ,csa_tree_add_51_79_groupi_n_7984 ,csa_tree_add_51_79_groupi_n_8241);
  and csa_tree_add_51_79_groupi_g37573(csa_tree_add_51_79_groupi_n_8578 ,csa_tree_add_51_79_groupi_n_8008 ,csa_tree_add_51_79_groupi_n_8190);
  or csa_tree_add_51_79_groupi_g37574(csa_tree_add_51_79_groupi_n_8576 ,csa_tree_add_51_79_groupi_n_7915 ,csa_tree_add_51_79_groupi_n_8193);
  or csa_tree_add_51_79_groupi_g37575(csa_tree_add_51_79_groupi_n_8574 ,csa_tree_add_51_79_groupi_n_7993 ,csa_tree_add_51_79_groupi_n_8245);
  and csa_tree_add_51_79_groupi_g37576(csa_tree_add_51_79_groupi_n_8572 ,csa_tree_add_51_79_groupi_n_7770 ,csa_tree_add_51_79_groupi_n_8262);
  or csa_tree_add_51_79_groupi_g37577(csa_tree_add_51_79_groupi_n_8571 ,csa_tree_add_51_79_groupi_n_7999 ,csa_tree_add_51_79_groupi_n_8248);
  and csa_tree_add_51_79_groupi_g37578(csa_tree_add_51_79_groupi_n_8569 ,csa_tree_add_51_79_groupi_n_7976 ,csa_tree_add_51_79_groupi_n_8243);
  and csa_tree_add_51_79_groupi_g37579(csa_tree_add_51_79_groupi_n_8567 ,csa_tree_add_51_79_groupi_n_7906 ,csa_tree_add_51_79_groupi_n_8186);
  not csa_tree_add_51_79_groupi_g37580(csa_tree_add_51_79_groupi_n_8504 ,csa_tree_add_51_79_groupi_n_8503);
  not csa_tree_add_51_79_groupi_g37581(csa_tree_add_51_79_groupi_n_8500 ,csa_tree_add_51_79_groupi_n_8499);
  not csa_tree_add_51_79_groupi_g37582(csa_tree_add_51_79_groupi_n_8493 ,csa_tree_add_51_79_groupi_n_8492);
  not csa_tree_add_51_79_groupi_g37583(csa_tree_add_51_79_groupi_n_8484 ,csa_tree_add_51_79_groupi_n_8483);
  not csa_tree_add_51_79_groupi_g37584(csa_tree_add_51_79_groupi_n_8482 ,csa_tree_add_51_79_groupi_n_8481);
  not csa_tree_add_51_79_groupi_g37585(csa_tree_add_51_79_groupi_n_8478 ,csa_tree_add_51_79_groupi_n_8479);
  not csa_tree_add_51_79_groupi_g37586(csa_tree_add_51_79_groupi_n_8476 ,csa_tree_add_51_79_groupi_n_8477);
  not csa_tree_add_51_79_groupi_g37587(csa_tree_add_51_79_groupi_n_8471 ,csa_tree_add_51_79_groupi_n_8470);
  not csa_tree_add_51_79_groupi_g37588(csa_tree_add_51_79_groupi_n_8469 ,csa_tree_add_51_79_groupi_n_8468);
  not csa_tree_add_51_79_groupi_g37589(csa_tree_add_51_79_groupi_n_8467 ,csa_tree_add_51_79_groupi_n_8466);
  not csa_tree_add_51_79_groupi_g37590(csa_tree_add_51_79_groupi_n_8463 ,csa_tree_add_51_79_groupi_n_8464);
  not csa_tree_add_51_79_groupi_g37591(csa_tree_add_51_79_groupi_n_8458 ,csa_tree_add_51_79_groupi_n_8459);
  not csa_tree_add_51_79_groupi_g37592(csa_tree_add_51_79_groupi_n_8457 ,csa_tree_add_51_79_groupi_n_8456);
  not csa_tree_add_51_79_groupi_g37593(csa_tree_add_51_79_groupi_n_8455 ,csa_tree_add_51_79_groupi_n_8454);
  not csa_tree_add_51_79_groupi_g37594(csa_tree_add_51_79_groupi_n_8451 ,csa_tree_add_51_79_groupi_n_8450);
  not csa_tree_add_51_79_groupi_g37595(csa_tree_add_51_79_groupi_n_8437 ,csa_tree_add_51_79_groupi_n_8438);
  not csa_tree_add_51_79_groupi_g37596(csa_tree_add_51_79_groupi_n_8432 ,csa_tree_add_51_79_groupi_n_8433);
  not csa_tree_add_51_79_groupi_g37597(csa_tree_add_51_79_groupi_n_8419 ,csa_tree_add_51_79_groupi_n_8420);
  not csa_tree_add_51_79_groupi_g37598(csa_tree_add_51_79_groupi_n_8416 ,csa_tree_add_51_79_groupi_n_8417);
  not csa_tree_add_51_79_groupi_g37599(csa_tree_add_51_79_groupi_n_8413 ,csa_tree_add_51_79_groupi_n_8414);
  not csa_tree_add_51_79_groupi_g37600(csa_tree_add_51_79_groupi_n_8411 ,csa_tree_add_51_79_groupi_n_8412);
  not csa_tree_add_51_79_groupi_g37601(csa_tree_add_51_79_groupi_n_8408 ,csa_tree_add_51_79_groupi_n_8409);
  not csa_tree_add_51_79_groupi_g37602(csa_tree_add_51_79_groupi_n_8405 ,csa_tree_add_51_79_groupi_n_8406);
  not csa_tree_add_51_79_groupi_g37603(csa_tree_add_51_79_groupi_n_8403 ,csa_tree_add_51_79_groupi_n_8402);
  not csa_tree_add_51_79_groupi_g37604(csa_tree_add_51_79_groupi_n_8397 ,csa_tree_add_51_79_groupi_n_8398);
  not csa_tree_add_51_79_groupi_g37605(csa_tree_add_51_79_groupi_n_8395 ,csa_tree_add_51_79_groupi_n_8396);
  not csa_tree_add_51_79_groupi_g37606(csa_tree_add_51_79_groupi_n_8390 ,csa_tree_add_51_79_groupi_n_8391);
  not csa_tree_add_51_79_groupi_g37607(csa_tree_add_51_79_groupi_n_8385 ,csa_tree_add_51_79_groupi_n_8386);
  not csa_tree_add_51_79_groupi_g37608(csa_tree_add_51_79_groupi_n_8382 ,csa_tree_add_51_79_groupi_n_8383);
  not csa_tree_add_51_79_groupi_g37609(csa_tree_add_51_79_groupi_n_8380 ,csa_tree_add_51_79_groupi_n_8379);
  not csa_tree_add_51_79_groupi_g37610(csa_tree_add_51_79_groupi_n_8376 ,csa_tree_add_51_79_groupi_n_8377);
  not csa_tree_add_51_79_groupi_g37611(csa_tree_add_51_79_groupi_n_8374 ,csa_tree_add_51_79_groupi_n_8375);
  not csa_tree_add_51_79_groupi_g37612(csa_tree_add_51_79_groupi_n_8370 ,csa_tree_add_51_79_groupi_n_8371);
  and csa_tree_add_51_79_groupi_g37613(csa_tree_add_51_79_groupi_n_8369 ,csa_tree_add_51_79_groupi_n_8173 ,csa_tree_add_51_79_groupi_n_8170);
  or csa_tree_add_51_79_groupi_g37614(csa_tree_add_51_79_groupi_n_8368 ,csa_tree_add_51_79_groupi_n_8168 ,csa_tree_add_51_79_groupi_n_8154);
  and csa_tree_add_51_79_groupi_g37615(csa_tree_add_51_79_groupi_n_8367 ,csa_tree_add_51_79_groupi_n_8168 ,csa_tree_add_51_79_groupi_n_8154);
  or csa_tree_add_51_79_groupi_g37616(csa_tree_add_51_79_groupi_n_8366 ,csa_tree_add_51_79_groupi_n_8166 ,csa_tree_add_51_79_groupi_n_8153);
  and csa_tree_add_51_79_groupi_g37617(csa_tree_add_51_79_groupi_n_8365 ,csa_tree_add_51_79_groupi_n_8166 ,csa_tree_add_51_79_groupi_n_8153);
  or csa_tree_add_51_79_groupi_g37618(csa_tree_add_51_79_groupi_n_8364 ,csa_tree_add_51_79_groupi_n_8167 ,csa_tree_add_51_79_groupi_n_8174);
  and csa_tree_add_51_79_groupi_g37619(csa_tree_add_51_79_groupi_n_8363 ,csa_tree_add_51_79_groupi_n_8167 ,csa_tree_add_51_79_groupi_n_8174);
  or csa_tree_add_51_79_groupi_g37620(csa_tree_add_51_79_groupi_n_8362 ,csa_tree_add_51_79_groupi_n_7237 ,csa_tree_add_51_79_groupi_n_8156);
  and csa_tree_add_51_79_groupi_g37621(csa_tree_add_51_79_groupi_n_8361 ,csa_tree_add_51_79_groupi_n_7237 ,csa_tree_add_51_79_groupi_n_8156);
  or csa_tree_add_51_79_groupi_g37622(csa_tree_add_51_79_groupi_n_8360 ,csa_tree_add_51_79_groupi_n_7372 ,csa_tree_add_51_79_groupi_n_8119);
  or csa_tree_add_51_79_groupi_g37623(csa_tree_add_51_79_groupi_n_8359 ,csa_tree_add_51_79_groupi_n_8018 ,csa_tree_add_51_79_groupi_n_8163);
  nor csa_tree_add_51_79_groupi_g37624(csa_tree_add_51_79_groupi_n_8358 ,csa_tree_add_51_79_groupi_n_8019 ,csa_tree_add_51_79_groupi_n_8162);
  or csa_tree_add_51_79_groupi_g37625(csa_tree_add_51_79_groupi_n_8357 ,csa_tree_add_51_79_groupi_n_8173 ,csa_tree_add_51_79_groupi_n_8170);
  xnor csa_tree_add_51_79_groupi_g37626(csa_tree_add_51_79_groupi_n_8356 ,csa_tree_add_51_79_groupi_n_7809 ,csa_tree_add_51_79_groupi_n_7628);
  xnor csa_tree_add_51_79_groupi_g37627(csa_tree_add_51_79_groupi_n_8355 ,csa_tree_add_51_79_groupi_n_8025 ,csa_tree_add_51_79_groupi_n_7814);
  xnor csa_tree_add_51_79_groupi_g37628(csa_tree_add_51_79_groupi_n_8354 ,csa_tree_add_51_79_groupi_n_7277 ,csa_tree_add_51_79_groupi_n_7828);
  xnor csa_tree_add_51_79_groupi_g37629(csa_tree_add_51_79_groupi_n_8353 ,csa_tree_add_51_79_groupi_n_8015 ,csa_tree_add_51_79_groupi_n_7236);
  xnor csa_tree_add_51_79_groupi_g37630(csa_tree_add_51_79_groupi_n_8352 ,csa_tree_add_51_79_groupi_n_7380 ,csa_tree_add_51_79_groupi_n_7815);
  xnor csa_tree_add_51_79_groupi_g37631(csa_tree_add_51_79_groupi_n_8351 ,csa_tree_add_51_79_groupi_n_7319 ,csa_tree_add_51_79_groupi_n_8022);
  xnor csa_tree_add_51_79_groupi_g37632(csa_tree_add_51_79_groupi_n_8350 ,csa_tree_add_51_79_groupi_n_6430 ,csa_tree_add_51_79_groupi_n_7812);
  xnor csa_tree_add_51_79_groupi_g37633(csa_tree_add_51_79_groupi_n_8349 ,csa_tree_add_51_79_groupi_n_7317 ,csa_tree_add_51_79_groupi_n_7817);
  xnor csa_tree_add_51_79_groupi_g37634(csa_tree_add_51_79_groupi_n_8348 ,csa_tree_add_51_79_groupi_n_7831 ,csa_tree_add_51_79_groupi_n_7270);
  xnor csa_tree_add_51_79_groupi_g37635(csa_tree_add_51_79_groupi_n_8347 ,csa_tree_add_51_79_groupi_n_7810 ,csa_tree_add_51_79_groupi_n_7832);
  xnor csa_tree_add_51_79_groupi_g37636(csa_tree_add_51_79_groupi_n_8346 ,csa_tree_add_51_79_groupi_n_7807 ,csa_tree_add_51_79_groupi_n_8026);
  xnor csa_tree_add_51_79_groupi_g37637(csa_tree_add_51_79_groupi_n_8345 ,csa_tree_add_51_79_groupi_n_7830 ,csa_tree_add_51_79_groupi_n_7598);
  xnor csa_tree_add_51_79_groupi_g37638(csa_tree_add_51_79_groupi_n_8344 ,csa_tree_add_51_79_groupi_n_7816 ,csa_tree_add_51_79_groupi_n_6818);
  and csa_tree_add_51_79_groupi_g37639(csa_tree_add_51_79_groupi_n_8506 ,csa_tree_add_51_79_groupi_n_7767 ,csa_tree_add_51_79_groupi_n_8134);
  and csa_tree_add_51_79_groupi_g37640(csa_tree_add_51_79_groupi_n_8505 ,csa_tree_add_51_79_groupi_n_7754 ,csa_tree_add_51_79_groupi_n_8131);
  xnor csa_tree_add_51_79_groupi_g37641(csa_tree_add_51_79_groupi_n_8503 ,csa_tree_add_51_79_groupi_n_7603 ,csa_tree_add_51_79_groupi_n_7695);
  and csa_tree_add_51_79_groupi_g37642(csa_tree_add_51_79_groupi_n_8502 ,csa_tree_add_51_79_groupi_n_7752 ,csa_tree_add_51_79_groupi_n_8130);
  and csa_tree_add_51_79_groupi_g37643(csa_tree_add_51_79_groupi_n_8501 ,csa_tree_add_51_79_groupi_n_7747 ,csa_tree_add_51_79_groupi_n_8128);
  xnor csa_tree_add_51_79_groupi_g37644(csa_tree_add_51_79_groupi_n_8499 ,csa_tree_add_51_79_groupi_n_7046 ,csa_tree_add_51_79_groupi_n_7699);
  and csa_tree_add_51_79_groupi_g37645(csa_tree_add_51_79_groupi_n_8498 ,csa_tree_add_51_79_groupi_n_7739 ,csa_tree_add_51_79_groupi_n_8126);
  xnor csa_tree_add_51_79_groupi_g37646(csa_tree_add_51_79_groupi_n_8497 ,csa_tree_add_51_79_groupi_n_6890 ,csa_tree_add_51_79_groupi_n_7683);
  xnor csa_tree_add_51_79_groupi_g37647(csa_tree_add_51_79_groupi_n_8496 ,csa_tree_add_51_79_groupi_n_6963 ,csa_tree_add_51_79_groupi_n_7678);
  and csa_tree_add_51_79_groupi_g37648(csa_tree_add_51_79_groupi_n_8495 ,csa_tree_add_51_79_groupi_n_7740 ,csa_tree_add_51_79_groupi_n_8124);
  xnor csa_tree_add_51_79_groupi_g37649(csa_tree_add_51_79_groupi_n_8494 ,csa_tree_add_51_79_groupi_n_7001 ,csa_tree_add_51_79_groupi_n_7705);
  xnor csa_tree_add_51_79_groupi_g37650(csa_tree_add_51_79_groupi_n_8492 ,csa_tree_add_51_79_groupi_n_6752 ,csa_tree_add_51_79_groupi_n_28);
  xnor csa_tree_add_51_79_groupi_g37651(csa_tree_add_51_79_groupi_n_8491 ,csa_tree_add_51_79_groupi_n_6827 ,csa_tree_add_51_79_groupi_n_7643);
  and csa_tree_add_51_79_groupi_g37652(csa_tree_add_51_79_groupi_n_8490 ,csa_tree_add_51_79_groupi_n_7738 ,csa_tree_add_51_79_groupi_n_8123);
  xnor csa_tree_add_51_79_groupi_g37653(csa_tree_add_51_79_groupi_n_8489 ,csa_tree_add_51_79_groupi_n_7098 ,csa_tree_add_51_79_groupi_n_7646);
  and csa_tree_add_51_79_groupi_g37654(csa_tree_add_51_79_groupi_n_8488 ,csa_tree_add_51_79_groupi_n_7892 ,csa_tree_add_51_79_groupi_n_8120);
  xnor csa_tree_add_51_79_groupi_g37655(csa_tree_add_51_79_groupi_n_8487 ,csa_tree_add_51_79_groupi_n_7047 ,csa_tree_add_51_79_groupi_n_7664);
  xnor csa_tree_add_51_79_groupi_g37656(csa_tree_add_51_79_groupi_n_8486 ,csa_tree_add_51_79_groupi_n_7052 ,csa_tree_add_51_79_groupi_n_7711);
  xnor csa_tree_add_51_79_groupi_g37657(csa_tree_add_51_79_groupi_n_8485 ,csa_tree_add_51_79_groupi_n_7067 ,csa_tree_add_51_79_groupi_n_7714);
  xnor csa_tree_add_51_79_groupi_g37658(csa_tree_add_51_79_groupi_n_8483 ,csa_tree_add_51_79_groupi_n_6861 ,csa_tree_add_51_79_groupi_n_7710);
  xnor csa_tree_add_51_79_groupi_g37659(csa_tree_add_51_79_groupi_n_8481 ,csa_tree_add_51_79_groupi_n_6722 ,csa_tree_add_51_79_groupi_n_7698);
  and csa_tree_add_51_79_groupi_g37660(csa_tree_add_51_79_groupi_n_8480 ,csa_tree_add_51_79_groupi_n_7749 ,csa_tree_add_51_79_groupi_n_8129);
  and csa_tree_add_51_79_groupi_g37661(csa_tree_add_51_79_groupi_n_8479 ,csa_tree_add_51_79_groupi_n_7727 ,csa_tree_add_51_79_groupi_n_8136);
  or csa_tree_add_51_79_groupi_g37662(csa_tree_add_51_79_groupi_n_8477 ,csa_tree_add_51_79_groupi_n_7863 ,csa_tree_add_51_79_groupi_n_8137);
  and csa_tree_add_51_79_groupi_g37663(csa_tree_add_51_79_groupi_n_8475 ,csa_tree_add_51_79_groupi_n_7758 ,csa_tree_add_51_79_groupi_n_8132);
  and csa_tree_add_51_79_groupi_g37664(csa_tree_add_51_79_groupi_n_8474 ,csa_tree_add_51_79_groupi_n_7744 ,csa_tree_add_51_79_groupi_n_8127);
  xnor csa_tree_add_51_79_groupi_g37665(csa_tree_add_51_79_groupi_n_8473 ,csa_tree_add_51_79_groupi_n_7097 ,csa_tree_add_51_79_groupi_n_7694);
  xnor csa_tree_add_51_79_groupi_g37666(csa_tree_add_51_79_groupi_n_8472 ,csa_tree_add_51_79_groupi_n_6846 ,csa_tree_add_51_79_groupi_n_7693);
  xnor csa_tree_add_51_79_groupi_g37667(csa_tree_add_51_79_groupi_n_8470 ,csa_tree_add_51_79_groupi_n_6877 ,csa_tree_add_51_79_groupi_n_7644);
  xnor csa_tree_add_51_79_groupi_g37668(csa_tree_add_51_79_groupi_n_8468 ,csa_tree_add_51_79_groupi_n_7066 ,csa_tree_add_51_79_groupi_n_7703);
  xnor csa_tree_add_51_79_groupi_g37669(csa_tree_add_51_79_groupi_n_8466 ,csa_tree_add_51_79_groupi_n_6930 ,csa_tree_add_51_79_groupi_n_7692);
  xnor csa_tree_add_51_79_groupi_g37670(csa_tree_add_51_79_groupi_n_8465 ,csa_tree_add_51_79_groupi_n_6136 ,csa_tree_add_51_79_groupi_n_7642);
  xnor csa_tree_add_51_79_groupi_g37671(csa_tree_add_51_79_groupi_n_8464 ,csa_tree_add_51_79_groupi_n_6131 ,csa_tree_add_51_79_groupi_n_7637);
  xnor csa_tree_add_51_79_groupi_g37672(csa_tree_add_51_79_groupi_n_8462 ,csa_tree_add_51_79_groupi_n_7063 ,csa_tree_add_51_79_groupi_n_7691);
  xnor csa_tree_add_51_79_groupi_g37673(csa_tree_add_51_79_groupi_n_8461 ,csa_tree_add_51_79_groupi_n_6839 ,csa_tree_add_51_79_groupi_n_7690);
  xnor csa_tree_add_51_79_groupi_g37674(csa_tree_add_51_79_groupi_n_8460 ,csa_tree_add_51_79_groupi_n_7074 ,csa_tree_add_51_79_groupi_n_7704);
  xnor csa_tree_add_51_79_groupi_g37675(csa_tree_add_51_79_groupi_n_8459 ,csa_tree_add_51_79_groupi_n_6745 ,csa_tree_add_51_79_groupi_n_7660);
  xnor csa_tree_add_51_79_groupi_g37676(csa_tree_add_51_79_groupi_n_8456 ,csa_tree_add_51_79_groupi_n_6836 ,csa_tree_add_51_79_groupi_n_7689);
  xnor csa_tree_add_51_79_groupi_g37677(csa_tree_add_51_79_groupi_n_8454 ,csa_tree_add_51_79_groupi_n_6939 ,csa_tree_add_51_79_groupi_n_7688);
  and csa_tree_add_51_79_groupi_g37678(csa_tree_add_51_79_groupi_n_8453 ,csa_tree_add_51_79_groupi_n_7772 ,csa_tree_add_51_79_groupi_n_8135);
  xnor csa_tree_add_51_79_groupi_g37679(csa_tree_add_51_79_groupi_n_8452 ,csa_tree_add_51_79_groupi_n_6736 ,csa_tree_add_51_79_groupi_n_27);
  xnor csa_tree_add_51_79_groupi_g37680(csa_tree_add_51_79_groupi_n_8450 ,csa_tree_add_51_79_groupi_n_7040 ,csa_tree_add_51_79_groupi_n_7686);
  xnor csa_tree_add_51_79_groupi_g37681(csa_tree_add_51_79_groupi_n_8449 ,csa_tree_add_51_79_groupi_n_6831 ,csa_tree_add_51_79_groupi_n_7685);
  xnor csa_tree_add_51_79_groupi_g37682(csa_tree_add_51_79_groupi_n_8448 ,csa_tree_add_51_79_groupi_n_7069 ,csa_tree_add_51_79_groupi_n_7684);
  xnor csa_tree_add_51_79_groupi_g37683(csa_tree_add_51_79_groupi_n_8447 ,csa_tree_add_51_79_groupi_n_6934 ,csa_tree_add_51_79_groupi_n_7682);
  xnor csa_tree_add_51_79_groupi_g37684(csa_tree_add_51_79_groupi_n_8446 ,csa_tree_add_51_79_groupi_n_6128 ,csa_tree_add_51_79_groupi_n_7661);
  xnor csa_tree_add_51_79_groupi_g37685(csa_tree_add_51_79_groupi_n_8445 ,csa_tree_add_51_79_groupi_n_6895 ,csa_tree_add_51_79_groupi_n_7681);
  xnor csa_tree_add_51_79_groupi_g37686(csa_tree_add_51_79_groupi_n_8444 ,csa_tree_add_51_79_groupi_n_6828 ,csa_tree_add_51_79_groupi_n_7680);
  xnor csa_tree_add_51_79_groupi_g37687(csa_tree_add_51_79_groupi_n_8443 ,csa_tree_add_51_79_groupi_n_7071 ,csa_tree_add_51_79_groupi_n_7679);
  xnor csa_tree_add_51_79_groupi_g37688(csa_tree_add_51_79_groupi_n_8442 ,csa_tree_add_51_79_groupi_n_5851 ,csa_tree_add_51_79_groupi_n_7687);
  xnor csa_tree_add_51_79_groupi_g37689(csa_tree_add_51_79_groupi_n_8441 ,csa_tree_add_51_79_groupi_n_7105 ,csa_tree_add_51_79_groupi_n_7677);
  xnor csa_tree_add_51_79_groupi_g37690(csa_tree_add_51_79_groupi_n_8440 ,csa_tree_add_51_79_groupi_n_7096 ,csa_tree_add_51_79_groupi_n_7675);
  xnor csa_tree_add_51_79_groupi_g37691(csa_tree_add_51_79_groupi_n_8439 ,csa_tree_add_51_79_groupi_n_7202 ,csa_tree_add_51_79_groupi_n_7674);
  xnor csa_tree_add_51_79_groupi_g37692(csa_tree_add_51_79_groupi_n_8438 ,csa_tree_add_51_79_groupi_n_6134 ,csa_tree_add_51_79_groupi_n_7717);
  xnor csa_tree_add_51_79_groupi_g37693(csa_tree_add_51_79_groupi_n_8436 ,csa_tree_add_51_79_groupi_n_6969 ,csa_tree_add_51_79_groupi_n_7672);
  xnor csa_tree_add_51_79_groupi_g37694(csa_tree_add_51_79_groupi_n_8435 ,csa_tree_add_51_79_groupi_n_6907 ,csa_tree_add_51_79_groupi_n_7668);
  xnor csa_tree_add_51_79_groupi_g37695(csa_tree_add_51_79_groupi_n_8434 ,csa_tree_add_51_79_groupi_n_6905 ,csa_tree_add_51_79_groupi_n_7676);
  xnor csa_tree_add_51_79_groupi_g37696(csa_tree_add_51_79_groupi_n_8433 ,csa_tree_add_51_79_groupi_n_7025 ,csa_tree_add_51_79_groupi_n_7669);
  xnor csa_tree_add_51_79_groupi_g37697(csa_tree_add_51_79_groupi_n_8431 ,csa_tree_add_51_79_groupi_n_6883 ,csa_tree_add_51_79_groupi_n_7671);
  xnor csa_tree_add_51_79_groupi_g37698(csa_tree_add_51_79_groupi_n_8430 ,csa_tree_add_51_79_groupi_n_6917 ,csa_tree_add_51_79_groupi_n_7670);
  xnor csa_tree_add_51_79_groupi_g37699(csa_tree_add_51_79_groupi_n_8429 ,csa_tree_add_51_79_groupi_n_6863 ,csa_tree_add_51_79_groupi_n_7667);
  xnor csa_tree_add_51_79_groupi_g37700(csa_tree_add_51_79_groupi_n_8428 ,csa_tree_add_51_79_groupi_n_6910 ,csa_tree_add_51_79_groupi_n_7666);
  xnor csa_tree_add_51_79_groupi_g37701(csa_tree_add_51_79_groupi_n_8427 ,csa_tree_add_51_79_groupi_n_6894 ,csa_tree_add_51_79_groupi_n_7654);
  xnor csa_tree_add_51_79_groupi_g37702(csa_tree_add_51_79_groupi_n_8426 ,csa_tree_add_51_79_groupi_n_6931 ,csa_tree_add_51_79_groupi_n_7653);
  xnor csa_tree_add_51_79_groupi_g37703(csa_tree_add_51_79_groupi_n_8425 ,csa_tree_add_51_79_groupi_n_7050 ,csa_tree_add_51_79_groupi_n_7647);
  xnor csa_tree_add_51_79_groupi_g37704(csa_tree_add_51_79_groupi_n_8424 ,csa_tree_add_51_79_groupi_n_7109 ,csa_tree_add_51_79_groupi_n_7641);
  xnor csa_tree_add_51_79_groupi_g37705(csa_tree_add_51_79_groupi_n_8423 ,csa_tree_add_51_79_groupi_n_6986 ,csa_tree_add_51_79_groupi_n_7639);
  xnor csa_tree_add_51_79_groupi_g37706(csa_tree_add_51_79_groupi_n_8422 ,csa_tree_add_51_79_groupi_n_7039 ,csa_tree_add_51_79_groupi_n_7716);
  xnor csa_tree_add_51_79_groupi_g37707(csa_tree_add_51_79_groupi_n_8421 ,csa_tree_add_51_79_groupi_n_6902 ,csa_tree_add_51_79_groupi_n_7713);
  xnor csa_tree_add_51_79_groupi_g37708(csa_tree_add_51_79_groupi_n_8420 ,csa_tree_add_51_79_groupi_n_7008 ,csa_tree_add_51_79_groupi_n_7707);
  xnor csa_tree_add_51_79_groupi_g37709(csa_tree_add_51_79_groupi_n_8418 ,csa_tree_add_51_79_groupi_n_6431 ,csa_tree_add_51_79_groupi_n_7658);
  xnor csa_tree_add_51_79_groupi_g37710(csa_tree_add_51_79_groupi_n_8417 ,csa_tree_add_51_79_groupi_n_7079 ,csa_tree_add_51_79_groupi_n_7721);
  xnor csa_tree_add_51_79_groupi_g37711(csa_tree_add_51_79_groupi_n_8415 ,csa_tree_add_51_79_groupi_n_7617 ,csa_tree_add_51_79_groupi_n_7665);
  xnor csa_tree_add_51_79_groupi_g37713(csa_tree_add_51_79_groupi_n_8414 ,csa_tree_add_51_79_groupi_n_7164 ,csa_tree_add_51_79_groupi_n_7673);
  xnor csa_tree_add_51_79_groupi_g37714(csa_tree_add_51_79_groupi_n_8412 ,csa_tree_add_51_79_groupi_n_6862 ,csa_tree_add_51_79_groupi_n_7656);
  xnor csa_tree_add_51_79_groupi_g37715(csa_tree_add_51_79_groupi_n_8410 ,csa_tree_add_51_79_groupi_n_6819 ,csa_tree_add_51_79_groupi_n_7655);
  xnor csa_tree_add_51_79_groupi_g37716(csa_tree_add_51_79_groupi_n_8409 ,csa_tree_add_51_79_groupi_n_7087 ,csa_tree_add_51_79_groupi_n_7652);
  xnor csa_tree_add_51_79_groupi_g37717(csa_tree_add_51_79_groupi_n_8407 ,csa_tree_add_51_79_groupi_n_6875 ,csa_tree_add_51_79_groupi_n_7651);
  xnor csa_tree_add_51_79_groupi_g37718(csa_tree_add_51_79_groupi_n_8406 ,csa_tree_add_51_79_groupi_n_6899 ,csa_tree_add_51_79_groupi_n_7650);
  xnor csa_tree_add_51_79_groupi_g37719(csa_tree_add_51_79_groupi_n_8404 ,csa_tree_add_51_79_groupi_n_6993 ,csa_tree_add_51_79_groupi_n_7648);
  xnor csa_tree_add_51_79_groupi_g37720(csa_tree_add_51_79_groupi_n_8402 ,csa_tree_add_51_79_groupi_n_7085 ,csa_tree_add_51_79_groupi_n_7697);
  xnor csa_tree_add_51_79_groupi_g37721(csa_tree_add_51_79_groupi_n_8401 ,csa_tree_add_51_79_groupi_n_6872 ,csa_tree_add_51_79_groupi_n_7645);
  and csa_tree_add_51_79_groupi_g37722(csa_tree_add_51_79_groupi_n_8400 ,csa_tree_add_51_79_groupi_n_7742 ,csa_tree_add_51_79_groupi_n_8125);
  xnor csa_tree_add_51_79_groupi_g37723(csa_tree_add_51_79_groupi_n_8399 ,csa_tree_add_51_79_groupi_n_6965 ,csa_tree_add_51_79_groupi_n_7640);
  xnor csa_tree_add_51_79_groupi_g37724(csa_tree_add_51_79_groupi_n_8398 ,csa_tree_add_51_79_groupi_n_7032 ,csa_tree_add_51_79_groupi_n_7638);
  xnor csa_tree_add_51_79_groupi_g37725(csa_tree_add_51_79_groupi_n_8396 ,csa_tree_add_51_79_groupi_n_7064 ,csa_tree_add_51_79_groupi_n_7636);
  xnor csa_tree_add_51_79_groupi_g37726(csa_tree_add_51_79_groupi_n_8394 ,csa_tree_add_51_79_groupi_n_7112 ,csa_tree_add_51_79_groupi_n_7715);
  xnor csa_tree_add_51_79_groupi_g37727(csa_tree_add_51_79_groupi_n_8393 ,csa_tree_add_51_79_groupi_n_7014 ,csa_tree_add_51_79_groupi_n_7657);
  xnor csa_tree_add_51_79_groupi_g37728(csa_tree_add_51_79_groupi_n_8392 ,csa_tree_add_51_79_groupi_n_7094 ,csa_tree_add_51_79_groupi_n_7659);
  xnor csa_tree_add_51_79_groupi_g37729(csa_tree_add_51_79_groupi_n_8391 ,csa_tree_add_51_79_groupi_n_6897 ,csa_tree_add_51_79_groupi_n_7708);
  xnor csa_tree_add_51_79_groupi_g37730(csa_tree_add_51_79_groupi_n_8389 ,csa_tree_add_51_79_groupi_n_6990 ,csa_tree_add_51_79_groupi_n_7662);
  xnor csa_tree_add_51_79_groupi_g37731(csa_tree_add_51_79_groupi_n_8388 ,csa_tree_add_51_79_groupi_n_7168 ,csa_tree_add_51_79_groupi_n_7702);
  xnor csa_tree_add_51_79_groupi_g37732(csa_tree_add_51_79_groupi_n_8387 ,csa_tree_add_51_79_groupi_n_7113 ,csa_tree_add_51_79_groupi_n_7663);
  xnor csa_tree_add_51_79_groupi_g37733(csa_tree_add_51_79_groupi_n_8386 ,csa_tree_add_51_79_groupi_n_7089 ,csa_tree_add_51_79_groupi_n_7696);
  xnor csa_tree_add_51_79_groupi_g37734(csa_tree_add_51_79_groupi_n_8384 ,csa_tree_add_51_79_groupi_n_7073 ,csa_tree_add_51_79_groupi_n_7701);
  xnor csa_tree_add_51_79_groupi_g37735(csa_tree_add_51_79_groupi_n_8383 ,csa_tree_add_51_79_groupi_n_7624 ,csa_tree_add_51_79_groupi_n_7709);
  xnor csa_tree_add_51_79_groupi_g37736(csa_tree_add_51_79_groupi_n_8381 ,csa_tree_add_51_79_groupi_n_6976 ,csa_tree_add_51_79_groupi_n_7706);
  xnor csa_tree_add_51_79_groupi_g37737(csa_tree_add_51_79_groupi_n_8379 ,csa_tree_add_51_79_groupi_n_7065 ,csa_tree_add_51_79_groupi_n_7700);
  and csa_tree_add_51_79_groupi_g37738(csa_tree_add_51_79_groupi_n_8378 ,csa_tree_add_51_79_groupi_n_7759 ,csa_tree_add_51_79_groupi_n_8133);
  xnor csa_tree_add_51_79_groupi_g37739(csa_tree_add_51_79_groupi_n_8377 ,csa_tree_add_51_79_groupi_n_7030 ,csa_tree_add_51_79_groupi_n_7649);
  xnor csa_tree_add_51_79_groupi_g37740(csa_tree_add_51_79_groupi_n_8375 ,csa_tree_add_51_79_groupi_n_6991 ,csa_tree_add_51_79_groupi_n_7718);
  xnor csa_tree_add_51_79_groupi_g37741(csa_tree_add_51_79_groupi_n_8373 ,csa_tree_add_51_79_groupi_n_6878 ,csa_tree_add_51_79_groupi_n_7712);
  xnor csa_tree_add_51_79_groupi_g37742(csa_tree_add_51_79_groupi_n_8372 ,csa_tree_add_51_79_groupi_n_6858 ,csa_tree_add_51_79_groupi_n_7719);
  xnor csa_tree_add_51_79_groupi_g37743(csa_tree_add_51_79_groupi_n_8371 ,csa_tree_add_51_79_groupi_n_7027 ,csa_tree_add_51_79_groupi_n_7720);
  not csa_tree_add_51_79_groupi_g37744(csa_tree_add_51_79_groupi_n_8329 ,csa_tree_add_51_79_groupi_n_8328);
  not csa_tree_add_51_79_groupi_g37745(csa_tree_add_51_79_groupi_n_8306 ,csa_tree_add_51_79_groupi_n_8307);
  not csa_tree_add_51_79_groupi_g37746(csa_tree_add_51_79_groupi_n_8303 ,csa_tree_add_51_79_groupi_n_8304);
  not csa_tree_add_51_79_groupi_g37747(csa_tree_add_51_79_groupi_n_8294 ,csa_tree_add_51_79_groupi_n_8295);
  not csa_tree_add_51_79_groupi_g37748(csa_tree_add_51_79_groupi_n_8281 ,csa_tree_add_51_79_groupi_n_8282);
  not csa_tree_add_51_79_groupi_g37749(csa_tree_add_51_79_groupi_n_8275 ,csa_tree_add_51_79_groupi_n_8274);
  not csa_tree_add_51_79_groupi_g37750(csa_tree_add_51_79_groupi_n_8272 ,csa_tree_add_51_79_groupi_n_8271);
  not csa_tree_add_51_79_groupi_g37751(csa_tree_add_51_79_groupi_n_8266 ,csa_tree_add_51_79_groupi_n_8267);
  or csa_tree_add_51_79_groupi_g37752(csa_tree_add_51_79_groupi_n_8264 ,csa_tree_add_51_79_groupi_n_7342 ,csa_tree_add_51_79_groupi_n_7918);
  or csa_tree_add_51_79_groupi_g37753(csa_tree_add_51_79_groupi_n_8263 ,csa_tree_add_51_79_groupi_n_7318 ,csa_tree_add_51_79_groupi_n_7795);
  or csa_tree_add_51_79_groupi_g37754(csa_tree_add_51_79_groupi_n_8262 ,csa_tree_add_51_79_groupi_n_7341 ,csa_tree_add_51_79_groupi_n_7769);
  or csa_tree_add_51_79_groupi_g37755(csa_tree_add_51_79_groupi_n_8261 ,csa_tree_add_51_79_groupi_n_7360 ,csa_tree_add_51_79_groupi_n_7762);
  or csa_tree_add_51_79_groupi_g37756(csa_tree_add_51_79_groupi_n_8260 ,csa_tree_add_51_79_groupi_n_7388 ,csa_tree_add_51_79_groupi_n_7722);
  or csa_tree_add_51_79_groupi_g37757(csa_tree_add_51_79_groupi_n_8259 ,csa_tree_add_51_79_groupi_n_7361 ,csa_tree_add_51_79_groupi_n_7974);
  or csa_tree_add_51_79_groupi_g37758(csa_tree_add_51_79_groupi_n_8258 ,csa_tree_add_51_79_groupi_n_7362 ,csa_tree_add_51_79_groupi_n_7933);
  and csa_tree_add_51_79_groupi_g37759(csa_tree_add_51_79_groupi_n_8257 ,csa_tree_add_51_79_groupi_n_8023 ,csa_tree_add_51_79_groupi_n_7820);
  or csa_tree_add_51_79_groupi_g37760(csa_tree_add_51_79_groupi_n_8256 ,csa_tree_add_51_79_groupi_n_7339 ,csa_tree_add_51_79_groupi_n_8003);
  or csa_tree_add_51_79_groupi_g37761(csa_tree_add_51_79_groupi_n_8255 ,csa_tree_add_51_79_groupi_n_7236 ,csa_tree_add_51_79_groupi_n_8015);
  or csa_tree_add_51_79_groupi_g37762(csa_tree_add_51_79_groupi_n_8254 ,csa_tree_add_51_79_groupi_n_8023 ,csa_tree_add_51_79_groupi_n_7820);
  and csa_tree_add_51_79_groupi_g37763(csa_tree_add_51_79_groupi_n_8253 ,csa_tree_add_51_79_groupi_n_7343 ,csa_tree_add_51_79_groupi_n_7837);
  and csa_tree_add_51_79_groupi_g37764(csa_tree_add_51_79_groupi_n_8252 ,csa_tree_add_51_79_groupi_n_6818 ,csa_tree_add_51_79_groupi_n_7816);
  and csa_tree_add_51_79_groupi_g37765(csa_tree_add_51_79_groupi_n_8251 ,csa_tree_add_51_79_groupi_n_7236 ,csa_tree_add_51_79_groupi_n_8015);
  or csa_tree_add_51_79_groupi_g37766(csa_tree_add_51_79_groupi_n_8250 ,csa_tree_add_51_79_groupi_n_6818 ,csa_tree_add_51_79_groupi_n_7816);
  and csa_tree_add_51_79_groupi_g37767(csa_tree_add_51_79_groupi_n_8249 ,csa_tree_add_51_79_groupi_n_7330 ,csa_tree_add_51_79_groupi_n_7835);
  and csa_tree_add_51_79_groupi_g37768(csa_tree_add_51_79_groupi_n_8248 ,csa_tree_add_51_79_groupi_n_7630 ,csa_tree_add_51_79_groupi_n_7997);
  or csa_tree_add_51_79_groupi_g37769(csa_tree_add_51_79_groupi_n_8247 ,csa_tree_add_51_79_groupi_n_7338 ,csa_tree_add_51_79_groupi_n_7994);
  or csa_tree_add_51_79_groupi_g37770(csa_tree_add_51_79_groupi_n_8246 ,csa_tree_add_51_79_groupi_n_7320 ,csa_tree_add_51_79_groupi_n_7839);
  and csa_tree_add_51_79_groupi_g37771(csa_tree_add_51_79_groupi_n_8245 ,csa_tree_add_51_79_groupi_n_7629 ,csa_tree_add_51_79_groupi_n_7990);
  or csa_tree_add_51_79_groupi_g37772(csa_tree_add_51_79_groupi_n_8244 ,csa_tree_add_51_79_groupi_n_7828 ,csa_tree_add_51_79_groupi_n_7988);
  or csa_tree_add_51_79_groupi_g37773(csa_tree_add_51_79_groupi_n_8243 ,csa_tree_add_51_79_groupi_n_7321 ,csa_tree_add_51_79_groupi_n_7842);
  or csa_tree_add_51_79_groupi_g37774(csa_tree_add_51_79_groupi_n_8242 ,csa_tree_add_51_79_groupi_n_7337 ,csa_tree_add_51_79_groupi_n_7985);
  or csa_tree_add_51_79_groupi_g37775(csa_tree_add_51_79_groupi_n_8241 ,csa_tree_add_51_79_groupi_n_7386 ,csa_tree_add_51_79_groupi_n_7983);
  or csa_tree_add_51_79_groupi_g37776(csa_tree_add_51_79_groupi_n_8240 ,csa_tree_add_51_79_groupi_n_8021 ,csa_tree_add_51_79_groupi_n_7821);
  or csa_tree_add_51_79_groupi_g37777(csa_tree_add_51_79_groupi_n_8239 ,csa_tree_add_51_79_groupi_n_7385 ,csa_tree_add_51_79_groupi_n_7981);
  or csa_tree_add_51_79_groupi_g37778(csa_tree_add_51_79_groupi_n_8238 ,csa_tree_add_51_79_groupi_n_7357 ,csa_tree_add_51_79_groupi_n_7978);
  or csa_tree_add_51_79_groupi_g37779(csa_tree_add_51_79_groupi_n_8237 ,csa_tree_add_51_79_groupi_n_8025 ,csa_tree_add_51_79_groupi_n_7813);
  nor csa_tree_add_51_79_groupi_g37780(csa_tree_add_51_79_groupi_n_8236 ,csa_tree_add_51_79_groupi_n_8024 ,csa_tree_add_51_79_groupi_n_7814);
  and csa_tree_add_51_79_groupi_g37781(csa_tree_add_51_79_groupi_n_8235 ,csa_tree_add_51_79_groupi_n_8026 ,csa_tree_add_51_79_groupi_n_7807);
  or csa_tree_add_51_79_groupi_g37782(csa_tree_add_51_79_groupi_n_8234 ,csa_tree_add_51_79_groupi_n_8026 ,csa_tree_add_51_79_groupi_n_7807);
  or csa_tree_add_51_79_groupi_g37783(csa_tree_add_51_79_groupi_n_8233 ,csa_tree_add_51_79_groupi_n_7368 ,csa_tree_add_51_79_groupi_n_7869);
  or csa_tree_add_51_79_groupi_g37784(csa_tree_add_51_79_groupi_n_8232 ,csa_tree_add_51_79_groupi_n_7827 ,csa_tree_add_51_79_groupi_n_7849);
  and csa_tree_add_51_79_groupi_g37785(csa_tree_add_51_79_groupi_n_8231 ,csa_tree_add_51_79_groupi_n_7626 ,csa_tree_add_51_79_groupi_n_7967);
  or csa_tree_add_51_79_groupi_g37786(csa_tree_add_51_79_groupi_n_8230 ,csa_tree_add_51_79_groupi_n_7322 ,csa_tree_add_51_79_groupi_n_7783);
  or csa_tree_add_51_79_groupi_g37787(csa_tree_add_51_79_groupi_n_8229 ,csa_tree_add_51_79_groupi_n_6918 ,csa_tree_add_51_79_groupi_n_7860);
  or csa_tree_add_51_79_groupi_g37788(csa_tree_add_51_79_groupi_n_8228 ,csa_tree_add_51_79_groupi_n_7107 ,csa_tree_add_51_79_groupi_n_7962);
  or csa_tree_add_51_79_groupi_g37789(csa_tree_add_51_79_groupi_n_8227 ,csa_tree_add_51_79_groupi_n_7336 ,csa_tree_add_51_79_groupi_n_7963);
  or csa_tree_add_51_79_groupi_g37790(csa_tree_add_51_79_groupi_n_8226 ,csa_tree_add_51_79_groupi_n_7335 ,csa_tree_add_51_79_groupi_n_7781);
  or csa_tree_add_51_79_groupi_g37791(csa_tree_add_51_79_groupi_n_8225 ,csa_tree_add_51_79_groupi_n_7334 ,csa_tree_add_51_79_groupi_n_7764);
  or csa_tree_add_51_79_groupi_g37792(csa_tree_add_51_79_groupi_n_8224 ,csa_tree_add_51_79_groupi_n_7333 ,csa_tree_add_51_79_groupi_n_7958);
  or csa_tree_add_51_79_groupi_g37793(csa_tree_add_51_79_groupi_n_8223 ,csa_tree_add_51_79_groupi_n_7383 ,csa_tree_add_51_79_groupi_n_7956);
  or csa_tree_add_51_79_groupi_g37794(csa_tree_add_51_79_groupi_n_8222 ,csa_tree_add_51_79_groupi_n_6906 ,csa_tree_add_51_79_groupi_n_7725);
  nor csa_tree_add_51_79_groupi_g37795(csa_tree_add_51_79_groupi_n_8221 ,csa_tree_add_51_79_groupi_n_7625 ,csa_tree_add_51_79_groupi_n_7954);
  or csa_tree_add_51_79_groupi_g37796(csa_tree_add_51_79_groupi_n_8220 ,csa_tree_add_51_79_groupi_n_7332 ,csa_tree_add_51_79_groupi_n_29);
  and csa_tree_add_51_79_groupi_g37797(csa_tree_add_51_79_groupi_n_8219 ,csa_tree_add_51_79_groupi_n_7344 ,csa_tree_add_51_79_groupi_n_7864);
  nor csa_tree_add_51_79_groupi_g37798(csa_tree_add_51_79_groupi_n_8218 ,csa_tree_add_51_79_groupi_n_7623 ,csa_tree_add_51_79_groupi_n_7945);
  or csa_tree_add_51_79_groupi_g37799(csa_tree_add_51_79_groupi_n_8217 ,csa_tree_add_51_79_groupi_n_7382 ,csa_tree_add_51_79_groupi_n_7944);
  or csa_tree_add_51_79_groupi_g37800(csa_tree_add_51_79_groupi_n_8216 ,csa_tree_add_51_79_groupi_n_7331 ,csa_tree_add_51_79_groupi_n_7761);
  or csa_tree_add_51_79_groupi_g37801(csa_tree_add_51_79_groupi_n_8215 ,csa_tree_add_51_79_groupi_n_7622 ,csa_tree_add_51_79_groupi_n_7939);
  and csa_tree_add_51_79_groupi_g37802(csa_tree_add_51_79_groupi_n_8214 ,csa_tree_add_51_79_groupi_n_7633 ,csa_tree_add_51_79_groupi_n_7941);
  or csa_tree_add_51_79_groupi_g37803(csa_tree_add_51_79_groupi_n_8213 ,csa_tree_add_51_79_groupi_n_7809 ,csa_tree_add_51_79_groupi_n_7169);
  or csa_tree_add_51_79_groupi_g37804(csa_tree_add_51_79_groupi_n_8212 ,csa_tree_add_51_79_groupi_n_7329 ,csa_tree_add_51_79_groupi_n_7867);
  or csa_tree_add_51_79_groupi_g37805(csa_tree_add_51_79_groupi_n_8211 ,csa_tree_add_51_79_groupi_n_7777 ,csa_tree_add_51_79_groupi_n_8027);
  nor csa_tree_add_51_79_groupi_g37806(csa_tree_add_51_79_groupi_n_8210 ,csa_tree_add_51_79_groupi_n_7808 ,csa_tree_add_51_79_groupi_n_7170);
  or csa_tree_add_51_79_groupi_g37807(csa_tree_add_51_79_groupi_n_8209 ,csa_tree_add_51_79_groupi_n_7620 ,csa_tree_add_51_79_groupi_n_7871);
  or csa_tree_add_51_79_groupi_g37808(csa_tree_add_51_79_groupi_n_8208 ,csa_tree_add_51_79_groupi_n_7354 ,csa_tree_add_51_79_groupi_n_7874);
  or csa_tree_add_51_79_groupi_g37809(csa_tree_add_51_79_groupi_n_8207 ,csa_tree_add_51_79_groupi_n_7632 ,csa_tree_add_51_79_groupi_n_7949);
  or csa_tree_add_51_79_groupi_g37810(csa_tree_add_51_79_groupi_n_8206 ,csa_tree_add_51_79_groupi_n_6900 ,csa_tree_add_51_79_groupi_n_7876);
  or csa_tree_add_51_79_groupi_g37811(csa_tree_add_51_79_groupi_n_8205 ,csa_tree_add_51_79_groupi_n_7323 ,csa_tree_add_51_79_groupi_n_7750);
  or csa_tree_add_51_79_groupi_g37812(csa_tree_add_51_79_groupi_n_8204 ,csa_tree_add_51_79_groupi_n_7325 ,csa_tree_add_51_79_groupi_n_7881);
  or csa_tree_add_51_79_groupi_g37813(csa_tree_add_51_79_groupi_n_8203 ,csa_tree_add_51_79_groupi_n_7381 ,csa_tree_add_51_79_groupi_n_7930);
  or csa_tree_add_51_79_groupi_g37814(csa_tree_add_51_79_groupi_n_8202 ,csa_tree_add_51_79_groupi_n_7815 ,csa_tree_add_51_79_groupi_n_7204);
  or csa_tree_add_51_79_groupi_g37815(csa_tree_add_51_79_groupi_n_8201 ,csa_tree_add_51_79_groupi_n_7346 ,csa_tree_add_51_79_groupi_n_7883);
  and csa_tree_add_51_79_groupi_g37816(csa_tree_add_51_79_groupi_n_8200 ,csa_tree_add_51_79_groupi_n_7815 ,csa_tree_add_51_79_groupi_n_7204);
  or csa_tree_add_51_79_groupi_g37817(csa_tree_add_51_79_groupi_n_8199 ,csa_tree_add_51_79_groupi_n_7090 ,csa_tree_add_51_79_groupi_n_7926);
  or csa_tree_add_51_79_groupi_g37818(csa_tree_add_51_79_groupi_n_8198 ,csa_tree_add_51_79_groupi_n_7378 ,csa_tree_add_51_79_groupi_n_7922);
  or csa_tree_add_51_79_groupi_g37819(csa_tree_add_51_79_groupi_n_8197 ,csa_tree_add_51_79_groupi_n_7634 ,csa_tree_add_51_79_groupi_n_7919);
  or csa_tree_add_51_79_groupi_g37820(csa_tree_add_51_79_groupi_n_8196 ,csa_tree_add_51_79_groupi_n_7377 ,csa_tree_add_51_79_groupi_n_7920);
  and csa_tree_add_51_79_groupi_g37821(csa_tree_add_51_79_groupi_n_8195 ,csa_tree_add_51_79_groupi_n_7347 ,csa_tree_add_51_79_groupi_n_7885);
  and csa_tree_add_51_79_groupi_g37822(csa_tree_add_51_79_groupi_n_8194 ,csa_tree_add_51_79_groupi_n_7618 ,csa_tree_add_51_79_groupi_n_7916);
  and csa_tree_add_51_79_groupi_g37823(csa_tree_add_51_79_groupi_n_8193 ,csa_tree_add_51_79_groupi_n_7635 ,csa_tree_add_51_79_groupi_n_7913);
  and csa_tree_add_51_79_groupi_g37824(csa_tree_add_51_79_groupi_n_8192 ,csa_tree_add_51_79_groupi_n_7359 ,csa_tree_add_51_79_groupi_n_7888);
  or csa_tree_add_51_79_groupi_g37825(csa_tree_add_51_79_groupi_n_8191 ,csa_tree_add_51_79_groupi_n_7328 ,csa_tree_add_51_79_groupi_n_7911);
  or csa_tree_add_51_79_groupi_g37826(csa_tree_add_51_79_groupi_n_8190 ,csa_tree_add_51_79_groupi_n_7326 ,csa_tree_add_51_79_groupi_n_7890);
  and csa_tree_add_51_79_groupi_g37827(csa_tree_add_51_79_groupi_n_8189 ,csa_tree_add_51_79_groupi_n_7348 ,csa_tree_add_51_79_groupi_n_7891);
  or csa_tree_add_51_79_groupi_g37828(csa_tree_add_51_79_groupi_n_8188 ,csa_tree_add_51_79_groupi_n_7324 ,csa_tree_add_51_79_groupi_n_7868);
  or csa_tree_add_51_79_groupi_g37829(csa_tree_add_51_79_groupi_n_8187 ,csa_tree_add_51_79_groupi_n_7327 ,csa_tree_add_51_79_groupi_n_7755);
  or csa_tree_add_51_79_groupi_g37830(csa_tree_add_51_79_groupi_n_8186 ,csa_tree_add_51_79_groupi_n_7376 ,csa_tree_add_51_79_groupi_n_7904);
  or csa_tree_add_51_79_groupi_g37831(csa_tree_add_51_79_groupi_n_8343 ,csa_tree_add_51_79_groupi_n_6953 ,csa_tree_add_51_79_groupi_n_7893);
  and csa_tree_add_51_79_groupi_g37832(csa_tree_add_51_79_groupi_n_8342 ,csa_tree_add_51_79_groupi_n_7480 ,csa_tree_add_51_79_groupi_n_7898);
  and csa_tree_add_51_79_groupi_g37833(csa_tree_add_51_79_groupi_n_8341 ,csa_tree_add_51_79_groupi_n_7479 ,csa_tree_add_51_79_groupi_n_7900);
  and csa_tree_add_51_79_groupi_g37834(csa_tree_add_51_79_groupi_n_8340 ,csa_tree_add_51_79_groupi_n_7478 ,csa_tree_add_51_79_groupi_n_7897);
  and csa_tree_add_51_79_groupi_g37835(csa_tree_add_51_79_groupi_n_8339 ,csa_tree_add_51_79_groupi_n_7501 ,csa_tree_add_51_79_groupi_n_7848);
  and csa_tree_add_51_79_groupi_g37836(csa_tree_add_51_79_groupi_n_8338 ,csa_tree_add_51_79_groupi_n_7498 ,csa_tree_add_51_79_groupi_n_7894);
  and csa_tree_add_51_79_groupi_g37837(csa_tree_add_51_79_groupi_n_8337 ,csa_tree_add_51_79_groupi_n_7473 ,csa_tree_add_51_79_groupi_n_7879);
  and csa_tree_add_51_79_groupi_g37838(csa_tree_add_51_79_groupi_n_8336 ,csa_tree_add_51_79_groupi_n_7525 ,csa_tree_add_51_79_groupi_n_7908);
  and csa_tree_add_51_79_groupi_g37839(csa_tree_add_51_79_groupi_n_8335 ,csa_tree_add_51_79_groupi_n_7414 ,csa_tree_add_51_79_groupi_n_7843);
  and csa_tree_add_51_79_groupi_g37840(csa_tree_add_51_79_groupi_n_8334 ,csa_tree_add_51_79_groupi_n_7500 ,csa_tree_add_51_79_groupi_n_7914);
  and csa_tree_add_51_79_groupi_g37841(csa_tree_add_51_79_groupi_n_8333 ,csa_tree_add_51_79_groupi_n_7509 ,csa_tree_add_51_79_groupi_n_7925);
  and csa_tree_add_51_79_groupi_g37842(csa_tree_add_51_79_groupi_n_8332 ,csa_tree_add_51_79_groupi_n_7513 ,csa_tree_add_51_79_groupi_n_7932);
  and csa_tree_add_51_79_groupi_g37843(csa_tree_add_51_79_groupi_n_8331 ,csa_tree_add_51_79_groupi_n_7515 ,csa_tree_add_51_79_groupi_n_7936);
  or csa_tree_add_51_79_groupi_g37844(csa_tree_add_51_79_groupi_n_8330 ,csa_tree_add_51_79_groupi_n_7505 ,csa_tree_add_51_79_groupi_n_7846);
  and csa_tree_add_51_79_groupi_g37845(csa_tree_add_51_79_groupi_n_8328 ,csa_tree_add_51_79_groupi_n_6760 ,csa_tree_add_51_79_groupi_n_8029);
  and csa_tree_add_51_79_groupi_g37846(csa_tree_add_51_79_groupi_n_8327 ,csa_tree_add_51_79_groupi_n_7531 ,csa_tree_add_51_79_groupi_n_7964);
  and csa_tree_add_51_79_groupi_g37847(csa_tree_add_51_79_groupi_n_8326 ,csa_tree_add_51_79_groupi_n_7456 ,csa_tree_add_51_79_groupi_n_7854);
  and csa_tree_add_51_79_groupi_g37848(csa_tree_add_51_79_groupi_n_8325 ,csa_tree_add_51_79_groupi_n_7538 ,csa_tree_add_51_79_groupi_n_7969);
  and csa_tree_add_51_79_groupi_g37849(csa_tree_add_51_79_groupi_n_8324 ,csa_tree_add_51_79_groupi_n_7541 ,csa_tree_add_51_79_groupi_n_7972);
  or csa_tree_add_51_79_groupi_g37850(csa_tree_add_51_79_groupi_n_8323 ,csa_tree_add_51_79_groupi_n_7545 ,csa_tree_add_51_79_groupi_n_7960);
  and csa_tree_add_51_79_groupi_g37851(csa_tree_add_51_79_groupi_n_8322 ,csa_tree_add_51_79_groupi_n_7546 ,csa_tree_add_51_79_groupi_n_7952);
  and csa_tree_add_51_79_groupi_g37852(csa_tree_add_51_79_groupi_n_8321 ,csa_tree_add_51_79_groupi_n_7549 ,csa_tree_add_51_79_groupi_n_7975);
  and csa_tree_add_51_79_groupi_g37853(csa_tree_add_51_79_groupi_n_8320 ,csa_tree_add_51_79_groupi_n_7554 ,csa_tree_add_51_79_groupi_n_7995);
  and csa_tree_add_51_79_groupi_g37854(csa_tree_add_51_79_groupi_n_8319 ,csa_tree_add_51_79_groupi_n_7438 ,csa_tree_add_51_79_groupi_n_7850);
  and csa_tree_add_51_79_groupi_g37855(csa_tree_add_51_79_groupi_n_8318 ,csa_tree_add_51_79_groupi_n_7562 ,csa_tree_add_51_79_groupi_n_8001);
  and csa_tree_add_51_79_groupi_g37856(csa_tree_add_51_79_groupi_n_8317 ,csa_tree_add_51_79_groupi_n_7434 ,csa_tree_add_51_79_groupi_n_7858);
  and csa_tree_add_51_79_groupi_g37857(csa_tree_add_51_79_groupi_n_8316 ,csa_tree_add_51_79_groupi_n_7430 ,csa_tree_add_51_79_groupi_n_7870);
  or csa_tree_add_51_79_groupi_g37858(csa_tree_add_51_79_groupi_n_8315 ,csa_tree_add_51_79_groupi_n_7569 ,csa_tree_add_51_79_groupi_n_7986);
  and csa_tree_add_51_79_groupi_g37859(csa_tree_add_51_79_groupi_n_8314 ,csa_tree_add_51_79_groupi_n_7421 ,csa_tree_add_51_79_groupi_n_7799);
  and csa_tree_add_51_79_groupi_g37860(csa_tree_add_51_79_groupi_n_8313 ,csa_tree_add_51_79_groupi_n_7570 ,csa_tree_add_51_79_groupi_n_8010);
  and csa_tree_add_51_79_groupi_g37861(csa_tree_add_51_79_groupi_n_8312 ,csa_tree_add_51_79_groupi_n_7572 ,csa_tree_add_51_79_groupi_n_8009);
  and csa_tree_add_51_79_groupi_g37862(csa_tree_add_51_79_groupi_n_8311 ,csa_tree_add_51_79_groupi_n_7463 ,csa_tree_add_51_79_groupi_n_7859);
  and csa_tree_add_51_79_groupi_g37863(csa_tree_add_51_79_groupi_n_8310 ,csa_tree_add_51_79_groupi_n_7534 ,csa_tree_add_51_79_groupi_n_7968);
  and csa_tree_add_51_79_groupi_g37864(csa_tree_add_51_79_groupi_n_8309 ,csa_tree_add_51_79_groupi_n_7462 ,csa_tree_add_51_79_groupi_n_7856);
  and csa_tree_add_51_79_groupi_g37865(csa_tree_add_51_79_groupi_n_8308 ,csa_tree_add_51_79_groupi_n_7537 ,csa_tree_add_51_79_groupi_n_7970);
  and csa_tree_add_51_79_groupi_g37866(csa_tree_add_51_79_groupi_n_8307 ,csa_tree_add_51_79_groupi_n_7485 ,csa_tree_add_51_79_groupi_n_7895);
  and csa_tree_add_51_79_groupi_g37867(csa_tree_add_51_79_groupi_n_8305 ,csa_tree_add_51_79_groupi_n_7483 ,csa_tree_add_51_79_groupi_n_7903);
  or csa_tree_add_51_79_groupi_g37868(csa_tree_add_51_79_groupi_n_8304 ,csa_tree_add_51_79_groupi_n_7506 ,csa_tree_add_51_79_groupi_n_7927);
  and csa_tree_add_51_79_groupi_g37869(csa_tree_add_51_79_groupi_n_8302 ,csa_tree_add_51_79_groupi_n_7450 ,csa_tree_add_51_79_groupi_n_8014);
  and csa_tree_add_51_79_groupi_g37870(csa_tree_add_51_79_groupi_n_8301 ,csa_tree_add_51_79_groupi_n_7492 ,csa_tree_add_51_79_groupi_n_7905);
  and csa_tree_add_51_79_groupi_g37871(csa_tree_add_51_79_groupi_n_8300 ,csa_tree_add_51_79_groupi_n_7543 ,csa_tree_add_51_79_groupi_n_7973);
  and csa_tree_add_51_79_groupi_g37872(csa_tree_add_51_79_groupi_n_8299 ,csa_tree_add_51_79_groupi_n_7493 ,csa_tree_add_51_79_groupi_n_7907);
  and csa_tree_add_51_79_groupi_g37873(csa_tree_add_51_79_groupi_n_8298 ,csa_tree_add_51_79_groupi_n_7458 ,csa_tree_add_51_79_groupi_n_7852);
  and csa_tree_add_51_79_groupi_g37874(csa_tree_add_51_79_groupi_n_8297 ,csa_tree_add_51_79_groupi_n_7547 ,csa_tree_add_51_79_groupi_n_7977);
  and csa_tree_add_51_79_groupi_g37875(csa_tree_add_51_79_groupi_n_8296 ,csa_tree_add_51_79_groupi_n_7445 ,csa_tree_add_51_79_groupi_n_7836);
  and csa_tree_add_51_79_groupi_g37876(csa_tree_add_51_79_groupi_n_8295 ,csa_tree_add_51_79_groupi_n_7517 ,csa_tree_add_51_79_groupi_n_7928);
  and csa_tree_add_51_79_groupi_g37877(csa_tree_add_51_79_groupi_n_8293 ,csa_tree_add_51_79_groupi_n_7552 ,csa_tree_add_51_79_groupi_n_7992);
  and csa_tree_add_51_79_groupi_g37878(csa_tree_add_51_79_groupi_n_8292 ,csa_tree_add_51_79_groupi_n_7518 ,csa_tree_add_51_79_groupi_n_7938);
  and csa_tree_add_51_79_groupi_g37879(csa_tree_add_51_79_groupi_n_8291 ,csa_tree_add_51_79_groupi_n_7556 ,csa_tree_add_51_79_groupi_n_7991);
  and csa_tree_add_51_79_groupi_g37880(csa_tree_add_51_79_groupi_n_8290 ,csa_tree_add_51_79_groupi_n_7557 ,csa_tree_add_51_79_groupi_n_7998);
  and csa_tree_add_51_79_groupi_g37881(csa_tree_add_51_79_groupi_n_8289 ,csa_tree_add_51_79_groupi_n_7560 ,csa_tree_add_51_79_groupi_n_8000);
  and csa_tree_add_51_79_groupi_g37882(csa_tree_add_51_79_groupi_n_8288 ,csa_tree_add_51_79_groupi_n_7455 ,csa_tree_add_51_79_groupi_n_7851);
  and csa_tree_add_51_79_groupi_g37883(csa_tree_add_51_79_groupi_n_8287 ,csa_tree_add_51_79_groupi_n_7519 ,csa_tree_add_51_79_groupi_n_7937);
  and csa_tree_add_51_79_groupi_g37884(csa_tree_add_51_79_groupi_n_8286 ,csa_tree_add_51_79_groupi_n_7470 ,csa_tree_add_51_79_groupi_n_7872);
  and csa_tree_add_51_79_groupi_g37885(csa_tree_add_51_79_groupi_n_8285 ,csa_tree_add_51_79_groupi_n_7521 ,csa_tree_add_51_79_groupi_n_7935);
  and csa_tree_add_51_79_groupi_g37886(csa_tree_add_51_79_groupi_n_8284 ,csa_tree_add_51_79_groupi_n_7496 ,csa_tree_add_51_79_groupi_n_7909);
  and csa_tree_add_51_79_groupi_g37887(csa_tree_add_51_79_groupi_n_8283 ,csa_tree_add_51_79_groupi_n_7433 ,csa_tree_add_51_79_groupi_n_7853);
  or csa_tree_add_51_79_groupi_g37888(csa_tree_add_51_79_groupi_n_8282 ,csa_tree_add_51_79_groupi_n_7432 ,csa_tree_add_51_79_groupi_n_7798);
  and csa_tree_add_51_79_groupi_g37889(csa_tree_add_51_79_groupi_n_8280 ,csa_tree_add_51_79_groupi_n_7522 ,csa_tree_add_51_79_groupi_n_7940);
  and csa_tree_add_51_79_groupi_g37890(csa_tree_add_51_79_groupi_n_8279 ,csa_tree_add_51_79_groupi_n_7566 ,csa_tree_add_51_79_groupi_n_8006);
  and csa_tree_add_51_79_groupi_g37891(csa_tree_add_51_79_groupi_n_8278 ,csa_tree_add_51_79_groupi_n_7567 ,csa_tree_add_51_79_groupi_n_8004);
  and csa_tree_add_51_79_groupi_g37892(csa_tree_add_51_79_groupi_n_8277 ,csa_tree_add_51_79_groupi_n_7397 ,csa_tree_add_51_79_groupi_n_8007);
  and csa_tree_add_51_79_groupi_g37893(csa_tree_add_51_79_groupi_n_8276 ,csa_tree_add_51_79_groupi_n_7472 ,csa_tree_add_51_79_groupi_n_7884);
  and csa_tree_add_51_79_groupi_g37894(csa_tree_add_51_79_groupi_n_8274 ,csa_tree_add_51_79_groupi_n_7419 ,csa_tree_add_51_79_groupi_n_7787);
  and csa_tree_add_51_79_groupi_g37895(csa_tree_add_51_79_groupi_n_8273 ,csa_tree_add_51_79_groupi_n_7424 ,csa_tree_add_51_79_groupi_n_7801);
  and csa_tree_add_51_79_groupi_g37896(csa_tree_add_51_79_groupi_n_8271 ,csa_tree_add_51_79_groupi_n_7423 ,csa_tree_add_51_79_groupi_n_7800);
  and csa_tree_add_51_79_groupi_g37897(csa_tree_add_51_79_groupi_n_8270 ,csa_tree_add_51_79_groupi_n_7527 ,csa_tree_add_51_79_groupi_n_7953);
  and csa_tree_add_51_79_groupi_g37898(csa_tree_add_51_79_groupi_n_8269 ,csa_tree_add_51_79_groupi_n_7416 ,csa_tree_add_51_79_groupi_n_7796);
  and csa_tree_add_51_79_groupi_g37899(csa_tree_add_51_79_groupi_n_8268 ,csa_tree_add_51_79_groupi_n_7497 ,csa_tree_add_51_79_groupi_n_7910);
  or csa_tree_add_51_79_groupi_g37900(csa_tree_add_51_79_groupi_n_8267 ,csa_tree_add_51_79_groupi_n_7428 ,csa_tree_add_51_79_groupi_n_7980);
  and csa_tree_add_51_79_groupi_g37901(csa_tree_add_51_79_groupi_n_8265 ,csa_tree_add_51_79_groupi_n_7447 ,csa_tree_add_51_79_groupi_n_7855);
  not csa_tree_add_51_79_groupi_g37902(csa_tree_add_51_79_groupi_n_8171 ,csa_tree_add_51_79_groupi_n_8172);
  not csa_tree_add_51_79_groupi_g37903(csa_tree_add_51_79_groupi_n_8164 ,csa_tree_add_51_79_groupi_n_8165);
  not csa_tree_add_51_79_groupi_g37904(csa_tree_add_51_79_groupi_n_8163 ,csa_tree_add_51_79_groupi_n_8162);
  not csa_tree_add_51_79_groupi_g37905(csa_tree_add_51_79_groupi_n_8159 ,csa_tree_add_51_79_groupi_n_8158);
  or csa_tree_add_51_79_groupi_g37906(csa_tree_add_51_79_groupi_n_8150 ,csa_tree_add_51_79_groupi_n_6924 ,csa_tree_add_51_79_groupi_n_7790);
  nor csa_tree_add_51_79_groupi_g37907(csa_tree_add_51_79_groupi_n_8149 ,csa_tree_add_51_79_groupi_n_8022 ,csa_tree_add_51_79_groupi_n_7822);
  or csa_tree_add_51_79_groupi_g37908(csa_tree_add_51_79_groupi_n_8148 ,csa_tree_add_51_79_groupi_n_6922 ,csa_tree_add_51_79_groupi_n_7792);
  or csa_tree_add_51_79_groupi_g37909(csa_tree_add_51_79_groupi_n_8147 ,csa_tree_add_51_79_groupi_n_7352 ,csa_tree_add_51_79_groupi_n_7789);
  and csa_tree_add_51_79_groupi_g37910(csa_tree_add_51_79_groupi_n_8146 ,csa_tree_add_51_79_groupi_n_7387 ,csa_tree_add_51_79_groupi_n_7786);
  or csa_tree_add_51_79_groupi_g37911(csa_tree_add_51_79_groupi_n_8145 ,csa_tree_add_51_79_groupi_n_7282 ,csa_tree_add_51_79_groupi_n_7805);
  and csa_tree_add_51_79_groupi_g37912(csa_tree_add_51_79_groupi_n_8144 ,csa_tree_add_51_79_groupi_n_7282 ,csa_tree_add_51_79_groupi_n_7805);
  or csa_tree_add_51_79_groupi_g37913(csa_tree_add_51_79_groupi_n_8143 ,csa_tree_add_51_79_groupi_n_7103 ,csa_tree_add_51_79_groupi_n_7948);
  or csa_tree_add_51_79_groupi_g37914(csa_tree_add_51_79_groupi_n_8142 ,csa_tree_add_51_79_groupi_n_7363 ,csa_tree_add_51_79_groupi_n_7779);
  or csa_tree_add_51_79_groupi_g37915(csa_tree_add_51_79_groupi_n_8141 ,csa_tree_add_51_79_groupi_n_7270 ,csa_tree_add_51_79_groupi_n_7826);
  and csa_tree_add_51_79_groupi_g37916(csa_tree_add_51_79_groupi_n_8140 ,csa_tree_add_51_79_groupi_n_7270 ,csa_tree_add_51_79_groupi_n_7826);
  xor csa_tree_add_51_79_groupi_g37917(out1[0] ,csa_tree_add_51_79_groupi_n_2 ,csa_tree_add_51_79_groupi_n_7118);
  or csa_tree_add_51_79_groupi_g37918(csa_tree_add_51_79_groupi_n_8138 ,csa_tree_add_51_79_groupi_n_7817 ,csa_tree_add_51_79_groupi_n_7317);
  nor csa_tree_add_51_79_groupi_g37919(csa_tree_add_51_79_groupi_n_8137 ,csa_tree_add_51_79_groupi_n_7351 ,csa_tree_add_51_79_groupi_n_7861);
  or csa_tree_add_51_79_groupi_g37920(csa_tree_add_51_79_groupi_n_8136 ,csa_tree_add_51_79_groupi_n_7353 ,csa_tree_add_51_79_groupi_n_7726);
  or csa_tree_add_51_79_groupi_g37921(csa_tree_add_51_79_groupi_n_8135 ,csa_tree_add_51_79_groupi_n_7371 ,csa_tree_add_51_79_groupi_n_7771);
  or csa_tree_add_51_79_groupi_g37922(csa_tree_add_51_79_groupi_n_8134 ,csa_tree_add_51_79_groupi_n_7384 ,csa_tree_add_51_79_groupi_n_7766);
  or csa_tree_add_51_79_groupi_g37923(csa_tree_add_51_79_groupi_n_8133 ,csa_tree_add_51_79_groupi_n_7379 ,csa_tree_add_51_79_groupi_n_7763);
  or csa_tree_add_51_79_groupi_g37924(csa_tree_add_51_79_groupi_n_8132 ,csa_tree_add_51_79_groupi_n_7355 ,csa_tree_add_51_79_groupi_n_7757);
  or csa_tree_add_51_79_groupi_g37925(csa_tree_add_51_79_groupi_n_8131 ,csa_tree_add_51_79_groupi_n_7375 ,csa_tree_add_51_79_groupi_n_7753);
  or csa_tree_add_51_79_groupi_g37926(csa_tree_add_51_79_groupi_n_8130 ,csa_tree_add_51_79_groupi_n_7374 ,csa_tree_add_51_79_groupi_n_7760);
  or csa_tree_add_51_79_groupi_g37927(csa_tree_add_51_79_groupi_n_8129 ,csa_tree_add_51_79_groupi_n_7829 ,csa_tree_add_51_79_groupi_n_7748);
  or csa_tree_add_51_79_groupi_g37928(csa_tree_add_51_79_groupi_n_8128 ,csa_tree_add_51_79_groupi_n_7373 ,csa_tree_add_51_79_groupi_n_7746);
  or csa_tree_add_51_79_groupi_g37929(csa_tree_add_51_79_groupi_n_8127 ,csa_tree_add_51_79_groupi_n_7369 ,csa_tree_add_51_79_groupi_n_7745);
  or csa_tree_add_51_79_groupi_g37930(csa_tree_add_51_79_groupi_n_8126 ,csa_tree_add_51_79_groupi_n_7367 ,csa_tree_add_51_79_groupi_n_7743);
  or csa_tree_add_51_79_groupi_g37931(csa_tree_add_51_79_groupi_n_8125 ,csa_tree_add_51_79_groupi_n_7366 ,csa_tree_add_51_79_groupi_n_7741);
  or csa_tree_add_51_79_groupi_g37932(csa_tree_add_51_79_groupi_n_8124 ,csa_tree_add_51_79_groupi_n_7365 ,csa_tree_add_51_79_groupi_n_7768);
  or csa_tree_add_51_79_groupi_g37933(csa_tree_add_51_79_groupi_n_8123 ,csa_tree_add_51_79_groupi_n_7358 ,csa_tree_add_51_79_groupi_n_7737);
  or csa_tree_add_51_79_groupi_g37934(csa_tree_add_51_79_groupi_n_8122 ,csa_tree_add_51_79_groupi_n_6429 ,csa_tree_add_51_79_groupi_n_7812);
  nor csa_tree_add_51_79_groupi_g37935(csa_tree_add_51_79_groupi_n_8121 ,csa_tree_add_51_79_groupi_n_6430 ,csa_tree_add_51_79_groupi_n_7811);
  or csa_tree_add_51_79_groupi_g37936(csa_tree_add_51_79_groupi_n_8120 ,csa_tree_add_51_79_groupi_n_6919 ,csa_tree_add_51_79_groupi_n_7847);
  and csa_tree_add_51_79_groupi_g37937(csa_tree_add_51_79_groupi_n_8119 ,csa_tree_add_51_79_groupi_n_7817 ,csa_tree_add_51_79_groupi_n_7317);
  xnor csa_tree_add_51_79_groupi_g37938(csa_tree_add_51_79_groupi_n_8118 ,csa_tree_add_51_79_groupi_n_7199 ,csa_tree_add_51_79_groupi_n_7191);
  xnor csa_tree_add_51_79_groupi_g37939(csa_tree_add_51_79_groupi_n_8117 ,csa_tree_add_51_79_groupi_n_7221 ,csa_tree_add_51_79_groupi_n_7222);
  xor csa_tree_add_51_79_groupi_g37940(csa_tree_add_51_79_groupi_n_8116 ,csa_tree_add_51_79_groupi_n_6405 ,csa_tree_add_51_79_groupi_n_7623);
  xnor csa_tree_add_51_79_groupi_g37941(csa_tree_add_51_79_groupi_n_8115 ,csa_tree_add_51_79_groupi_n_7268 ,csa_tree_add_51_79_groupi_n_7147);
  xor csa_tree_add_51_79_groupi_g37942(csa_tree_add_51_79_groupi_n_8114 ,csa_tree_add_51_79_groupi_n_7151 ,csa_tree_add_51_79_groupi_n_7388);
  xnor csa_tree_add_51_79_groupi_g37943(csa_tree_add_51_79_groupi_n_8113 ,csa_tree_add_51_79_groupi_n_6418 ,csa_tree_add_51_79_groupi_n_7240);
  xnor csa_tree_add_51_79_groupi_g37944(csa_tree_add_51_79_groupi_n_8112 ,csa_tree_add_51_79_groupi_n_6426 ,csa_tree_add_51_79_groupi_n_7137);
  xnor csa_tree_add_51_79_groupi_g37945(csa_tree_add_51_79_groupi_n_8111 ,csa_tree_add_51_79_groupi_n_7595 ,csa_tree_add_51_79_groupi_n_7209);
  xnor csa_tree_add_51_79_groupi_g37946(csa_tree_add_51_79_groupi_n_8110 ,csa_tree_add_51_79_groupi_n_7338 ,csa_tree_add_51_79_groupi_n_7616);
  xnor csa_tree_add_51_79_groupi_g37947(csa_tree_add_51_79_groupi_n_8109 ,csa_tree_add_51_79_groupi_n_7232 ,csa_tree_add_51_79_groupi_n_7629);
  xnor csa_tree_add_51_79_groupi_g37948(csa_tree_add_51_79_groupi_n_8108 ,csa_tree_add_51_79_groupi_n_7635 ,csa_tree_add_51_79_groupi_n_7194);
  xnor csa_tree_add_51_79_groupi_g37949(csa_tree_add_51_79_groupi_n_8107 ,csa_tree_add_51_79_groupi_n_7359 ,csa_tree_add_51_79_groupi_n_7181);
  xnor csa_tree_add_51_79_groupi_g37950(csa_tree_add_51_79_groupi_n_8106 ,csa_tree_add_51_79_groupi_n_6437 ,csa_tree_add_51_79_groupi_n_10);
  xnor csa_tree_add_51_79_groupi_g37951(csa_tree_add_51_79_groupi_n_8105 ,csa_tree_add_51_79_groupi_n_7332 ,csa_tree_add_51_79_groupi_n_7599);
  xnor csa_tree_add_51_79_groupi_g37952(csa_tree_add_51_79_groupi_n_8104 ,csa_tree_add_51_79_groupi_n_6409 ,csa_tree_add_51_79_groupi_n_7626);
  xnor csa_tree_add_51_79_groupi_g37953(csa_tree_add_51_79_groupi_n_8103 ,csa_tree_add_51_79_groupi_n_7287 ,csa_tree_add_51_79_groupi_n_7179);
  xnor csa_tree_add_51_79_groupi_g37954(csa_tree_add_51_79_groupi_n_8102 ,csa_tree_add_51_79_groupi_n_7587 ,csa_tree_add_51_79_groupi_n_7320);
  xnor csa_tree_add_51_79_groupi_g37955(csa_tree_add_51_79_groupi_n_8101 ,csa_tree_add_51_79_groupi_n_0 ,csa_tree_add_51_79_groupi_n_7187);
  xnor csa_tree_add_51_79_groupi_g37956(csa_tree_add_51_79_groupi_n_8100 ,csa_tree_add_51_79_groupi_n_7350 ,csa_tree_add_51_79_groupi_n_7167);
  xnor csa_tree_add_51_79_groupi_g37957(csa_tree_add_51_79_groupi_n_8099 ,csa_tree_add_51_79_groupi_n_7354 ,csa_tree_add_51_79_groupi_n_7310);
  xnor csa_tree_add_51_79_groupi_g37958(csa_tree_add_51_79_groupi_n_8098 ,csa_tree_add_51_79_groupi_n_7627 ,csa_tree_add_51_79_groupi_n_7282);
  xnor csa_tree_add_51_79_groupi_g37959(csa_tree_add_51_79_groupi_n_8097 ,csa_tree_add_51_79_groupi_n_5844 ,csa_tree_add_51_79_groupi_n_7364);
  xnor csa_tree_add_51_79_groupi_g37960(csa_tree_add_51_79_groupi_n_8096 ,csa_tree_add_51_79_groupi_n_7198 ,csa_tree_add_51_79_groupi_n_7159);
  xnor csa_tree_add_51_79_groupi_g37961(csa_tree_add_51_79_groupi_n_8095 ,csa_tree_add_51_79_groupi_n_6923 ,csa_tree_add_51_79_groupi_n_7256);
  xnor csa_tree_add_51_79_groupi_g37962(csa_tree_add_51_79_groupi_n_8094 ,csa_tree_add_51_79_groupi_n_7183 ,csa_tree_add_51_79_groupi_n_6971);
  xnor csa_tree_add_51_79_groupi_g37963(csa_tree_add_51_79_groupi_n_8093 ,csa_tree_add_51_79_groupi_n_6407 ,csa_tree_add_51_79_groupi_n_7589);
  xnor csa_tree_add_51_79_groupi_g37964(csa_tree_add_51_79_groupi_n_8092 ,csa_tree_add_51_79_groupi_n_7612 ,csa_tree_add_51_79_groupi_n_7322);
  xnor csa_tree_add_51_79_groupi_g37965(csa_tree_add_51_79_groupi_n_8091 ,csa_tree_add_51_79_groupi_n_7313 ,csa_tree_add_51_79_groupi_n_6906);
  xnor csa_tree_add_51_79_groupi_g37966(csa_tree_add_51_79_groupi_n_8090 ,csa_tree_add_51_79_groupi_n_7353 ,csa_tree_add_51_79_groupi_n_7262);
  xnor csa_tree_add_51_79_groupi_g37967(csa_tree_add_51_79_groupi_n_8089 ,csa_tree_add_51_79_groupi_n_7140 ,csa_tree_add_51_79_groupi_n_7352);
  xnor csa_tree_add_51_79_groupi_g37968(csa_tree_add_51_79_groupi_n_8088 ,csa_tree_add_51_79_groupi_n_7284 ,csa_tree_add_51_79_groupi_n_7360);
  xnor csa_tree_add_51_79_groupi_g37969(csa_tree_add_51_79_groupi_n_8087 ,csa_tree_add_51_79_groupi_n_7153 ,csa_tree_add_51_79_groupi_n_7362);
  xnor csa_tree_add_51_79_groupi_g37970(csa_tree_add_51_79_groupi_n_8086 ,csa_tree_add_51_79_groupi_n_7150 ,csa_tree_add_51_79_groupi_n_7361);
  xnor csa_tree_add_51_79_groupi_g37971(csa_tree_add_51_79_groupi_n_8085 ,csa_tree_add_51_79_groupi_n_7278 ,csa_tree_add_51_79_groupi_n_7283);
  xnor csa_tree_add_51_79_groupi_g37972(csa_tree_add_51_79_groupi_n_8084 ,csa_tree_add_51_79_groupi_n_7210 ,csa_tree_add_51_79_groupi_n_7213);
  xnor csa_tree_add_51_79_groupi_g37973(csa_tree_add_51_79_groupi_n_8083 ,csa_tree_add_51_79_groupi_n_7358 ,csa_tree_add_51_79_groupi_n_7285);
  xnor csa_tree_add_51_79_groupi_g37974(csa_tree_add_51_79_groupi_n_8082 ,csa_tree_add_51_79_groupi_n_7384 ,csa_tree_add_51_79_groupi_n_7258);
  xnor csa_tree_add_51_79_groupi_g37975(csa_tree_add_51_79_groupi_n_8081 ,csa_tree_add_51_79_groupi_n_7223 ,csa_tree_add_51_79_groupi_n_7357);
  xnor csa_tree_add_51_79_groupi_g37976(csa_tree_add_51_79_groupi_n_8080 ,csa_tree_add_51_79_groupi_n_7224 ,csa_tree_add_51_79_groupi_n_7272);
  xnor csa_tree_add_51_79_groupi_g37977(csa_tree_add_51_79_groupi_n_8079 ,csa_tree_add_51_79_groupi_n_7238 ,csa_tree_add_51_79_groupi_n_7280);
  xnor csa_tree_add_51_79_groupi_g37978(csa_tree_add_51_79_groupi_n_8078 ,csa_tree_add_51_79_groupi_n_7225 ,csa_tree_add_51_79_groupi_n_7386);
  xnor csa_tree_add_51_79_groupi_g37979(csa_tree_add_51_79_groupi_n_8077 ,csa_tree_add_51_79_groupi_n_7335 ,csa_tree_add_51_79_groupi_n_7254);
  xnor csa_tree_add_51_79_groupi_g37980(csa_tree_add_51_79_groupi_n_8076 ,csa_tree_add_51_79_groupi_n_7383 ,csa_tree_add_51_79_groupi_n_7252);
  xnor csa_tree_add_51_79_groupi_g37981(csa_tree_add_51_79_groupi_n_8075 ,csa_tree_add_51_79_groupi_n_7356 ,csa_tree_add_51_79_groupi_n_7237);
  xnor csa_tree_add_51_79_groupi_g37982(csa_tree_add_51_79_groupi_n_8074 ,csa_tree_add_51_79_groupi_n_7331 ,csa_tree_add_51_79_groupi_n_7242);
  xnor csa_tree_add_51_79_groupi_g37983(csa_tree_add_51_79_groupi_n_8073 ,csa_tree_add_51_79_groupi_n_7273 ,csa_tree_add_51_79_groupi_n_7253);
  xnor csa_tree_add_51_79_groupi_g37984(csa_tree_add_51_79_groupi_n_8072 ,csa_tree_add_51_79_groupi_n_7248 ,csa_tree_add_51_79_groupi_n_7382);
  xnor csa_tree_add_51_79_groupi_g37985(csa_tree_add_51_79_groupi_n_8071 ,csa_tree_add_51_79_groupi_n_7203 ,csa_tree_add_51_79_groupi_n_7378);
  xnor csa_tree_add_51_79_groupi_g37986(csa_tree_add_51_79_groupi_n_8070 ,csa_tree_add_51_79_groupi_n_7192 ,csa_tree_add_51_79_groupi_n_6442);
  xnor csa_tree_add_51_79_groupi_g37987(csa_tree_add_51_79_groupi_n_8069 ,csa_tree_add_51_79_groupi_n_7205 ,csa_tree_add_51_79_groupi_n_7271);
  xnor csa_tree_add_51_79_groupi_g37988(csa_tree_add_51_79_groupi_n_8068 ,csa_tree_add_51_79_groupi_n_7233 ,csa_tree_add_51_79_groupi_n_7376);
  xnor csa_tree_add_51_79_groupi_g37989(csa_tree_add_51_79_groupi_n_8067 ,csa_tree_add_51_79_groupi_n_7269 ,csa_tree_add_51_79_groupi_n_7355);
  xnor csa_tree_add_51_79_groupi_g37990(csa_tree_add_51_79_groupi_n_8066 ,csa_tree_add_51_79_groupi_n_7375 ,csa_tree_add_51_79_groupi_n_7172);
  xnor csa_tree_add_51_79_groupi_g37991(csa_tree_add_51_79_groupi_n_8065 ,csa_tree_add_51_79_groupi_n_7266 ,csa_tree_add_51_79_groupi_n_7173);
  xnor csa_tree_add_51_79_groupi_g37992(csa_tree_add_51_79_groupi_n_8064 ,csa_tree_add_51_79_groupi_n_7162 ,csa_tree_add_51_79_groupi_n_7279);
  xnor csa_tree_add_51_79_groupi_g37993(csa_tree_add_51_79_groupi_n_8063 ,csa_tree_add_51_79_groupi_n_7323 ,csa_tree_add_51_79_groupi_n_7265);
  xnor csa_tree_add_51_79_groupi_g37994(csa_tree_add_51_79_groupi_n_8062 ,csa_tree_add_51_79_groupi_n_7371 ,csa_tree_add_51_79_groupi_n_7017);
  xnor csa_tree_add_51_79_groupi_g37995(csa_tree_add_51_79_groupi_n_8061 ,csa_tree_add_51_79_groupi_n_7260 ,csa_tree_add_51_79_groupi_n_7373);
  xnor csa_tree_add_51_79_groupi_g37996(csa_tree_add_51_79_groupi_n_8060 ,csa_tree_add_51_79_groupi_n_7308 ,csa_tree_add_51_79_groupi_n_7610);
  xnor csa_tree_add_51_79_groupi_g37997(csa_tree_add_51_79_groupi_n_8059 ,csa_tree_add_51_79_groupi_n_7369 ,csa_tree_add_51_79_groupi_n_7305);
  xnor csa_tree_add_51_79_groupi_g37998(csa_tree_add_51_79_groupi_n_8058 ,csa_tree_add_51_79_groupi_n_7302 ,csa_tree_add_51_79_groupi_n_6857);
  xnor csa_tree_add_51_79_groupi_g37999(csa_tree_add_51_79_groupi_n_8057 ,csa_tree_add_51_79_groupi_n_7583 ,csa_tree_add_51_79_groupi_n_7220);
  xnor csa_tree_add_51_79_groupi_g38000(csa_tree_add_51_79_groupi_n_8056 ,csa_tree_add_51_79_groupi_n_7365 ,csa_tree_add_51_79_groupi_n_7294);
  xnor csa_tree_add_51_79_groupi_g38001(csa_tree_add_51_79_groupi_n_8055 ,csa_tree_add_51_79_groupi_n_7298 ,csa_tree_add_51_79_groupi_n_7299);
  xnor csa_tree_add_51_79_groupi_g38002(csa_tree_add_51_79_groupi_n_8054 ,csa_tree_add_51_79_groupi_n_7297 ,csa_tree_add_51_79_groupi_n_7366);
  xnor csa_tree_add_51_79_groupi_g38003(csa_tree_add_51_79_groupi_n_8053 ,csa_tree_add_51_79_groupi_n_7264 ,csa_tree_add_51_79_groupi_n_7227);
  xnor csa_tree_add_51_79_groupi_g38004(csa_tree_add_51_79_groupi_n_8052 ,csa_tree_add_51_79_groupi_n_7330 ,csa_tree_add_51_79_groupi_n_7157);
  xnor csa_tree_add_51_79_groupi_g38005(csa_tree_add_51_79_groupi_n_8051 ,csa_tree_add_51_79_groupi_n_6412 ,csa_tree_add_51_79_groupi_n_7618);
  xnor csa_tree_add_51_79_groupi_g38006(csa_tree_add_51_79_groupi_n_8050 ,csa_tree_add_51_79_groupi_n_7171 ,csa_tree_add_51_79_groupi_n_6900);
  xnor csa_tree_add_51_79_groupi_g38007(csa_tree_add_51_79_groupi_n_8049 ,csa_tree_add_51_79_groupi_n_6850 ,csa_tree_add_51_79_groupi_n_7609);
  xnor csa_tree_add_51_79_groupi_g38008(csa_tree_add_51_79_groupi_n_8048 ,csa_tree_add_51_79_groupi_n_7333 ,csa_tree_add_51_79_groupi_n_7217);
  xnor csa_tree_add_51_79_groupi_g38009(csa_tree_add_51_79_groupi_n_8047 ,csa_tree_add_51_79_groupi_n_7176 ,csa_tree_add_51_79_groupi_n_7177);
  xnor csa_tree_add_51_79_groupi_g38010(csa_tree_add_51_79_groupi_n_8046 ,csa_tree_add_51_79_groupi_n_7155 ,csa_tree_add_51_79_groupi_n_7325);
  xnor csa_tree_add_51_79_groupi_g38011(csa_tree_add_51_79_groupi_n_8045 ,csa_tree_add_51_79_groupi_n_7200 ,csa_tree_add_51_79_groupi_n_7634);
  xnor csa_tree_add_51_79_groupi_g38012(csa_tree_add_51_79_groupi_n_8044 ,csa_tree_add_51_79_groupi_n_7143 ,csa_tree_add_51_79_groupi_n_6922);
  xnor csa_tree_add_51_79_groupi_g38013(csa_tree_add_51_79_groupi_n_8043 ,csa_tree_add_51_79_groupi_n_7342 ,csa_tree_add_51_79_groupi_n_6399);
  xnor csa_tree_add_51_79_groupi_g38014(csa_tree_add_51_79_groupi_n_8042 ,csa_tree_add_51_79_groupi_n_7251 ,csa_tree_add_51_79_groupi_n_7387);
  xnor csa_tree_add_51_79_groupi_g38015(csa_tree_add_51_79_groupi_n_8041 ,csa_tree_add_51_79_groupi_n_9 ,csa_tree_add_51_79_groupi_n_7296);
  xnor csa_tree_add_51_79_groupi_g38016(csa_tree_add_51_79_groupi_n_8040 ,csa_tree_add_51_79_groupi_n_6420 ,csa_tree_add_51_79_groupi_n_7304);
  xnor csa_tree_add_51_79_groupi_g38017(csa_tree_add_51_79_groupi_n_8039 ,csa_tree_add_51_79_groupi_n_7321 ,csa_tree_add_51_79_groupi_n_7244);
  xnor csa_tree_add_51_79_groupi_g38018(csa_tree_add_51_79_groupi_n_8038 ,csa_tree_add_51_79_groupi_n_7229 ,csa_tree_add_51_79_groupi_n_7337);
  xnor csa_tree_add_51_79_groupi_g38019(csa_tree_add_51_79_groupi_n_8037 ,csa_tree_add_51_79_groupi_n_6415 ,csa_tree_add_51_79_groupi_n_7189);
  xnor csa_tree_add_51_79_groupi_g38020(csa_tree_add_51_79_groupi_n_8036 ,csa_tree_add_51_79_groupi_n_7275 ,csa_tree_add_51_79_groupi_n_7578);
  xnor csa_tree_add_51_79_groupi_g38021(csa_tree_add_51_79_groupi_n_8035 ,csa_tree_add_51_79_groupi_n_6961 ,csa_tree_add_51_79_groupi_n_7585);
  xnor csa_tree_add_51_79_groupi_g38022(csa_tree_add_51_79_groupi_n_8034 ,csa_tree_add_51_79_groupi_n_6402 ,csa_tree_add_51_79_groupi_n_7630);
  xor csa_tree_add_51_79_groupi_g38023(csa_tree_add_51_79_groupi_n_8033 ,csa_tree_add_51_79_groupi_n_7601 ,csa_tree_add_51_79_groupi_n_7625);
  xnor csa_tree_add_51_79_groupi_g38024(csa_tree_add_51_79_groupi_n_8032 ,csa_tree_add_51_79_groupi_n_6424 ,csa_tree_add_51_79_groupi_n_7348);
  and csa_tree_add_51_79_groupi_g38025(csa_tree_add_51_79_groupi_n_8185 ,csa_tree_add_51_79_groupi_n_7410 ,csa_tree_add_51_79_groupi_n_7775);
  xnor csa_tree_add_51_79_groupi_g38026(csa_tree_add_51_79_groupi_n_8184 ,csa_tree_add_51_79_groupi_n_6753 ,csa_tree_add_51_79_groupi_n_7123);
  xnor csa_tree_add_51_79_groupi_g38027(csa_tree_add_51_79_groupi_n_8183 ,csa_tree_add_51_79_groupi_n_7115 ,csa_tree_add_51_79_groupi_n_7135);
  xnor csa_tree_add_51_79_groupi_g38028(csa_tree_add_51_79_groupi_n_8182 ,csa_tree_add_51_79_groupi_n_7070 ,csa_tree_add_51_79_groupi_n_7125);
  and csa_tree_add_51_79_groupi_g38029(csa_tree_add_51_79_groupi_n_8181 ,csa_tree_add_51_79_groupi_n_7487 ,csa_tree_add_51_79_groupi_n_7736);
  xnor csa_tree_add_51_79_groupi_g38030(csa_tree_add_51_79_groupi_n_8180 ,csa_tree_add_51_79_groupi_n_6454 ,csa_tree_add_51_79_groupi_n_7129);
  and csa_tree_add_51_79_groupi_g38031(csa_tree_add_51_79_groupi_n_8179 ,csa_tree_add_51_79_groupi_n_7406 ,csa_tree_add_51_79_groupi_n_7773);
  and csa_tree_add_51_79_groupi_g38032(csa_tree_add_51_79_groupi_n_8178 ,csa_tree_add_51_79_groupi_n_7412 ,csa_tree_add_51_79_groupi_n_7776);
  xnor csa_tree_add_51_79_groupi_g38033(csa_tree_add_51_79_groupi_n_8177 ,csa_tree_add_51_79_groupi_n_6938 ,csa_tree_add_51_79_groupi_n_7121);
  xnor csa_tree_add_51_79_groupi_g38034(csa_tree_add_51_79_groupi_n_8176 ,csa_tree_add_51_79_groupi_n_6441 ,csa_tree_add_51_79_groupi_n_7132);
  and csa_tree_add_51_79_groupi_g38035(csa_tree_add_51_79_groupi_n_8175 ,csa_tree_add_51_79_groupi_n_7503 ,csa_tree_add_51_79_groupi_n_7729);
  xnor csa_tree_add_51_79_groupi_g38036(csa_tree_add_51_79_groupi_n_8174 ,csa_tree_add_51_79_groupi_n_6397 ,csa_tree_add_51_79_groupi_n_7130);
  and csa_tree_add_51_79_groupi_g38037(csa_tree_add_51_79_groupi_n_8173 ,csa_tree_add_51_79_groupi_n_7399 ,csa_tree_add_51_79_groupi_n_7735);
  xnor csa_tree_add_51_79_groupi_g38038(csa_tree_add_51_79_groupi_n_8172 ,csa_tree_add_51_79_groupi_n_7349 ,csa_tree_add_51_79_groupi_n_7119);
  xnor csa_tree_add_51_79_groupi_g38039(csa_tree_add_51_79_groupi_n_8170 ,csa_tree_add_51_79_groupi_n_6761 ,csa_tree_add_51_79_groupi_n_7128);
  xnor csa_tree_add_51_79_groupi_g38040(csa_tree_add_51_79_groupi_n_8169 ,csa_tree_add_51_79_groupi_n_6459 ,csa_tree_add_51_79_groupi_n_7127);
  and csa_tree_add_51_79_groupi_g38041(csa_tree_add_51_79_groupi_n_8168 ,csa_tree_add_51_79_groupi_n_7392 ,csa_tree_add_51_79_groupi_n_7733);
  and csa_tree_add_51_79_groupi_g38042(csa_tree_add_51_79_groupi_n_8167 ,csa_tree_add_51_79_groupi_n_7425 ,csa_tree_add_51_79_groupi_n_7734);
  and csa_tree_add_51_79_groupi_g38043(csa_tree_add_51_79_groupi_n_8166 ,csa_tree_add_51_79_groupi_n_7426 ,csa_tree_add_51_79_groupi_n_7732);
  and csa_tree_add_51_79_groupi_g38044(csa_tree_add_51_79_groupi_n_8165 ,csa_tree_add_51_79_groupi_n_6782 ,csa_tree_add_51_79_groupi_n_7724);
  and csa_tree_add_51_79_groupi_g38045(csa_tree_add_51_79_groupi_n_8162 ,csa_tree_add_51_79_groupi_n_7529 ,csa_tree_add_51_79_groupi_n_7723);
  and csa_tree_add_51_79_groupi_g38046(csa_tree_add_51_79_groupi_n_8161 ,csa_tree_add_51_79_groupi_n_7390 ,csa_tree_add_51_79_groupi_n_7731);
  and csa_tree_add_51_79_groupi_g38047(csa_tree_add_51_79_groupi_n_8160 ,csa_tree_add_51_79_groupi_n_7446 ,csa_tree_add_51_79_groupi_n_7730);
  xnor csa_tree_add_51_79_groupi_g38048(csa_tree_add_51_79_groupi_n_8158 ,csa_tree_add_51_79_groupi_n_6912 ,csa_tree_add_51_79_groupi_n_7126);
  xnor csa_tree_add_51_79_groupi_g38049(csa_tree_add_51_79_groupi_n_8157 ,csa_tree_add_51_79_groupi_n_6904 ,csa_tree_add_51_79_groupi_n_7124);
  xnor csa_tree_add_51_79_groupi_g38050(csa_tree_add_51_79_groupi_n_8156 ,csa_tree_add_51_79_groupi_n_6732 ,csa_tree_add_51_79_groupi_n_7134);
  xnor csa_tree_add_51_79_groupi_g38051(csa_tree_add_51_79_groupi_n_8155 ,csa_tree_add_51_79_groupi_n_6458 ,csa_tree_add_51_79_groupi_n_7122);
  xnor csa_tree_add_51_79_groupi_g38052(csa_tree_add_51_79_groupi_n_8154 ,csa_tree_add_51_79_groupi_n_6456 ,csa_tree_add_51_79_groupi_n_7133);
  xnor csa_tree_add_51_79_groupi_g38053(csa_tree_add_51_79_groupi_n_8153 ,csa_tree_add_51_79_groupi_n_6724 ,csa_tree_add_51_79_groupi_n_7131);
  xnor csa_tree_add_51_79_groupi_g38054(csa_tree_add_51_79_groupi_n_8152 ,csa_tree_add_51_79_groupi_n_6453 ,csa_tree_add_51_79_groupi_n_7120);
  and csa_tree_add_51_79_groupi_g38055(csa_tree_add_51_79_groupi_n_8151 ,csa_tree_add_51_79_groupi_n_7409 ,csa_tree_add_51_79_groupi_n_7774);
  not csa_tree_add_51_79_groupi_g38056(csa_tree_add_51_79_groupi_n_8029 ,csa_tree_add_51_79_groupi_n_8028);
  not csa_tree_add_51_79_groupi_g38057(csa_tree_add_51_79_groupi_n_8024 ,csa_tree_add_51_79_groupi_n_8025);
  not csa_tree_add_51_79_groupi_g38058(csa_tree_add_51_79_groupi_n_8021 ,csa_tree_add_51_79_groupi_n_8022);
  not csa_tree_add_51_79_groupi_g38059(csa_tree_add_51_79_groupi_n_8018 ,csa_tree_add_51_79_groupi_n_8019);
  or csa_tree_add_51_79_groupi_g38060(csa_tree_add_51_79_groupi_n_8014 ,csa_tree_add_51_79_groupi_n_6901 ,csa_tree_add_51_79_groupi_n_7466);
  nor csa_tree_add_51_79_groupi_g38061(csa_tree_add_51_79_groupi_n_8013 ,csa_tree_add_51_79_groupi_n_7156 ,csa_tree_add_51_79_groupi_n_7161);
  or csa_tree_add_51_79_groupi_g38062(csa_tree_add_51_79_groupi_n_8012 ,csa_tree_add_51_79_groupi_n_6960 ,csa_tree_add_51_79_groupi_n_7584);
  nor csa_tree_add_51_79_groupi_g38063(csa_tree_add_51_79_groupi_n_8011 ,csa_tree_add_51_79_groupi_n_6961 ,csa_tree_add_51_79_groupi_n_7585);
  or csa_tree_add_51_79_groupi_g38064(csa_tree_add_51_79_groupi_n_8010 ,csa_tree_add_51_79_groupi_n_7064 ,csa_tree_add_51_79_groupi_n_7568);
  or csa_tree_add_51_79_groupi_g38065(csa_tree_add_51_79_groupi_n_8009 ,csa_tree_add_51_79_groupi_n_7066 ,csa_tree_add_51_79_groupi_n_7565);
  or csa_tree_add_51_79_groupi_g38066(csa_tree_add_51_79_groupi_n_8008 ,csa_tree_add_51_79_groupi_n_6971 ,csa_tree_add_51_79_groupi_n_7183);
  or csa_tree_add_51_79_groupi_g38067(csa_tree_add_51_79_groupi_n_8007 ,csa_tree_add_51_79_groupi_n_7069 ,csa_tree_add_51_79_groupi_n_7396);
  or csa_tree_add_51_79_groupi_g38068(csa_tree_add_51_79_groupi_n_8006 ,csa_tree_add_51_79_groupi_n_7071 ,csa_tree_add_51_79_groupi_n_7564);
  or csa_tree_add_51_79_groupi_g38069(csa_tree_add_51_79_groupi_n_8005 ,csa_tree_add_51_79_groupi_n_7280 ,csa_tree_add_51_79_groupi_n_7238);
  or csa_tree_add_51_79_groupi_g38070(csa_tree_add_51_79_groupi_n_8004 ,csa_tree_add_51_79_groupi_n_7077 ,csa_tree_add_51_79_groupi_n_7563);
  and csa_tree_add_51_79_groupi_g38071(csa_tree_add_51_79_groupi_n_8003 ,csa_tree_add_51_79_groupi_n_7280 ,csa_tree_add_51_79_groupi_n_7238);
  or csa_tree_add_51_79_groupi_g38072(csa_tree_add_51_79_groupi_n_8002 ,csa_tree_add_51_79_groupi_n_7284 ,csa_tree_add_51_79_groupi_n_7148);
  or csa_tree_add_51_79_groupi_g38073(csa_tree_add_51_79_groupi_n_8001 ,csa_tree_add_51_79_groupi_n_7078 ,csa_tree_add_51_79_groupi_n_7559);
  or csa_tree_add_51_79_groupi_g38074(csa_tree_add_51_79_groupi_n_8000 ,csa_tree_add_51_79_groupi_n_7080 ,csa_tree_add_51_79_groupi_n_7558);
  nor csa_tree_add_51_79_groupi_g38075(csa_tree_add_51_79_groupi_n_7999 ,csa_tree_add_51_79_groupi_n_6401 ,csa_tree_add_51_79_groupi_n_7235);
  or csa_tree_add_51_79_groupi_g38076(csa_tree_add_51_79_groupi_n_7998 ,csa_tree_add_51_79_groupi_n_7088 ,csa_tree_add_51_79_groupi_n_7555);
  or csa_tree_add_51_79_groupi_g38077(csa_tree_add_51_79_groupi_n_7997 ,csa_tree_add_51_79_groupi_n_6402 ,csa_tree_add_51_79_groupi_n_7234);
  or csa_tree_add_51_79_groupi_g38078(csa_tree_add_51_79_groupi_n_7996 ,csa_tree_add_51_79_groupi_n_7579 ,csa_tree_add_51_79_groupi_n_7615);
  or csa_tree_add_51_79_groupi_g38079(csa_tree_add_51_79_groupi_n_7995 ,csa_tree_add_51_79_groupi_n_7098 ,csa_tree_add_51_79_groupi_n_7553);
  nor csa_tree_add_51_79_groupi_g38080(csa_tree_add_51_79_groupi_n_7994 ,csa_tree_add_51_79_groupi_n_7580 ,csa_tree_add_51_79_groupi_n_7616);
  nor csa_tree_add_51_79_groupi_g38081(csa_tree_add_51_79_groupi_n_7993 ,csa_tree_add_51_79_groupi_n_7613 ,csa_tree_add_51_79_groupi_n_7232);
  or csa_tree_add_51_79_groupi_g38082(csa_tree_add_51_79_groupi_n_7992 ,csa_tree_add_51_79_groupi_n_7100 ,csa_tree_add_51_79_groupi_n_7551);
  or csa_tree_add_51_79_groupi_g38083(csa_tree_add_51_79_groupi_n_7991 ,csa_tree_add_51_79_groupi_n_7106 ,csa_tree_add_51_79_groupi_n_7550);
  or csa_tree_add_51_79_groupi_g38084(csa_tree_add_51_79_groupi_n_7990 ,csa_tree_add_51_79_groupi_n_7614 ,csa_tree_add_51_79_groupi_n_7231);
  or csa_tree_add_51_79_groupi_g38085(csa_tree_add_51_79_groupi_n_7989 ,csa_tree_add_51_79_groupi_n_7277 ,csa_tree_add_51_79_groupi_n_7230);
  and csa_tree_add_51_79_groupi_g38086(csa_tree_add_51_79_groupi_n_7988 ,csa_tree_add_51_79_groupi_n_7277 ,csa_tree_add_51_79_groupi_n_7230);
  or csa_tree_add_51_79_groupi_g38087(csa_tree_add_51_79_groupi_n_7987 ,csa_tree_add_51_79_groupi_n_7229 ,csa_tree_add_51_79_groupi_n_7228);
  and csa_tree_add_51_79_groupi_g38088(csa_tree_add_51_79_groupi_n_7986 ,csa_tree_add_51_79_groupi_n_7085 ,csa_tree_add_51_79_groupi_n_7548);
  and csa_tree_add_51_79_groupi_g38089(csa_tree_add_51_79_groupi_n_7985 ,csa_tree_add_51_79_groupi_n_7229 ,csa_tree_add_51_79_groupi_n_7228);
  or csa_tree_add_51_79_groupi_g38090(csa_tree_add_51_79_groupi_n_7984 ,csa_tree_add_51_79_groupi_n_7226 ,csa_tree_add_51_79_groupi_n_7225);
  and csa_tree_add_51_79_groupi_g38091(csa_tree_add_51_79_groupi_n_7983 ,csa_tree_add_51_79_groupi_n_7226 ,csa_tree_add_51_79_groupi_n_7225);
  or csa_tree_add_51_79_groupi_g38092(csa_tree_add_51_79_groupi_n_7982 ,csa_tree_add_51_79_groupi_n_7272 ,csa_tree_add_51_79_groupi_n_7224);
  and csa_tree_add_51_79_groupi_g38093(csa_tree_add_51_79_groupi_n_7981 ,csa_tree_add_51_79_groupi_n_7272 ,csa_tree_add_51_79_groupi_n_7224);
  nor csa_tree_add_51_79_groupi_g38094(csa_tree_add_51_79_groupi_n_7980 ,csa_tree_add_51_79_groupi_n_7114 ,csa_tree_add_51_79_groupi_n_7507);
  or csa_tree_add_51_79_groupi_g38095(csa_tree_add_51_79_groupi_n_7979 ,csa_tree_add_51_79_groupi_n_7263 ,csa_tree_add_51_79_groupi_n_7223);
  and csa_tree_add_51_79_groupi_g38096(csa_tree_add_51_79_groupi_n_7978 ,csa_tree_add_51_79_groupi_n_7263 ,csa_tree_add_51_79_groupi_n_7223);
  or csa_tree_add_51_79_groupi_g38097(csa_tree_add_51_79_groupi_n_7977 ,csa_tree_add_51_79_groupi_n_7116 ,csa_tree_add_51_79_groupi_n_7544);
  or csa_tree_add_51_79_groupi_g38098(csa_tree_add_51_79_groupi_n_7976 ,csa_tree_add_51_79_groupi_n_7244 ,csa_tree_add_51_79_groupi_n_7288);
  or csa_tree_add_51_79_groupi_g38099(csa_tree_add_51_79_groupi_n_7975 ,csa_tree_add_51_79_groupi_n_7089 ,csa_tree_add_51_79_groupi_n_7536);
  and csa_tree_add_51_79_groupi_g38100(csa_tree_add_51_79_groupi_n_7974 ,csa_tree_add_51_79_groupi_n_7150 ,csa_tree_add_51_79_groupi_n_7149);
  or csa_tree_add_51_79_groupi_g38101(csa_tree_add_51_79_groupi_n_7973 ,csa_tree_add_51_79_groupi_n_7113 ,csa_tree_add_51_79_groupi_n_7540);
  or csa_tree_add_51_79_groupi_g38102(csa_tree_add_51_79_groupi_n_7972 ,csa_tree_add_51_79_groupi_n_7112 ,csa_tree_add_51_79_groupi_n_7539);
  nor csa_tree_add_51_79_groupi_g38103(csa_tree_add_51_79_groupi_n_7971 ,csa_tree_add_51_79_groupi_n_6409 ,csa_tree_add_51_79_groupi_n_7604);
  or csa_tree_add_51_79_groupi_g38104(csa_tree_add_51_79_groupi_n_7970 ,csa_tree_add_51_79_groupi_n_7111 ,csa_tree_add_51_79_groupi_n_7535);
  or csa_tree_add_51_79_groupi_g38105(csa_tree_add_51_79_groupi_n_7969 ,csa_tree_add_51_79_groupi_n_7110 ,csa_tree_add_51_79_groupi_n_7533);
  or csa_tree_add_51_79_groupi_g38106(csa_tree_add_51_79_groupi_n_7968 ,csa_tree_add_51_79_groupi_n_7109 ,csa_tree_add_51_79_groupi_n_7532);
  or csa_tree_add_51_79_groupi_g38107(csa_tree_add_51_79_groupi_n_7967 ,csa_tree_add_51_79_groupi_n_6408 ,csa_tree_add_51_79_groupi_n_7605);
  or csa_tree_add_51_79_groupi_g38108(csa_tree_add_51_79_groupi_n_7966 ,csa_tree_add_51_79_groupi_n_6742 ,csa_tree_add_51_79_groupi_n_7602);
  or csa_tree_add_51_79_groupi_g38109(csa_tree_add_51_79_groupi_n_7965 ,csa_tree_add_51_79_groupi_n_7222 ,csa_tree_add_51_79_groupi_n_7221);
  or csa_tree_add_51_79_groupi_g38110(csa_tree_add_51_79_groupi_n_7964 ,csa_tree_add_51_79_groupi_n_7108 ,csa_tree_add_51_79_groupi_n_7530);
  and csa_tree_add_51_79_groupi_g38111(csa_tree_add_51_79_groupi_n_7963 ,csa_tree_add_51_79_groupi_n_7222 ,csa_tree_add_51_79_groupi_n_7221);
  nor csa_tree_add_51_79_groupi_g38112(csa_tree_add_51_79_groupi_n_7962 ,csa_tree_add_51_79_groupi_n_6741 ,csa_tree_add_51_79_groupi_n_7603);
  or csa_tree_add_51_79_groupi_g38113(csa_tree_add_51_79_groupi_n_7961 ,csa_tree_add_51_79_groupi_n_6403 ,csa_tree_add_51_79_groupi_n_7217);
  and csa_tree_add_51_79_groupi_g38114(csa_tree_add_51_79_groupi_n_7960 ,csa_tree_add_51_79_groupi_n_7624 ,csa_tree_add_51_79_groupi_n_7528);
  or csa_tree_add_51_79_groupi_g38115(csa_tree_add_51_79_groupi_n_7959 ,csa_tree_add_51_79_groupi_n_7252 ,csa_tree_add_51_79_groupi_n_7212);
  nor csa_tree_add_51_79_groupi_g38116(csa_tree_add_51_79_groupi_n_7958 ,csa_tree_add_51_79_groupi_n_6404 ,csa_tree_add_51_79_groupi_n_7216);
  and csa_tree_add_51_79_groupi_g38117(csa_tree_add_51_79_groupi_n_7957 ,csa_tree_add_51_79_groupi_n_7601 ,csa_tree_add_51_79_groupi_n_7600);
  and csa_tree_add_51_79_groupi_g38118(csa_tree_add_51_79_groupi_n_7956 ,csa_tree_add_51_79_groupi_n_7252 ,csa_tree_add_51_79_groupi_n_7212);
  or csa_tree_add_51_79_groupi_g38119(csa_tree_add_51_79_groupi_n_7955 ,csa_tree_add_51_79_groupi_n_1530 ,csa_tree_add_51_79_groupi_n_7211);
  nor csa_tree_add_51_79_groupi_g38120(csa_tree_add_51_79_groupi_n_7954 ,csa_tree_add_51_79_groupi_n_7601 ,csa_tree_add_51_79_groupi_n_7600);
  or csa_tree_add_51_79_groupi_g38121(csa_tree_add_51_79_groupi_n_7953 ,csa_tree_add_51_79_groupi_n_7105 ,csa_tree_add_51_79_groupi_n_7526);
  or csa_tree_add_51_79_groupi_g38122(csa_tree_add_51_79_groupi_n_7952 ,csa_tree_add_51_79_groupi_n_7104 ,csa_tree_add_51_79_groupi_n_7523);
  and csa_tree_add_51_79_groupi_g38124(csa_tree_add_51_79_groupi_n_7951 ,csa_tree_add_51_79_groupi_n_6405 ,csa_tree_add_51_79_groupi_n_7593);
  or csa_tree_add_51_79_groupi_g38125(csa_tree_add_51_79_groupi_n_7950 ,csa_tree_add_51_79_groupi_n_7594 ,csa_tree_add_51_79_groupi_n_7209);
  nor csa_tree_add_51_79_groupi_g38126(csa_tree_add_51_79_groupi_n_7949 ,csa_tree_add_51_79_groupi_n_6418 ,csa_tree_add_51_79_groupi_n_7239);
  nor csa_tree_add_51_79_groupi_g38127(csa_tree_add_51_79_groupi_n_7948 ,csa_tree_add_51_79_groupi_n_7595 ,csa_tree_add_51_79_groupi_n_7208);
  nor csa_tree_add_51_79_groupi_g38128(csa_tree_add_51_79_groupi_n_7947 ,csa_tree_add_51_79_groupi_n_6423 ,csa_tree_add_51_79_groupi_n_7185);
  or csa_tree_add_51_79_groupi_g38129(csa_tree_add_51_79_groupi_n_7946 ,csa_tree_add_51_79_groupi_n_7248 ,csa_tree_add_51_79_groupi_n_7207);
  nor csa_tree_add_51_79_groupi_g38130(csa_tree_add_51_79_groupi_n_7945 ,csa_tree_add_51_79_groupi_n_6405 ,csa_tree_add_51_79_groupi_n_7593);
  and csa_tree_add_51_79_groupi_g38131(csa_tree_add_51_79_groupi_n_7944 ,csa_tree_add_51_79_groupi_n_7248 ,csa_tree_add_51_79_groupi_n_7207);
  or csa_tree_add_51_79_groupi_g38132(csa_tree_add_51_79_groupi_n_7943 ,csa_tree_add_51_79_groupi_n_6406 ,csa_tree_add_51_79_groupi_n_7588);
  nor csa_tree_add_51_79_groupi_g38133(csa_tree_add_51_79_groupi_n_7942 ,csa_tree_add_51_79_groupi_n_6437 ,csa_tree_add_51_79_groupi_n_7590);
  or csa_tree_add_51_79_groupi_g38134(csa_tree_add_51_79_groupi_n_7941 ,csa_tree_add_51_79_groupi_n_6436 ,csa_tree_add_51_79_groupi_n_10);
  or csa_tree_add_51_79_groupi_g38135(csa_tree_add_51_79_groupi_n_7940 ,csa_tree_add_51_79_groupi_n_7099 ,csa_tree_add_51_79_groupi_n_7520);
  nor csa_tree_add_51_79_groupi_g38136(csa_tree_add_51_79_groupi_n_7939 ,csa_tree_add_51_79_groupi_n_6407 ,csa_tree_add_51_79_groupi_n_7589);
  or csa_tree_add_51_79_groupi_g38137(csa_tree_add_51_79_groupi_n_7938 ,csa_tree_add_51_79_groupi_n_7096 ,csa_tree_add_51_79_groupi_n_7516);
  or csa_tree_add_51_79_groupi_g38138(csa_tree_add_51_79_groupi_n_7937 ,csa_tree_add_51_79_groupi_n_7095 ,csa_tree_add_51_79_groupi_n_7514);
  or csa_tree_add_51_79_groupi_g38139(csa_tree_add_51_79_groupi_n_7936 ,csa_tree_add_51_79_groupi_n_7094 ,csa_tree_add_51_79_groupi_n_7512);
  or csa_tree_add_51_79_groupi_g38140(csa_tree_add_51_79_groupi_n_7935 ,csa_tree_add_51_79_groupi_n_7093 ,csa_tree_add_51_79_groupi_n_7510);
  or csa_tree_add_51_79_groupi_g38141(csa_tree_add_51_79_groupi_n_7934 ,csa_tree_add_51_79_groupi_n_7150 ,csa_tree_add_51_79_groupi_n_7149);
  and csa_tree_add_51_79_groupi_g38142(csa_tree_add_51_79_groupi_n_7933 ,csa_tree_add_51_79_groupi_n_7596 ,csa_tree_add_51_79_groupi_n_7153);
  or csa_tree_add_51_79_groupi_g38143(csa_tree_add_51_79_groupi_n_7932 ,csa_tree_add_51_79_groupi_n_7092 ,csa_tree_add_51_79_groupi_n_7508);
  or csa_tree_add_51_79_groupi_g38144(csa_tree_add_51_79_groupi_n_7931 ,csa_tree_add_51_79_groupi_n_7271 ,csa_tree_add_51_79_groupi_n_7205);
  and csa_tree_add_51_79_groupi_g38145(csa_tree_add_51_79_groupi_n_7930 ,csa_tree_add_51_79_groupi_n_7271 ,csa_tree_add_51_79_groupi_n_7205);
  or csa_tree_add_51_79_groupi_g38146(csa_tree_add_51_79_groupi_n_7929 ,csa_tree_add_51_79_groupi_n_7022 ,csa_tree_add_51_79_groupi_n_7202);
  or csa_tree_add_51_79_groupi_g38147(csa_tree_add_51_79_groupi_n_7928 ,csa_tree_add_51_79_groupi_n_7087 ,csa_tree_add_51_79_groupi_n_7484);
  and csa_tree_add_51_79_groupi_g38148(csa_tree_add_51_79_groupi_n_7927 ,csa_tree_add_51_79_groupi_n_7091 ,csa_tree_add_51_79_groupi_n_7504);
  and csa_tree_add_51_79_groupi_g38149(csa_tree_add_51_79_groupi_n_7926 ,csa_tree_add_51_79_groupi_n_7022 ,csa_tree_add_51_79_groupi_n_7202);
  or csa_tree_add_51_79_groupi_g38150(csa_tree_add_51_79_groupi_n_7925 ,csa_tree_add_51_79_groupi_n_7117 ,csa_tree_add_51_79_groupi_n_7502);
  or csa_tree_add_51_79_groupi_g38151(csa_tree_add_51_79_groupi_n_7924 ,csa_tree_add_51_79_groupi_n_7165 ,csa_tree_add_51_79_groupi_n_7200);
  or csa_tree_add_51_79_groupi_g38152(csa_tree_add_51_79_groupi_n_7923 ,csa_tree_add_51_79_groupi_n_7203 ,csa_tree_add_51_79_groupi_n_7201);
  and csa_tree_add_51_79_groupi_g38153(csa_tree_add_51_79_groupi_n_7922 ,csa_tree_add_51_79_groupi_n_7203 ,csa_tree_add_51_79_groupi_n_7201);
  or csa_tree_add_51_79_groupi_g38154(csa_tree_add_51_79_groupi_n_7921 ,csa_tree_add_51_79_groupi_n_7191 ,csa_tree_add_51_79_groupi_n_7199);
  and csa_tree_add_51_79_groupi_g38155(csa_tree_add_51_79_groupi_n_7920 ,csa_tree_add_51_79_groupi_n_7191 ,csa_tree_add_51_79_groupi_n_7199);
  and csa_tree_add_51_79_groupi_g38156(csa_tree_add_51_79_groupi_n_7919 ,csa_tree_add_51_79_groupi_n_7165 ,csa_tree_add_51_79_groupi_n_7200);
  nor csa_tree_add_51_79_groupi_g38157(csa_tree_add_51_79_groupi_n_7918 ,csa_tree_add_51_79_groupi_n_6398 ,csa_tree_add_51_79_groupi_n_7219);
  nor csa_tree_add_51_79_groupi_g38158(csa_tree_add_51_79_groupi_n_7917 ,csa_tree_add_51_79_groupi_n_6411 ,csa_tree_add_51_79_groupi_n_7196);
  or csa_tree_add_51_79_groupi_g38159(csa_tree_add_51_79_groupi_n_7916 ,csa_tree_add_51_79_groupi_n_6412 ,csa_tree_add_51_79_groupi_n_7195);
  nor csa_tree_add_51_79_groupi_g38160(csa_tree_add_51_79_groupi_n_7915 ,csa_tree_add_51_79_groupi_n_7581 ,csa_tree_add_51_79_groupi_n_7194);
  or csa_tree_add_51_79_groupi_g38161(csa_tree_add_51_79_groupi_n_7914 ,csa_tree_add_51_79_groupi_n_7086 ,csa_tree_add_51_79_groupi_n_7499);
  or csa_tree_add_51_79_groupi_g38162(csa_tree_add_51_79_groupi_n_7913 ,csa_tree_add_51_79_groupi_n_7582 ,csa_tree_add_51_79_groupi_n_7193);
  or csa_tree_add_51_79_groupi_g38163(csa_tree_add_51_79_groupi_n_7912 ,csa_tree_add_51_79_groupi_n_6442 ,csa_tree_add_51_79_groupi_n_7192);
  and csa_tree_add_51_79_groupi_g38164(csa_tree_add_51_79_groupi_n_7911 ,csa_tree_add_51_79_groupi_n_6442 ,csa_tree_add_51_79_groupi_n_7192);
  or csa_tree_add_51_79_groupi_g38165(csa_tree_add_51_79_groupi_n_7910 ,csa_tree_add_51_79_groupi_n_7081 ,csa_tree_add_51_79_groupi_n_7489);
  or csa_tree_add_51_79_groupi_g38166(csa_tree_add_51_79_groupi_n_7909 ,csa_tree_add_51_79_groupi_n_7083 ,csa_tree_add_51_79_groupi_n_7494);
  or csa_tree_add_51_79_groupi_g38167(csa_tree_add_51_79_groupi_n_7908 ,csa_tree_add_51_79_groupi_n_7617 ,csa_tree_add_51_79_groupi_n_7490);
  or csa_tree_add_51_79_groupi_g38168(csa_tree_add_51_79_groupi_n_7907 ,csa_tree_add_51_79_groupi_n_7079 ,csa_tree_add_51_79_groupi_n_7488);
  or csa_tree_add_51_79_groupi_g38169(csa_tree_add_51_79_groupi_n_7906 ,csa_tree_add_51_79_groupi_n_7233 ,csa_tree_add_51_79_groupi_n_7190);
  or csa_tree_add_51_79_groupi_g38170(csa_tree_add_51_79_groupi_n_7905 ,csa_tree_add_51_79_groupi_n_7076 ,csa_tree_add_51_79_groupi_n_7481);
  and csa_tree_add_51_79_groupi_g38171(csa_tree_add_51_79_groupi_n_7904 ,csa_tree_add_51_79_groupi_n_7233 ,csa_tree_add_51_79_groupi_n_7190);
  or csa_tree_add_51_79_groupi_g38172(csa_tree_add_51_79_groupi_n_7903 ,csa_tree_add_51_79_groupi_n_7073 ,csa_tree_add_51_79_groupi_n_7482);
  or csa_tree_add_51_79_groupi_g38173(csa_tree_add_51_79_groupi_n_7902 ,csa_tree_add_51_79_groupi_n_7206 ,csa_tree_add_51_79_groupi_n_7187);
  nor csa_tree_add_51_79_groupi_g38174(csa_tree_add_51_79_groupi_n_7901 ,csa_tree_add_51_79_groupi_n_0 ,csa_tree_add_51_79_groupi_n_7186);
  or csa_tree_add_51_79_groupi_g38175(csa_tree_add_51_79_groupi_n_7900 ,csa_tree_add_51_79_groupi_n_7072 ,csa_tree_add_51_79_groupi_n_7477);
  or csa_tree_add_51_79_groupi_g38176(csa_tree_add_51_79_groupi_n_7899 ,csa_tree_add_51_79_groupi_n_7152 ,csa_tree_add_51_79_groupi_n_7151);
  or csa_tree_add_51_79_groupi_g38177(csa_tree_add_51_79_groupi_n_7898 ,csa_tree_add_51_79_groupi_n_7067 ,csa_tree_add_51_79_groupi_n_7474);
  or csa_tree_add_51_79_groupi_g38178(csa_tree_add_51_79_groupi_n_7897 ,csa_tree_add_51_79_groupi_n_6909 ,csa_tree_add_51_79_groupi_n_7475);
  or csa_tree_add_51_79_groupi_g38179(csa_tree_add_51_79_groupi_n_7896 ,csa_tree_add_51_79_groupi_n_7596 ,csa_tree_add_51_79_groupi_n_7153);
  or csa_tree_add_51_79_groupi_g38180(csa_tree_add_51_79_groupi_n_7895 ,csa_tree_add_51_79_groupi_n_7065 ,csa_tree_add_51_79_groupi_n_7511);
  or csa_tree_add_51_79_groupi_g38181(csa_tree_add_51_79_groupi_n_7894 ,csa_tree_add_51_79_groupi_n_7062 ,csa_tree_add_51_79_groupi_n_7467);
  and csa_tree_add_51_79_groupi_g38182(csa_tree_add_51_79_groupi_n_7893 ,csa_tree_add_51_79_groupi_n_6957 ,csa_tree_add_51_79_groupi_n_7349);
  or csa_tree_add_51_79_groupi_g38183(csa_tree_add_51_79_groupi_n_7892 ,csa_tree_add_51_79_groupi_n_6755 ,csa_tree_add_51_79_groupi_n_7163);
  or csa_tree_add_51_79_groupi_g38184(csa_tree_add_51_79_groupi_n_7891 ,csa_tree_add_51_79_groupi_n_6424 ,csa_tree_add_51_79_groupi_n_7184);
  and csa_tree_add_51_79_groupi_g38185(csa_tree_add_51_79_groupi_n_7890 ,csa_tree_add_51_79_groupi_n_6971 ,csa_tree_add_51_79_groupi_n_7183);
  nor csa_tree_add_51_79_groupi_g38186(csa_tree_add_51_79_groupi_n_7889 ,csa_tree_add_51_79_groupi_n_7292 ,csa_tree_add_51_79_groupi_n_7181);
  or csa_tree_add_51_79_groupi_g38187(csa_tree_add_51_79_groupi_n_7888 ,csa_tree_add_51_79_groupi_n_7293 ,csa_tree_add_51_79_groupi_n_7180);
  nor csa_tree_add_51_79_groupi_g38188(csa_tree_add_51_79_groupi_n_7887 ,csa_tree_add_51_79_groupi_n_7286 ,csa_tree_add_51_79_groupi_n_7179);
  or csa_tree_add_51_79_groupi_g38189(csa_tree_add_51_79_groupi_n_7886 ,csa_tree_add_51_79_groupi_n_7177 ,csa_tree_add_51_79_groupi_n_7176);
  or csa_tree_add_51_79_groupi_g38190(csa_tree_add_51_79_groupi_n_7885 ,csa_tree_add_51_79_groupi_n_7287 ,csa_tree_add_51_79_groupi_n_7178);
  or csa_tree_add_51_79_groupi_g38191(csa_tree_add_51_79_groupi_n_7884 ,csa_tree_add_51_79_groupi_n_6907 ,csa_tree_add_51_79_groupi_n_7460);
  and csa_tree_add_51_79_groupi_g38192(csa_tree_add_51_79_groupi_n_7883 ,csa_tree_add_51_79_groupi_n_7177 ,csa_tree_add_51_79_groupi_n_7176);
  or csa_tree_add_51_79_groupi_g38193(csa_tree_add_51_79_groupi_n_7882 ,csa_tree_add_51_79_groupi_n_7246 ,csa_tree_add_51_79_groupi_n_7155);
  nor csa_tree_add_51_79_groupi_g38194(csa_tree_add_51_79_groupi_n_7881 ,csa_tree_add_51_79_groupi_n_7247 ,csa_tree_add_51_79_groupi_n_7154);
  or csa_tree_add_51_79_groupi_g38195(csa_tree_add_51_79_groupi_n_7880 ,csa_tree_add_51_79_groupi_n_6414 ,csa_tree_add_51_79_groupi_n_7188);
  or csa_tree_add_51_79_groupi_g38196(csa_tree_add_51_79_groupi_n_7879 ,csa_tree_add_51_79_groupi_n_6899 ,csa_tree_add_51_79_groupi_n_7471);
  or csa_tree_add_51_79_groupi_g38197(csa_tree_add_51_79_groupi_n_7878 ,csa_tree_add_51_79_groupi_n_7314 ,csa_tree_add_51_79_groupi_n_7171);
  or csa_tree_add_51_79_groupi_g38198(csa_tree_add_51_79_groupi_n_7877 ,csa_tree_add_51_79_groupi_n_6417 ,csa_tree_add_51_79_groupi_n_7240);
  and csa_tree_add_51_79_groupi_g38199(csa_tree_add_51_79_groupi_n_7876 ,csa_tree_add_51_79_groupi_n_7314 ,csa_tree_add_51_79_groupi_n_7171);
  or csa_tree_add_51_79_groupi_g38200(csa_tree_add_51_79_groupi_n_7875 ,csa_tree_add_51_79_groupi_n_1529 ,csa_tree_add_51_79_groupi_n_7306);
  nor csa_tree_add_51_79_groupi_g38201(csa_tree_add_51_79_groupi_n_7874 ,csa_tree_add_51_79_groupi_n_1070 ,csa_tree_add_51_79_groupi_n_7307);
  or csa_tree_add_51_79_groupi_g38202(csa_tree_add_51_79_groupi_n_7873 ,csa_tree_add_51_79_groupi_n_6419 ,csa_tree_add_51_79_groupi_n_7303);
  or csa_tree_add_51_79_groupi_g38203(csa_tree_add_51_79_groupi_n_7872 ,csa_tree_add_51_79_groupi_n_6902 ,csa_tree_add_51_79_groupi_n_7469);
  nor csa_tree_add_51_79_groupi_g38204(csa_tree_add_51_79_groupi_n_7871 ,csa_tree_add_51_79_groupi_n_6415 ,csa_tree_add_51_79_groupi_n_7189);
  or csa_tree_add_51_79_groupi_g38205(csa_tree_add_51_79_groupi_n_7870 ,csa_tree_add_51_79_groupi_n_6931 ,csa_tree_add_51_79_groupi_n_7427);
  and csa_tree_add_51_79_groupi_g38206(csa_tree_add_51_79_groupi_n_7869 ,csa_tree_add_51_79_groupi_n_6857 ,csa_tree_add_51_79_groupi_n_7302);
  nor csa_tree_add_51_79_groupi_g38207(csa_tree_add_51_79_groupi_n_7868 ,csa_tree_add_51_79_groupi_n_6426 ,csa_tree_add_51_79_groupi_n_7136);
  nor csa_tree_add_51_79_groupi_g38208(csa_tree_add_51_79_groupi_n_7867 ,csa_tree_add_51_79_groupi_n_6420 ,csa_tree_add_51_79_groupi_n_7304);
  and csa_tree_add_51_79_groupi_g38209(csa_tree_add_51_79_groupi_n_7866 ,csa_tree_add_51_79_groupi_n_9 ,csa_tree_add_51_79_groupi_n_7296);
  or csa_tree_add_51_79_groupi_g38210(csa_tree_add_51_79_groupi_n_7865 ,csa_tree_add_51_79_groupi_n_6728 ,csa_tree_add_51_79_groupi_n_7168);
  or csa_tree_add_51_79_groupi_g38211(csa_tree_add_51_79_groupi_n_7864 ,csa_tree_add_51_79_groupi_n_9 ,csa_tree_add_51_79_groupi_n_7296);
  nor csa_tree_add_51_79_groupi_g38212(csa_tree_add_51_79_groupi_n_7863 ,csa_tree_add_51_79_groupi_n_7291 ,csa_tree_add_51_79_groupi_n_7167);
  or csa_tree_add_51_79_groupi_g38213(csa_tree_add_51_79_groupi_n_7862 ,csa_tree_add_51_79_groupi_n_7274 ,csa_tree_add_51_79_groupi_n_7577);
  and csa_tree_add_51_79_groupi_g38214(csa_tree_add_51_79_groupi_n_7861 ,csa_tree_add_51_79_groupi_n_7291 ,csa_tree_add_51_79_groupi_n_7167);
  and csa_tree_add_51_79_groupi_g38215(csa_tree_add_51_79_groupi_n_7860 ,csa_tree_add_51_79_groupi_n_6728 ,csa_tree_add_51_79_groupi_n_7168);
  or csa_tree_add_51_79_groupi_g38216(csa_tree_add_51_79_groupi_n_7859 ,csa_tree_add_51_79_groupi_n_6910 ,csa_tree_add_51_79_groupi_n_7575);
  or csa_tree_add_51_79_groupi_g38217(csa_tree_add_51_79_groupi_n_7858 ,csa_tree_add_51_79_groupi_n_6932 ,csa_tree_add_51_79_groupi_n_7429);
  or csa_tree_add_51_79_groupi_g38218(csa_tree_add_51_79_groupi_n_7857 ,csa_tree_add_51_79_groupi_n_6857 ,csa_tree_add_51_79_groupi_n_7302);
  or csa_tree_add_51_79_groupi_g38219(csa_tree_add_51_79_groupi_n_7856 ,csa_tree_add_51_79_groupi_n_6908 ,csa_tree_add_51_79_groupi_n_7457);
  or csa_tree_add_51_79_groupi_g38220(csa_tree_add_51_79_groupi_n_7855 ,csa_tree_add_51_79_groupi_n_7084 ,csa_tree_add_51_79_groupi_n_7459);
  or csa_tree_add_51_79_groupi_g38221(csa_tree_add_51_79_groupi_n_7854 ,csa_tree_add_51_79_groupi_n_6911 ,csa_tree_add_51_79_groupi_n_7454);
  or csa_tree_add_51_79_groupi_g38222(csa_tree_add_51_79_groupi_n_7853 ,csa_tree_add_51_79_groupi_n_6933 ,csa_tree_add_51_79_groupi_n_7431);
  or csa_tree_add_51_79_groupi_g38223(csa_tree_add_51_79_groupi_n_7852 ,csa_tree_add_51_79_groupi_n_6914 ,csa_tree_add_51_79_groupi_n_7461);
  or csa_tree_add_51_79_groupi_g38224(csa_tree_add_51_79_groupi_n_7851 ,csa_tree_add_51_79_groupi_n_6936 ,csa_tree_add_51_79_groupi_n_7435);
  or csa_tree_add_51_79_groupi_g38225(csa_tree_add_51_79_groupi_n_7850 ,csa_tree_add_51_79_groupi_n_6937 ,csa_tree_add_51_79_groupi_n_7436);
  nor csa_tree_add_51_79_groupi_g38226(csa_tree_add_51_79_groupi_n_7849 ,csa_tree_add_51_79_groupi_n_7275 ,csa_tree_add_51_79_groupi_n_7578);
  or csa_tree_add_51_79_groupi_g38227(csa_tree_add_51_79_groupi_n_7848 ,csa_tree_add_51_79_groupi_n_6929 ,csa_tree_add_51_79_groupi_n_7448);
  nor csa_tree_add_51_79_groupi_g38228(csa_tree_add_51_79_groupi_n_7847 ,csa_tree_add_51_79_groupi_n_6754 ,csa_tree_add_51_79_groupi_n_7164);
  nor csa_tree_add_51_79_groupi_g38229(csa_tree_add_51_79_groupi_n_7846 ,csa_tree_add_51_79_groupi_n_6903 ,csa_tree_add_51_79_groupi_n_7571);
  or csa_tree_add_51_79_groupi_g38230(csa_tree_add_51_79_groupi_n_7845 ,csa_tree_add_51_79_groupi_n_7220 ,csa_tree_add_51_79_groupi_n_7583);
  and csa_tree_add_51_79_groupi_g38231(csa_tree_add_51_79_groupi_n_7844 ,csa_tree_add_51_79_groupi_n_7220 ,csa_tree_add_51_79_groupi_n_7583);
  or csa_tree_add_51_79_groupi_g38232(csa_tree_add_51_79_groupi_n_7843 ,csa_tree_add_51_79_groupi_n_6934 ,csa_tree_add_51_79_groupi_n_7444);
  nor csa_tree_add_51_79_groupi_g38233(csa_tree_add_51_79_groupi_n_7842 ,csa_tree_add_51_79_groupi_n_7243 ,csa_tree_add_51_79_groupi_n_7289);
  or csa_tree_add_51_79_groupi_g38234(csa_tree_add_51_79_groupi_n_7841 ,csa_tree_add_51_79_groupi_n_7586 ,csa_tree_add_51_79_groupi_n_7174);
  or csa_tree_add_51_79_groupi_g38235(csa_tree_add_51_79_groupi_n_7840 ,csa_tree_add_51_79_groupi_n_6425 ,csa_tree_add_51_79_groupi_n_7137);
  nor csa_tree_add_51_79_groupi_g38236(csa_tree_add_51_79_groupi_n_7839 ,csa_tree_add_51_79_groupi_n_7587 ,csa_tree_add_51_79_groupi_n_7175);
  nor csa_tree_add_51_79_groupi_g38237(csa_tree_add_51_79_groupi_n_7838 ,csa_tree_add_51_79_groupi_n_7197 ,csa_tree_add_51_79_groupi_n_7159);
  or csa_tree_add_51_79_groupi_g38238(csa_tree_add_51_79_groupi_n_7837 ,csa_tree_add_51_79_groupi_n_7198 ,csa_tree_add_51_79_groupi_n_7158);
  or csa_tree_add_51_79_groupi_g38239(csa_tree_add_51_79_groupi_n_7836 ,csa_tree_add_51_79_groupi_n_6915 ,csa_tree_add_51_79_groupi_n_7441);
  or csa_tree_add_51_79_groupi_g38240(csa_tree_add_51_79_groupi_n_7835 ,csa_tree_add_51_79_groupi_n_7157 ,csa_tree_add_51_79_groupi_n_7160);
  and csa_tree_add_51_79_groupi_g38241(csa_tree_add_51_79_groupi_n_8031 ,csa_tree_add_51_79_groupi_n_6815 ,csa_tree_add_51_79_groupi_n_7468);
  and csa_tree_add_51_79_groupi_g38242(csa_tree_add_51_79_groupi_n_8030 ,csa_tree_add_51_79_groupi_n_6958 ,csa_tree_add_51_79_groupi_n_7453);
  and csa_tree_add_51_79_groupi_g38243(csa_tree_add_51_79_groupi_n_8028 ,csa_tree_add_51_79_groupi_n_6512 ,csa_tree_add_51_79_groupi_n_7573);
  and csa_tree_add_51_79_groupi_g38244(csa_tree_add_51_79_groupi_n_8027 ,csa_tree_add_51_79_groupi_n_6949 ,csa_tree_add_51_79_groupi_n_7486);
  and csa_tree_add_51_79_groupi_g38245(csa_tree_add_51_79_groupi_n_8026 ,csa_tree_add_51_79_groupi_n_6795 ,csa_tree_add_51_79_groupi_n_7452);
  and csa_tree_add_51_79_groupi_g38246(csa_tree_add_51_79_groupi_n_8025 ,csa_tree_add_51_79_groupi_n_6809 ,csa_tree_add_51_79_groupi_n_7451);
  and csa_tree_add_51_79_groupi_g38247(csa_tree_add_51_79_groupi_n_8023 ,csa_tree_add_51_79_groupi_n_6781 ,csa_tree_add_51_79_groupi_n_7439);
  or csa_tree_add_51_79_groupi_g38248(csa_tree_add_51_79_groupi_n_8022 ,csa_tree_add_51_79_groupi_n_6780 ,csa_tree_add_51_79_groupi_n_7440);
  and csa_tree_add_51_79_groupi_g38249(csa_tree_add_51_79_groupi_n_8020 ,csa_tree_add_51_79_groupi_n_6955 ,csa_tree_add_51_79_groupi_n_7476);
  and csa_tree_add_51_79_groupi_g38250(csa_tree_add_51_79_groupi_n_8019 ,csa_tree_add_51_79_groupi_n_6945 ,csa_tree_add_51_79_groupi_n_7437);
  and csa_tree_add_51_79_groupi_g38251(csa_tree_add_51_79_groupi_n_8017 ,csa_tree_add_51_79_groupi_n_6521 ,csa_tree_add_51_79_groupi_n_7443);
  and csa_tree_add_51_79_groupi_g38252(csa_tree_add_51_79_groupi_n_8016 ,csa_tree_add_51_79_groupi_n_6940 ,csa_tree_add_51_79_groupi_n_7542);
  and csa_tree_add_51_79_groupi_g38253(csa_tree_add_51_79_groupi_n_8015 ,csa_tree_add_51_79_groupi_n_6951 ,csa_tree_add_51_79_groupi_n_7561);
  not csa_tree_add_51_79_groupi_g38254(csa_tree_add_51_79_groupi_n_7834 ,csa_tree_add_51_79_groupi_n_7833);
  not csa_tree_add_51_79_groupi_g38255(csa_tree_add_51_79_groupi_n_7824 ,csa_tree_add_51_79_groupi_n_7823);
  not csa_tree_add_51_79_groupi_g38256(csa_tree_add_51_79_groupi_n_7821 ,csa_tree_add_51_79_groupi_n_7822);
  not csa_tree_add_51_79_groupi_g38257(csa_tree_add_51_79_groupi_n_7818 ,csa_tree_add_51_79_groupi_n_7819);
  not csa_tree_add_51_79_groupi_g38258(csa_tree_add_51_79_groupi_n_7814 ,csa_tree_add_51_79_groupi_n_7813);
  not csa_tree_add_51_79_groupi_g38259(csa_tree_add_51_79_groupi_n_7812 ,csa_tree_add_51_79_groupi_n_7811);
  not csa_tree_add_51_79_groupi_g38260(csa_tree_add_51_79_groupi_n_7809 ,csa_tree_add_51_79_groupi_n_7808);
  or csa_tree_add_51_79_groupi_g38261(csa_tree_add_51_79_groupi_n_7802 ,csa_tree_add_51_79_groupi_n_7245 ,csa_tree_add_51_79_groupi_n_7242);
  or csa_tree_add_51_79_groupi_g38262(csa_tree_add_51_79_groupi_n_7801 ,csa_tree_add_51_79_groupi_n_6928 ,csa_tree_add_51_79_groupi_n_7422);
  or csa_tree_add_51_79_groupi_g38263(csa_tree_add_51_79_groupi_n_7800 ,csa_tree_add_51_79_groupi_n_6926 ,csa_tree_add_51_79_groupi_n_7417);
  or csa_tree_add_51_79_groupi_g38264(csa_tree_add_51_79_groupi_n_7799 ,csa_tree_add_51_79_groupi_n_6927 ,csa_tree_add_51_79_groupi_n_7418);
  and csa_tree_add_51_79_groupi_g38265(csa_tree_add_51_79_groupi_n_7798 ,csa_tree_add_51_79_groupi_n_6930 ,csa_tree_add_51_79_groupi_n_7420);
  or csa_tree_add_51_79_groupi_g38266(csa_tree_add_51_79_groupi_n_7797 ,csa_tree_add_51_79_groupi_n_7267 ,csa_tree_add_51_79_groupi_n_7147);
  or csa_tree_add_51_79_groupi_g38267(csa_tree_add_51_79_groupi_n_7796 ,csa_tree_add_51_79_groupi_n_6925 ,csa_tree_add_51_79_groupi_n_7415);
  nor csa_tree_add_51_79_groupi_g38268(csa_tree_add_51_79_groupi_n_7795 ,csa_tree_add_51_79_groupi_n_7268 ,csa_tree_add_51_79_groupi_n_7146);
  or csa_tree_add_51_79_groupi_g38269(csa_tree_add_51_79_groupi_n_7794 ,csa_tree_add_51_79_groupi_n_6427 ,csa_tree_add_51_79_groupi_n_7255);
  or csa_tree_add_51_79_groupi_g38270(csa_tree_add_51_79_groupi_n_7793 ,csa_tree_add_51_79_groupi_n_7143 ,csa_tree_add_51_79_groupi_n_7142);
  and csa_tree_add_51_79_groupi_g38271(csa_tree_add_51_79_groupi_n_7792 ,csa_tree_add_51_79_groupi_n_7143 ,csa_tree_add_51_79_groupi_n_7142);
  or csa_tree_add_51_79_groupi_g38272(csa_tree_add_51_79_groupi_n_7791 ,csa_tree_add_51_79_groupi_n_7141 ,csa_tree_add_51_79_groupi_n_7140);
  nor csa_tree_add_51_79_groupi_g38273(csa_tree_add_51_79_groupi_n_7790 ,csa_tree_add_51_79_groupi_n_6428 ,csa_tree_add_51_79_groupi_n_7256);
  and csa_tree_add_51_79_groupi_g38274(csa_tree_add_51_79_groupi_n_7789 ,csa_tree_add_51_79_groupi_n_7141 ,csa_tree_add_51_79_groupi_n_7140);
  nor csa_tree_add_51_79_groupi_g38275(csa_tree_add_51_79_groupi_n_7788 ,csa_tree_add_51_79_groupi_n_7250 ,csa_tree_add_51_79_groupi_n_7139);
  or csa_tree_add_51_79_groupi_g38276(csa_tree_add_51_79_groupi_n_7787 ,csa_tree_add_51_79_groupi_n_6920 ,csa_tree_add_51_79_groupi_n_7574);
  or csa_tree_add_51_79_groupi_g38277(csa_tree_add_51_79_groupi_n_7786 ,csa_tree_add_51_79_groupi_n_7251 ,csa_tree_add_51_79_groupi_n_7138);
  or csa_tree_add_51_79_groupi_g38278(csa_tree_add_51_79_groupi_n_7785 ,csa_tree_add_51_79_groupi_n_6399 ,csa_tree_add_51_79_groupi_n_7218);
  or csa_tree_add_51_79_groupi_g38279(csa_tree_add_51_79_groupi_n_7784 ,csa_tree_add_51_79_groupi_n_7611 ,csa_tree_add_51_79_groupi_n_7214);
  nor csa_tree_add_51_79_groupi_g38280(csa_tree_add_51_79_groupi_n_7783 ,csa_tree_add_51_79_groupi_n_7612 ,csa_tree_add_51_79_groupi_n_7215);
  or csa_tree_add_51_79_groupi_g38281(csa_tree_add_51_79_groupi_n_7782 ,csa_tree_add_51_79_groupi_n_7576 ,csa_tree_add_51_79_groupi_n_7254);
  and csa_tree_add_51_79_groupi_g38282(csa_tree_add_51_79_groupi_n_7781 ,csa_tree_add_51_79_groupi_n_7576 ,csa_tree_add_51_79_groupi_n_7254);
  or csa_tree_add_51_79_groupi_g38283(csa_tree_add_51_79_groupi_n_7780 ,csa_tree_add_51_79_groupi_n_7610 ,csa_tree_add_51_79_groupi_n_7308);
  and csa_tree_add_51_79_groupi_g38284(csa_tree_add_51_79_groupi_n_7779 ,csa_tree_add_51_79_groupi_n_7610 ,csa_tree_add_51_79_groupi_n_7308);
  or csa_tree_add_51_79_groupi_g38285(csa_tree_add_51_79_groupi_n_7778 ,csa_tree_add_51_79_groupi_n_6849 ,csa_tree_add_51_79_groupi_n_7608);
  nor csa_tree_add_51_79_groupi_g38286(csa_tree_add_51_79_groupi_n_7777 ,csa_tree_add_51_79_groupi_n_6850 ,csa_tree_add_51_79_groupi_n_7609);
  or csa_tree_add_51_79_groupi_g38287(csa_tree_add_51_79_groupi_n_7776 ,csa_tree_add_51_79_groupi_n_7068 ,csa_tree_add_51_79_groupi_n_7411);
  or csa_tree_add_51_79_groupi_g38288(csa_tree_add_51_79_groupi_n_7775 ,csa_tree_add_51_79_groupi_n_6905 ,csa_tree_add_51_79_groupi_n_7407);
  or csa_tree_add_51_79_groupi_g38289(csa_tree_add_51_79_groupi_n_7774 ,csa_tree_add_51_79_groupi_n_6917 ,csa_tree_add_51_79_groupi_n_7408);
  or csa_tree_add_51_79_groupi_g38290(csa_tree_add_51_79_groupi_n_7773 ,csa_tree_add_51_79_groupi_n_6916 ,csa_tree_add_51_79_groupi_n_7405);
  or csa_tree_add_51_79_groupi_g38291(csa_tree_add_51_79_groupi_n_7772 ,csa_tree_add_51_79_groupi_n_7017 ,csa_tree_add_51_79_groupi_n_7311);
  and csa_tree_add_51_79_groupi_g38292(csa_tree_add_51_79_groupi_n_7771 ,csa_tree_add_51_79_groupi_n_7017 ,csa_tree_add_51_79_groupi_n_7311);
  or csa_tree_add_51_79_groupi_g38293(csa_tree_add_51_79_groupi_n_7770 ,csa_tree_add_51_79_groupi_n_7283 ,csa_tree_add_51_79_groupi_n_7278);
  and csa_tree_add_51_79_groupi_g38294(csa_tree_add_51_79_groupi_n_7769 ,csa_tree_add_51_79_groupi_n_7283 ,csa_tree_add_51_79_groupi_n_7278);
  and csa_tree_add_51_79_groupi_g38295(csa_tree_add_51_79_groupi_n_7768 ,csa_tree_add_51_79_groupi_n_7295 ,csa_tree_add_51_79_groupi_n_7294);
  or csa_tree_add_51_79_groupi_g38296(csa_tree_add_51_79_groupi_n_7767 ,csa_tree_add_51_79_groupi_n_7258 ,csa_tree_add_51_79_groupi_n_7257);
  and csa_tree_add_51_79_groupi_g38297(csa_tree_add_51_79_groupi_n_7766 ,csa_tree_add_51_79_groupi_n_7258 ,csa_tree_add_51_79_groupi_n_7257);
  or csa_tree_add_51_79_groupi_g38298(csa_tree_add_51_79_groupi_n_7765 ,csa_tree_add_51_79_groupi_n_7253 ,csa_tree_add_51_79_groupi_n_7273);
  and csa_tree_add_51_79_groupi_g38299(csa_tree_add_51_79_groupi_n_7764 ,csa_tree_add_51_79_groupi_n_7253 ,csa_tree_add_51_79_groupi_n_7273);
  and csa_tree_add_51_79_groupi_g38300(csa_tree_add_51_79_groupi_n_7763 ,csa_tree_add_51_79_groupi_n_7213 ,csa_tree_add_51_79_groupi_n_7210);
  and csa_tree_add_51_79_groupi_g38301(csa_tree_add_51_79_groupi_n_7762 ,csa_tree_add_51_79_groupi_n_7284 ,csa_tree_add_51_79_groupi_n_7148);
  and csa_tree_add_51_79_groupi_g38302(csa_tree_add_51_79_groupi_n_7761 ,csa_tree_add_51_79_groupi_n_7245 ,csa_tree_add_51_79_groupi_n_7242);
  and csa_tree_add_51_79_groupi_g38303(csa_tree_add_51_79_groupi_n_7760 ,csa_tree_add_51_79_groupi_n_7279 ,csa_tree_add_51_79_groupi_n_7162);
  or csa_tree_add_51_79_groupi_g38304(csa_tree_add_51_79_groupi_n_7759 ,csa_tree_add_51_79_groupi_n_7213 ,csa_tree_add_51_79_groupi_n_7210);
  or csa_tree_add_51_79_groupi_g38305(csa_tree_add_51_79_groupi_n_7758 ,csa_tree_add_51_79_groupi_n_7182 ,csa_tree_add_51_79_groupi_n_7269);
  and csa_tree_add_51_79_groupi_g38306(csa_tree_add_51_79_groupi_n_7757 ,csa_tree_add_51_79_groupi_n_7182 ,csa_tree_add_51_79_groupi_n_7269);
  or csa_tree_add_51_79_groupi_g38307(csa_tree_add_51_79_groupi_n_7756 ,csa_tree_add_51_79_groupi_n_7173 ,csa_tree_add_51_79_groupi_n_7266);
  and csa_tree_add_51_79_groupi_g38308(csa_tree_add_51_79_groupi_n_7755 ,csa_tree_add_51_79_groupi_n_7173 ,csa_tree_add_51_79_groupi_n_7266);
  or csa_tree_add_51_79_groupi_g38309(csa_tree_add_51_79_groupi_n_7754 ,csa_tree_add_51_79_groupi_n_7172 ,csa_tree_add_51_79_groupi_n_7166);
  and csa_tree_add_51_79_groupi_g38310(csa_tree_add_51_79_groupi_n_7753 ,csa_tree_add_51_79_groupi_n_7172 ,csa_tree_add_51_79_groupi_n_7166);
  or csa_tree_add_51_79_groupi_g38311(csa_tree_add_51_79_groupi_n_7752 ,csa_tree_add_51_79_groupi_n_7279 ,csa_tree_add_51_79_groupi_n_7162);
  or csa_tree_add_51_79_groupi_g38312(csa_tree_add_51_79_groupi_n_7751 ,csa_tree_add_51_79_groupi_n_7276 ,csa_tree_add_51_79_groupi_n_7265);
  and csa_tree_add_51_79_groupi_g38313(csa_tree_add_51_79_groupi_n_7750 ,csa_tree_add_51_79_groupi_n_7276 ,csa_tree_add_51_79_groupi_n_7265);
  or csa_tree_add_51_79_groupi_g38314(csa_tree_add_51_79_groupi_n_7749 ,csa_tree_add_51_79_groupi_n_7227 ,csa_tree_add_51_79_groupi_n_7264);
  and csa_tree_add_51_79_groupi_g38315(csa_tree_add_51_79_groupi_n_7748 ,csa_tree_add_51_79_groupi_n_7227 ,csa_tree_add_51_79_groupi_n_7264);
  or csa_tree_add_51_79_groupi_g38316(csa_tree_add_51_79_groupi_n_7747 ,csa_tree_add_51_79_groupi_n_7309 ,csa_tree_add_51_79_groupi_n_7260);
  and csa_tree_add_51_79_groupi_g38317(csa_tree_add_51_79_groupi_n_7746 ,csa_tree_add_51_79_groupi_n_7309 ,csa_tree_add_51_79_groupi_n_7260);
  and csa_tree_add_51_79_groupi_g38318(csa_tree_add_51_79_groupi_n_7745 ,csa_tree_add_51_79_groupi_n_7305 ,csa_tree_add_51_79_groupi_n_7259);
  or csa_tree_add_51_79_groupi_g38319(csa_tree_add_51_79_groupi_n_7744 ,csa_tree_add_51_79_groupi_n_7305 ,csa_tree_add_51_79_groupi_n_7259);
  and csa_tree_add_51_79_groupi_g38320(csa_tree_add_51_79_groupi_n_7743 ,csa_tree_add_51_79_groupi_n_7299 ,csa_tree_add_51_79_groupi_n_7298);
  or csa_tree_add_51_79_groupi_g38321(csa_tree_add_51_79_groupi_n_7742 ,csa_tree_add_51_79_groupi_n_7241 ,csa_tree_add_51_79_groupi_n_7297);
  and csa_tree_add_51_79_groupi_g38322(csa_tree_add_51_79_groupi_n_7741 ,csa_tree_add_51_79_groupi_n_7241 ,csa_tree_add_51_79_groupi_n_7297);
  or csa_tree_add_51_79_groupi_g38323(csa_tree_add_51_79_groupi_n_7740 ,csa_tree_add_51_79_groupi_n_7295 ,csa_tree_add_51_79_groupi_n_7294);
  or csa_tree_add_51_79_groupi_g38324(csa_tree_add_51_79_groupi_n_7739 ,csa_tree_add_51_79_groupi_n_7299 ,csa_tree_add_51_79_groupi_n_7298);
  or csa_tree_add_51_79_groupi_g38325(csa_tree_add_51_79_groupi_n_7738 ,csa_tree_add_51_79_groupi_n_7285 ,csa_tree_add_51_79_groupi_n_7281);
  and csa_tree_add_51_79_groupi_g38326(csa_tree_add_51_79_groupi_n_7737 ,csa_tree_add_51_79_groupi_n_7285 ,csa_tree_add_51_79_groupi_n_7281);
  or csa_tree_add_51_79_groupi_g38327(csa_tree_add_51_79_groupi_n_7736 ,csa_tree_add_51_79_groupi_n_7075 ,csa_tree_add_51_79_groupi_n_7449);
  or csa_tree_add_51_79_groupi_g38328(csa_tree_add_51_79_groupi_n_7735 ,csa_tree_add_51_79_groupi_n_6148 ,csa_tree_add_51_79_groupi_n_7398);
  or csa_tree_add_51_79_groupi_g38329(csa_tree_add_51_79_groupi_n_7734 ,csa_tree_add_51_79_groupi_n_5867 ,csa_tree_add_51_79_groupi_n_7495);
  or csa_tree_add_51_79_groupi_g38330(csa_tree_add_51_79_groupi_n_7733 ,csa_tree_add_51_79_groupi_n_6154 ,csa_tree_add_51_79_groupi_n_7391);
  or csa_tree_add_51_79_groupi_g38331(csa_tree_add_51_79_groupi_n_7732 ,csa_tree_add_51_79_groupi_n_5868 ,csa_tree_add_51_79_groupi_n_7442);
  or csa_tree_add_51_79_groupi_g38332(csa_tree_add_51_79_groupi_n_7731 ,csa_tree_add_51_79_groupi_n_7097 ,csa_tree_add_51_79_groupi_n_7389);
  or csa_tree_add_51_79_groupi_g38333(csa_tree_add_51_79_groupi_n_7730 ,csa_tree_add_51_79_groupi_n_7063 ,csa_tree_add_51_79_groupi_n_7464);
  or csa_tree_add_51_79_groupi_g38334(csa_tree_add_51_79_groupi_n_7729 ,csa_tree_add_51_79_groupi_n_6939 ,csa_tree_add_51_79_groupi_n_7524);
  or csa_tree_add_51_79_groupi_g38335(csa_tree_add_51_79_groupi_n_7728 ,csa_tree_add_51_79_groupi_n_7313 ,csa_tree_add_51_79_groupi_n_7315);
  or csa_tree_add_51_79_groupi_g38336(csa_tree_add_51_79_groupi_n_7727 ,csa_tree_add_51_79_groupi_n_7262 ,csa_tree_add_51_79_groupi_n_7144);
  nor csa_tree_add_51_79_groupi_g38337(csa_tree_add_51_79_groupi_n_7726 ,csa_tree_add_51_79_groupi_n_7261 ,csa_tree_add_51_79_groupi_n_7145);
  nor csa_tree_add_51_79_groupi_g38338(csa_tree_add_51_79_groupi_n_7725 ,csa_tree_add_51_79_groupi_n_7312 ,csa_tree_add_51_79_groupi_n_7316);
  or csa_tree_add_51_79_groupi_g38339(csa_tree_add_51_79_groupi_n_7724 ,csa_tree_add_51_79_groupi_n_6779 ,csa_tree_add_51_79_groupi_n_7364);
  or csa_tree_add_51_79_groupi_g38340(csa_tree_add_51_79_groupi_n_7723 ,csa_tree_add_51_79_groupi_n_6921 ,csa_tree_add_51_79_groupi_n_7395);
  and csa_tree_add_51_79_groupi_g38341(csa_tree_add_51_79_groupi_n_7722 ,csa_tree_add_51_79_groupi_n_7152 ,csa_tree_add_51_79_groupi_n_7151);
  xnor csa_tree_add_51_79_groupi_g38342(csa_tree_add_51_79_groupi_n_7721 ,csa_tree_add_51_79_groupi_n_6869 ,csa_tree_add_51_79_groupi_n_6997);
  xnor csa_tree_add_51_79_groupi_g38343(csa_tree_add_51_79_groupi_n_7720 ,csa_tree_add_51_79_groupi_n_7026 ,csa_tree_add_51_79_groupi_n_7117);
  xnor csa_tree_add_51_79_groupi_g38344(csa_tree_add_51_79_groupi_n_7719 ,csa_tree_add_51_79_groupi_n_6908 ,csa_tree_add_51_79_groupi_n_6856);
  xnor csa_tree_add_51_79_groupi_g38345(csa_tree_add_51_79_groupi_n_7718 ,csa_tree_add_51_79_groupi_n_7076 ,csa_tree_add_51_79_groupi_n_6998);
  xnor csa_tree_add_51_79_groupi_g38346(csa_tree_add_51_79_groupi_n_7717 ,csa_tree_add_51_79_groupi_n_7081 ,csa_tree_add_51_79_groupi_n_7010);
  xnor csa_tree_add_51_79_groupi_g38347(csa_tree_add_51_79_groupi_n_7716 ,csa_tree_add_51_79_groupi_n_6992 ,csa_tree_add_51_79_groupi_n_7062);
  xnor csa_tree_add_51_79_groupi_g38348(csa_tree_add_51_79_groupi_n_7715 ,csa_tree_add_51_79_groupi_n_6994 ,csa_tree_add_51_79_groupi_n_7004);
  xnor csa_tree_add_51_79_groupi_g38349(csa_tree_add_51_79_groupi_n_7714 ,csa_tree_add_51_79_groupi_n_6970 ,csa_tree_add_51_79_groupi_n_6978);
  xnor csa_tree_add_51_79_groupi_g38350(csa_tree_add_51_79_groupi_n_7713 ,csa_tree_add_51_79_groupi_n_6821 ,csa_tree_add_51_79_groupi_n_6865);
  xnor csa_tree_add_51_79_groupi_g38351(csa_tree_add_51_79_groupi_n_7712 ,csa_tree_add_51_79_groupi_n_6901 ,csa_tree_add_51_79_groupi_n_6879);
  xnor csa_tree_add_51_79_groupi_g38352(csa_tree_add_51_79_groupi_n_7711 ,csa_tree_add_51_79_groupi_n_7099 ,csa_tree_add_51_79_groupi_n_7051);
  xnor csa_tree_add_51_79_groupi_g38353(csa_tree_add_51_79_groupi_n_7710 ,csa_tree_add_51_79_groupi_n_5841 ,csa_tree_add_51_79_groupi_n_6926);
  xnor csa_tree_add_51_79_groupi_g38354(csa_tree_add_51_79_groupi_n_7709 ,csa_tree_add_51_79_groupi_n_6740 ,csa_tree_add_51_79_groupi_n_6981);
  xnor csa_tree_add_51_79_groupi_g38355(csa_tree_add_51_79_groupi_n_7708 ,csa_tree_add_51_79_groupi_n_6823 ,csa_tree_add_51_79_groupi_n_6920);
  xnor csa_tree_add_51_79_groupi_g38356(csa_tree_add_51_79_groupi_n_7707 ,csa_tree_add_51_79_groupi_n_5309 ,csa_tree_add_51_79_groupi_n_7083);
  xnor csa_tree_add_51_79_groupi_g38357(csa_tree_add_51_79_groupi_n_7706 ,csa_tree_add_51_79_groupi_n_6974 ,csa_tree_add_51_79_groupi_n_6909);
  xnor csa_tree_add_51_79_groupi_g38358(csa_tree_add_51_79_groupi_n_7705 ,csa_tree_add_51_79_groupi_n_6929 ,csa_tree_add_51_79_groupi_n_6825);
  xnor csa_tree_add_51_79_groupi_g38359(csa_tree_add_51_79_groupi_n_7704 ,csa_tree_add_51_79_groupi_n_6867 ,csa_tree_add_51_79_groupi_n_6988);
  xnor csa_tree_add_51_79_groupi_g38360(csa_tree_add_51_79_groupi_n_7703 ,csa_tree_add_51_79_groupi_n_7020 ,csa_tree_add_51_79_groupi_n_6973);
  xnor csa_tree_add_51_79_groupi_g38361(csa_tree_add_51_79_groupi_n_7702 ,csa_tree_add_51_79_groupi_n_6918 ,csa_tree_add_51_79_groupi_n_6728);
  xnor csa_tree_add_51_79_groupi_g38362(csa_tree_add_51_79_groupi_n_7701 ,csa_tree_add_51_79_groupi_n_6982 ,csa_tree_add_51_79_groupi_n_6983);
  xnor csa_tree_add_51_79_groupi_g38363(csa_tree_add_51_79_groupi_n_7700 ,csa_tree_add_51_79_groupi_n_6979 ,csa_tree_add_51_79_groupi_n_6746);
  xnor csa_tree_add_51_79_groupi_g38364(csa_tree_add_51_79_groupi_n_7699 ,csa_tree_add_51_79_groupi_n_7042 ,csa_tree_add_51_79_groupi_n_7095);
  xnor csa_tree_add_51_79_groupi_g38365(csa_tree_add_51_79_groupi_n_7698 ,csa_tree_add_51_79_groupi_n_6853 ,csa_tree_add_51_79_groupi_n_7084);
  xnor csa_tree_add_51_79_groupi_g38366(csa_tree_add_51_79_groupi_n_7697 ,csa_tree_add_51_79_groupi_n_7003 ,csa_tree_add_51_79_groupi_n_7036);
  xnor csa_tree_add_51_79_groupi_g38367(csa_tree_add_51_79_groupi_n_7696 ,csa_tree_add_51_79_groupi_n_7021 ,csa_tree_add_51_79_groupi_n_7033);
  xnor csa_tree_add_51_79_groupi_g38368(csa_tree_add_51_79_groupi_n_7695 ,csa_tree_add_51_79_groupi_n_7107 ,csa_tree_add_51_79_groupi_n_6742);
  xnor csa_tree_add_51_79_groupi_g38369(csa_tree_add_51_79_groupi_n_7694 ,csa_tree_add_51_79_groupi_n_6845 ,csa_tree_add_51_79_groupi_n_6844);
  xnor csa_tree_add_51_79_groupi_g38370(csa_tree_add_51_79_groupi_n_7693 ,csa_tree_add_51_79_groupi_n_6154 ,csa_tree_add_51_79_groupi_n_6847);
  xnor csa_tree_add_51_79_groupi_g38371(csa_tree_add_51_79_groupi_n_7692 ,csa_tree_add_51_79_groupi_n_5853 ,csa_tree_add_51_79_groupi_n_6888);
  xnor csa_tree_add_51_79_groupi_g38372(csa_tree_add_51_79_groupi_n_7691 ,csa_tree_add_51_79_groupi_n_6841 ,csa_tree_add_51_79_groupi_n_6837);
  xnor csa_tree_add_51_79_groupi_g38373(csa_tree_add_51_79_groupi_n_7690 ,csa_tree_add_51_79_groupi_n_5868 ,csa_tree_add_51_79_groupi_n_6838);
  xnor csa_tree_add_51_79_groupi_g38374(csa_tree_add_51_79_groupi_n_7689 ,csa_tree_add_51_79_groupi_n_5867 ,csa_tree_add_51_79_groupi_n_6843);
  xnor csa_tree_add_51_79_groupi_g38375(csa_tree_add_51_79_groupi_n_7688 ,csa_tree_add_51_79_groupi_n_6848 ,csa_tree_add_51_79_groupi_n_6835);
  xor csa_tree_add_51_79_groupi_g38376(csa_tree_add_51_79_groupi_n_7687 ,csa_tree_add_51_79_groupi_n_7114 ,csa_tree_add_51_79_groupi_n_6820);
  xnor csa_tree_add_51_79_groupi_g38379(csa_tree_add_51_79_groupi_n_7686 ,csa_tree_add_51_79_groupi_n_7093 ,csa_tree_add_51_79_groupi_n_6743);
  xnor csa_tree_add_51_79_groupi_g38380(csa_tree_add_51_79_groupi_n_7685 ,csa_tree_add_51_79_groupi_n_6832 ,csa_tree_add_51_79_groupi_n_6148);
  xnor csa_tree_add_51_79_groupi_g38381(csa_tree_add_51_79_groupi_n_7684 ,csa_tree_add_51_79_groupi_n_6829 ,csa_tree_add_51_79_groupi_n_6830);
  xnor csa_tree_add_51_79_groupi_g38382(csa_tree_add_51_79_groupi_n_7683 ,csa_tree_add_51_79_groupi_n_6977 ,csa_tree_add_51_79_groupi_n_7072);
  xnor csa_tree_add_51_79_groupi_g38383(csa_tree_add_51_79_groupi_n_7682 ,csa_tree_add_51_79_groupi_n_6882 ,csa_tree_add_51_79_groupi_n_6891);
  xnor csa_tree_add_51_79_groupi_g38384(csa_tree_add_51_79_groupi_n_7681 ,csa_tree_add_51_79_groupi_n_6933 ,csa_tree_add_51_79_groupi_n_6824);
  xnor csa_tree_add_51_79_groupi_g38385(csa_tree_add_51_79_groupi_n_7680 ,csa_tree_add_51_79_groupi_n_6927 ,csa_tree_add_51_79_groupi_n_6859);
  xnor csa_tree_add_51_79_groupi_g38386(csa_tree_add_51_79_groupi_n_7679 ,csa_tree_add_51_79_groupi_n_7048 ,csa_tree_add_51_79_groupi_n_7053);
  xnor csa_tree_add_51_79_groupi_g38387(csa_tree_add_51_79_groupi_n_7678 ,csa_tree_add_51_79_groupi_n_6966 ,csa_tree_add_51_79_groupi_n_7088);
  xnor csa_tree_add_51_79_groupi_g38388(csa_tree_add_51_79_groupi_n_7677 ,csa_tree_add_51_79_groupi_n_7059 ,csa_tree_add_51_79_groupi_n_7060);
  xnor csa_tree_add_51_79_groupi_g38389(csa_tree_add_51_79_groupi_n_7676 ,csa_tree_add_51_79_groupi_n_6826 ,csa_tree_add_51_79_groupi_n_6880);
  xnor csa_tree_add_51_79_groupi_g38390(csa_tree_add_51_79_groupi_n_7675 ,csa_tree_add_51_79_groupi_n_7043 ,csa_tree_add_51_79_groupi_n_7044);
  xnor csa_tree_add_51_79_groupi_g38391(csa_tree_add_51_79_groupi_n_7674 ,csa_tree_add_51_79_groupi_n_7090 ,csa_tree_add_51_79_groupi_n_7022);
  xnor csa_tree_add_51_79_groupi_g38392(csa_tree_add_51_79_groupi_n_7673 ,csa_tree_add_51_79_groupi_n_6919 ,csa_tree_add_51_79_groupi_n_6755);
  xnor csa_tree_add_51_79_groupi_g38393(csa_tree_add_51_79_groupi_n_7672 ,csa_tree_add_51_79_groupi_n_6968 ,csa_tree_add_51_79_groupi_n_7068);
  xnor csa_tree_add_51_79_groupi_g38394(csa_tree_add_51_79_groupi_n_7671 ,csa_tree_add_51_79_groupi_n_6916 ,csa_tree_add_51_79_groupi_n_6881);
  xnor csa_tree_add_51_79_groupi_g38395(csa_tree_add_51_79_groupi_n_7670 ,csa_tree_add_51_79_groupi_n_6886 ,csa_tree_add_51_79_groupi_n_6842);
  xnor csa_tree_add_51_79_groupi_g38396(csa_tree_add_51_79_groupi_n_7669 ,csa_tree_add_51_79_groupi_n_6871 ,csa_tree_add_51_79_groupi_n_7091);
  xnor csa_tree_add_51_79_groupi_g38397(csa_tree_add_51_79_groupi_n_7668 ,csa_tree_add_51_79_groupi_n_7013 ,csa_tree_add_51_79_groupi_n_7054);
  xnor csa_tree_add_51_79_groupi_g38398(csa_tree_add_51_79_groupi_n_7667 ,csa_tree_add_51_79_groupi_n_6864 ,csa_tree_add_51_79_groupi_n_6911);
  xnor csa_tree_add_51_79_groupi_g38399(csa_tree_add_51_79_groupi_n_7666 ,csa_tree_add_51_79_groupi_n_6851 ,csa_tree_add_51_79_groupi_n_6840);
  xnor csa_tree_add_51_79_groupi_g38400(csa_tree_add_51_79_groupi_n_7665 ,csa_tree_add_51_79_groupi_n_6995 ,csa_tree_add_51_79_groupi_n_6999);
  xnor csa_tree_add_51_79_groupi_g38401(csa_tree_add_51_79_groupi_n_7664 ,csa_tree_add_51_79_groupi_n_7061 ,csa_tree_add_51_79_groupi_n_7077);
  xnor csa_tree_add_51_79_groupi_g38402(csa_tree_add_51_79_groupi_n_7663 ,csa_tree_add_51_79_groupi_n_7006 ,csa_tree_add_51_79_groupi_n_7018);
  xnor csa_tree_add_51_79_groupi_g38403(csa_tree_add_51_79_groupi_n_7662 ,csa_tree_add_51_79_groupi_n_6975 ,csa_tree_add_51_79_groupi_n_7110);
  xor csa_tree_add_51_79_groupi_g38404(csa_tree_add_51_79_groupi_n_7661 ,csa_tree_add_51_79_groupi_n_6903 ,csa_tree_add_51_79_groupi_n_7000);
  xnor csa_tree_add_51_79_groupi_g38405(csa_tree_add_51_79_groupi_n_7660 ,csa_tree_add_51_79_groupi_n_7106 ,csa_tree_add_51_79_groupi_n_7056);
  xnor csa_tree_add_51_79_groupi_g38406(csa_tree_add_51_79_groupi_n_7659 ,csa_tree_add_51_79_groupi_n_7034 ,csa_tree_add_51_79_groupi_n_7037);
  xnor csa_tree_add_51_79_groupi_g38407(csa_tree_add_51_79_groupi_n_7658 ,csa_tree_add_51_79_groupi_n_7082 ,csa_tree_add_51_79_groupi_n_6432);
  xnor csa_tree_add_51_79_groupi_g38408(csa_tree_add_51_79_groupi_n_7657 ,csa_tree_add_51_79_groupi_n_7086 ,csa_tree_add_51_79_groupi_n_7016);
  xnor csa_tree_add_51_79_groupi_g38409(csa_tree_add_51_79_groupi_n_7656 ,csa_tree_add_51_79_groupi_n_6873 ,csa_tree_add_51_79_groupi_n_6914);
  xnor csa_tree_add_51_79_groupi_g38410(csa_tree_add_51_79_groupi_n_7655 ,csa_tree_add_51_79_groupi_n_6816 ,csa_tree_add_51_79_groupi_n_6925);
  xnor csa_tree_add_51_79_groupi_g38411(csa_tree_add_51_79_groupi_n_7654 ,csa_tree_add_51_79_groupi_n_6893 ,csa_tree_add_51_79_groupi_n_6937);
  xnor csa_tree_add_51_79_groupi_g38412(csa_tree_add_51_79_groupi_n_7653 ,csa_tree_add_51_79_groupi_n_6889 ,csa_tree_add_51_79_groupi_n_6892);
  xnor csa_tree_add_51_79_groupi_g38413(csa_tree_add_51_79_groupi_n_7652 ,csa_tree_add_51_79_groupi_n_7023 ,csa_tree_add_51_79_groupi_n_7038);
  xnor csa_tree_add_51_79_groupi_g38414(csa_tree_add_51_79_groupi_n_7651 ,csa_tree_add_51_79_groupi_n_6874 ,csa_tree_add_51_79_groupi_n_6928);
  xnor csa_tree_add_51_79_groupi_g38415(csa_tree_add_51_79_groupi_n_7650 ,csa_tree_add_51_79_groupi_n_6817 ,csa_tree_add_51_79_groupi_n_6962);
  xnor csa_tree_add_51_79_groupi_g38416(csa_tree_add_51_79_groupi_n_7649 ,csa_tree_add_51_79_groupi_n_7092 ,csa_tree_add_51_79_groupi_n_7031);
  xnor csa_tree_add_51_79_groupi_g38417(csa_tree_add_51_79_groupi_n_7648 ,csa_tree_add_51_79_groupi_n_7080 ,csa_tree_add_51_79_groupi_n_7005);
  xnor csa_tree_add_51_79_groupi_g38418(csa_tree_add_51_79_groupi_n_7647 ,csa_tree_add_51_79_groupi_n_7049 ,csa_tree_add_51_79_groupi_n_7100);
  xnor csa_tree_add_51_79_groupi_g38419(csa_tree_add_51_79_groupi_n_7646 ,csa_tree_add_51_79_groupi_n_7057 ,csa_tree_add_51_79_groupi_n_7058);
  xnor csa_tree_add_51_79_groupi_g38420(csa_tree_add_51_79_groupi_n_7645 ,csa_tree_add_51_79_groupi_n_6932 ,csa_tree_add_51_79_groupi_n_6898);
  xnor csa_tree_add_51_79_groupi_g38421(csa_tree_add_51_79_groupi_n_7644 ,csa_tree_add_51_79_groupi_n_6885 ,csa_tree_add_51_79_groupi_n_6915);
  xnor csa_tree_add_51_79_groupi_g38422(csa_tree_add_51_79_groupi_n_7643 ,csa_tree_add_51_79_groupi_n_6936 ,csa_tree_add_51_79_groupi_n_7029);
  xnor csa_tree_add_51_79_groupi_g38423(csa_tree_add_51_79_groupi_n_7642 ,csa_tree_add_51_79_groupi_n_6985 ,csa_tree_add_51_79_groupi_n_7104);
  xnor csa_tree_add_51_79_groupi_g38424(csa_tree_add_51_79_groupi_n_7641 ,csa_tree_add_51_79_groupi_n_6967 ,csa_tree_add_51_79_groupi_n_6972);
  xnor csa_tree_add_51_79_groupi_g38425(csa_tree_add_51_79_groupi_n_7640 ,csa_tree_add_51_79_groupi_n_6964 ,csa_tree_add_51_79_groupi_n_7108);
  xnor csa_tree_add_51_79_groupi_g38426(csa_tree_add_51_79_groupi_n_7639 ,csa_tree_add_51_79_groupi_n_7111 ,csa_tree_add_51_79_groupi_n_6989);
  xnor csa_tree_add_51_79_groupi_g38427(csa_tree_add_51_79_groupi_n_7638 ,csa_tree_add_51_79_groupi_n_7116 ,csa_tree_add_51_79_groupi_n_7028);
  xnor csa_tree_add_51_79_groupi_g38428(csa_tree_add_51_79_groupi_n_7637 ,csa_tree_add_51_79_groupi_n_7078 ,csa_tree_add_51_79_groupi_n_7012);
  xnor csa_tree_add_51_79_groupi_g38429(csa_tree_add_51_79_groupi_n_7636 ,csa_tree_add_51_79_groupi_n_7015 ,csa_tree_add_51_79_groupi_n_7019);
  xnor csa_tree_add_51_79_groupi_g38430(csa_tree_add_51_79_groupi_n_7833 ,csa_tree_add_51_79_groupi_n_6451 ,csa_tree_add_51_79_groupi_n_6776);
  and csa_tree_add_51_79_groupi_g38431(csa_tree_add_51_79_groupi_n_7832 ,csa_tree_add_51_79_groupi_n_6794 ,csa_tree_add_51_79_groupi_n_7402);
  and csa_tree_add_51_79_groupi_g38432(csa_tree_add_51_79_groupi_n_7831 ,csa_tree_add_51_79_groupi_n_6801 ,csa_tree_add_51_79_groupi_n_7401);
  xnor csa_tree_add_51_79_groupi_g38433(csa_tree_add_51_79_groupi_n_7830 ,csa_tree_add_51_79_groupi_n_6452 ,csa_tree_add_51_79_groupi_n_6768);
  xnor csa_tree_add_51_79_groupi_g38434(csa_tree_add_51_79_groupi_n_7829 ,csa_tree_add_51_79_groupi_n_6149 ,csa_tree_add_51_79_groupi_n_6765);
  and csa_tree_add_51_79_groupi_g38435(csa_tree_add_51_79_groupi_n_7828 ,csa_tree_add_51_79_groupi_n_6804 ,csa_tree_add_51_79_groupi_n_7393);
  and csa_tree_add_51_79_groupi_g38436(csa_tree_add_51_79_groupi_n_7827 ,csa_tree_add_51_79_groupi_n_6812 ,csa_tree_add_51_79_groupi_n_7491);
  xnor csa_tree_add_51_79_groupi_g38437(csa_tree_add_51_79_groupi_n_7826 ,csa_tree_add_51_79_groupi_n_6144 ,csa_tree_add_51_79_groupi_n_6763);
  xnor csa_tree_add_51_79_groupi_g38438(csa_tree_add_51_79_groupi_n_7825 ,csa_tree_add_51_79_groupi_n_6445 ,csa_tree_add_51_79_groupi_n_6770);
  xnor csa_tree_add_51_79_groupi_g38439(csa_tree_add_51_79_groupi_n_7823 ,csa_tree_add_51_79_groupi_n_25 ,csa_tree_add_51_79_groupi_n_6771);
  xnor csa_tree_add_51_79_groupi_g38440(csa_tree_add_51_79_groupi_n_7822 ,csa_tree_add_51_79_groupi_n_6156 ,csa_tree_add_51_79_groupi_n_6775);
  xnor csa_tree_add_51_79_groupi_g38441(csa_tree_add_51_79_groupi_n_7820 ,csa_tree_add_51_79_groupi_n_6913 ,csa_tree_add_51_79_groupi_n_6772);
  xnor csa_tree_add_51_79_groupi_g38442(csa_tree_add_51_79_groupi_n_7819 ,csa_tree_add_51_79_groupi_n_7101 ,csa_tree_add_51_79_groupi_n_6774);
  and csa_tree_add_51_79_groupi_g38443(csa_tree_add_51_79_groupi_n_7817 ,csa_tree_add_51_79_groupi_n_6808 ,csa_tree_add_51_79_groupi_n_7465);
  xnor csa_tree_add_51_79_groupi_g38444(csa_tree_add_51_79_groupi_n_7816 ,csa_tree_add_51_79_groupi_n_5846 ,csa_tree_add_51_79_groupi_n_6764);
  and csa_tree_add_51_79_groupi_g38445(csa_tree_add_51_79_groupi_n_7815 ,csa_tree_add_51_79_groupi_n_6806 ,csa_tree_add_51_79_groupi_n_7413);
  xnor csa_tree_add_51_79_groupi_g38446(csa_tree_add_51_79_groupi_n_7813 ,csa_tree_add_51_79_groupi_n_6422 ,csa_tree_add_51_79_groupi_n_6773);
  or csa_tree_add_51_79_groupi_g38447(csa_tree_add_51_79_groupi_n_7811 ,csa_tree_add_51_79_groupi_n_6942 ,csa_tree_add_51_79_groupi_n_7394);
  xnor csa_tree_add_51_79_groupi_g38448(csa_tree_add_51_79_groupi_n_7810 ,csa_tree_add_51_79_groupi_n_5863 ,csa_tree_add_51_79_groupi_n_6777);
  and csa_tree_add_51_79_groupi_g38449(csa_tree_add_51_79_groupi_n_7808 ,csa_tree_add_51_79_groupi_n_6802 ,csa_tree_add_51_79_groupi_n_7400);
  xnor csa_tree_add_51_79_groupi_g38450(csa_tree_add_51_79_groupi_n_7807 ,csa_tree_add_51_79_groupi_n_6129 ,csa_tree_add_51_79_groupi_n_6766);
  and csa_tree_add_51_79_groupi_g38451(csa_tree_add_51_79_groupi_n_7806 ,csa_tree_add_51_79_groupi_n_6799 ,csa_tree_add_51_79_groupi_n_7403);
  xnor csa_tree_add_51_79_groupi_g38452(csa_tree_add_51_79_groupi_n_7805 ,csa_tree_add_51_79_groupi_n_6137 ,csa_tree_add_51_79_groupi_n_6767);
  and csa_tree_add_51_79_groupi_g38453(csa_tree_add_51_79_groupi_n_7804 ,csa_tree_add_51_79_groupi_n_6791 ,csa_tree_add_51_79_groupi_n_7404);
  xnor csa_tree_add_51_79_groupi_g38454(csa_tree_add_51_79_groupi_n_7803 ,csa_tree_add_51_79_groupi_n_5848 ,csa_tree_add_51_79_groupi_n_6769);
  not csa_tree_add_51_79_groupi_g38455(csa_tree_add_51_79_groupi_n_7632 ,csa_tree_add_51_79_groupi_n_7631);
  not csa_tree_add_51_79_groupi_g38456(csa_tree_add_51_79_groupi_n_7622 ,csa_tree_add_51_79_groupi_n_7621);
  not csa_tree_add_51_79_groupi_g38457(csa_tree_add_51_79_groupi_n_7620 ,csa_tree_add_51_79_groupi_n_7619);
  not csa_tree_add_51_79_groupi_g38458(csa_tree_add_51_79_groupi_n_7615 ,csa_tree_add_51_79_groupi_n_7616);
  not csa_tree_add_51_79_groupi_g38459(csa_tree_add_51_79_groupi_n_7613 ,csa_tree_add_51_79_groupi_n_7614);
  not csa_tree_add_51_79_groupi_g38460(csa_tree_add_51_79_groupi_n_7612 ,csa_tree_add_51_79_groupi_n_7611);
  not csa_tree_add_51_79_groupi_g38461(csa_tree_add_51_79_groupi_n_7608 ,csa_tree_add_51_79_groupi_n_7609);
  not csa_tree_add_51_79_groupi_g38462(csa_tree_add_51_79_groupi_n_7606 ,csa_tree_add_51_79_groupi_n_7607);
  not csa_tree_add_51_79_groupi_g38463(csa_tree_add_51_79_groupi_n_7604 ,csa_tree_add_51_79_groupi_n_7605);
  not csa_tree_add_51_79_groupi_g38464(csa_tree_add_51_79_groupi_n_7602 ,csa_tree_add_51_79_groupi_n_7603);
  not csa_tree_add_51_79_groupi_g38466(csa_tree_add_51_79_groupi_n_7597 ,csa_tree_add_51_79_groupi_n_7598);
  not csa_tree_add_51_79_groupi_g38467(csa_tree_add_51_79_groupi_n_7594 ,csa_tree_add_51_79_groupi_n_7595);
  not csa_tree_add_51_79_groupi_g38468(csa_tree_add_51_79_groupi_n_7591 ,csa_tree_add_51_79_groupi_n_7592);
  not csa_tree_add_51_79_groupi_g38469(csa_tree_add_51_79_groupi_n_7590 ,csa_tree_add_51_79_groupi_n_10);
  not csa_tree_add_51_79_groupi_g38470(csa_tree_add_51_79_groupi_n_7588 ,csa_tree_add_51_79_groupi_n_7589);
  not csa_tree_add_51_79_groupi_g38471(csa_tree_add_51_79_groupi_n_7586 ,csa_tree_add_51_79_groupi_n_7587);
  not csa_tree_add_51_79_groupi_g38472(csa_tree_add_51_79_groupi_n_7584 ,csa_tree_add_51_79_groupi_n_7585);
  not csa_tree_add_51_79_groupi_g38473(csa_tree_add_51_79_groupi_n_7581 ,csa_tree_add_51_79_groupi_n_7582);
  not csa_tree_add_51_79_groupi_g38474(csa_tree_add_51_79_groupi_n_7579 ,csa_tree_add_51_79_groupi_n_7580);
  not csa_tree_add_51_79_groupi_g38475(csa_tree_add_51_79_groupi_n_7577 ,csa_tree_add_51_79_groupi_n_7578);
  and csa_tree_add_51_79_groupi_g38476(csa_tree_add_51_79_groupi_n_7575 ,csa_tree_add_51_79_groupi_n_6840 ,csa_tree_add_51_79_groupi_n_6851);
  nor csa_tree_add_51_79_groupi_g38477(csa_tree_add_51_79_groupi_n_7574 ,csa_tree_add_51_79_groupi_n_6823 ,csa_tree_add_51_79_groupi_n_6897);
  or csa_tree_add_51_79_groupi_g38478(csa_tree_add_51_79_groupi_n_7573 ,csa_tree_add_51_79_groupi_n_6495 ,csa_tree_add_51_79_groupi_n_7101);
  or csa_tree_add_51_79_groupi_g38479(csa_tree_add_51_79_groupi_n_7572 ,csa_tree_add_51_79_groupi_n_6973 ,csa_tree_add_51_79_groupi_n_7020);
  nor csa_tree_add_51_79_groupi_g38480(csa_tree_add_51_79_groupi_n_7571 ,csa_tree_add_51_79_groupi_n_6128 ,csa_tree_add_51_79_groupi_n_7000);
  or csa_tree_add_51_79_groupi_g38481(csa_tree_add_51_79_groupi_n_7570 ,csa_tree_add_51_79_groupi_n_7019 ,csa_tree_add_51_79_groupi_n_7015);
  nor csa_tree_add_51_79_groupi_g38482(csa_tree_add_51_79_groupi_n_7569 ,csa_tree_add_51_79_groupi_n_7003 ,csa_tree_add_51_79_groupi_n_7035);
  and csa_tree_add_51_79_groupi_g38483(csa_tree_add_51_79_groupi_n_7568 ,csa_tree_add_51_79_groupi_n_7019 ,csa_tree_add_51_79_groupi_n_7015);
  or csa_tree_add_51_79_groupi_g38484(csa_tree_add_51_79_groupi_n_7567 ,csa_tree_add_51_79_groupi_n_7061 ,csa_tree_add_51_79_groupi_n_7047);
  or csa_tree_add_51_79_groupi_g38485(csa_tree_add_51_79_groupi_n_7566 ,csa_tree_add_51_79_groupi_n_7053 ,csa_tree_add_51_79_groupi_n_7048);
  and csa_tree_add_51_79_groupi_g38486(csa_tree_add_51_79_groupi_n_7565 ,csa_tree_add_51_79_groupi_n_6973 ,csa_tree_add_51_79_groupi_n_7020);
  and csa_tree_add_51_79_groupi_g38487(csa_tree_add_51_79_groupi_n_7564 ,csa_tree_add_51_79_groupi_n_7053 ,csa_tree_add_51_79_groupi_n_7048);
  and csa_tree_add_51_79_groupi_g38488(csa_tree_add_51_79_groupi_n_7563 ,csa_tree_add_51_79_groupi_n_7061 ,csa_tree_add_51_79_groupi_n_7047);
  or csa_tree_add_51_79_groupi_g38489(csa_tree_add_51_79_groupi_n_7562 ,csa_tree_add_51_79_groupi_n_6130 ,csa_tree_add_51_79_groupi_n_7012);
  or csa_tree_add_51_79_groupi_g38490(csa_tree_add_51_79_groupi_n_7561 ,csa_tree_add_51_79_groupi_n_6153 ,csa_tree_add_51_79_groupi_n_6948);
  or csa_tree_add_51_79_groupi_g38491(csa_tree_add_51_79_groupi_n_7560 ,csa_tree_add_51_79_groupi_n_7005 ,csa_tree_add_51_79_groupi_n_6993);
  nor csa_tree_add_51_79_groupi_g38492(csa_tree_add_51_79_groupi_n_7559 ,csa_tree_add_51_79_groupi_n_6131 ,csa_tree_add_51_79_groupi_n_7011);
  and csa_tree_add_51_79_groupi_g38493(csa_tree_add_51_79_groupi_n_7558 ,csa_tree_add_51_79_groupi_n_7005 ,csa_tree_add_51_79_groupi_n_6993);
  or csa_tree_add_51_79_groupi_g38494(csa_tree_add_51_79_groupi_n_7557 ,csa_tree_add_51_79_groupi_n_6966 ,csa_tree_add_51_79_groupi_n_6963);
  or csa_tree_add_51_79_groupi_g38495(csa_tree_add_51_79_groupi_n_7556 ,csa_tree_add_51_79_groupi_n_6744 ,csa_tree_add_51_79_groupi_n_7056);
  and csa_tree_add_51_79_groupi_g38496(csa_tree_add_51_79_groupi_n_7555 ,csa_tree_add_51_79_groupi_n_6966 ,csa_tree_add_51_79_groupi_n_6963);
  or csa_tree_add_51_79_groupi_g38497(csa_tree_add_51_79_groupi_n_7554 ,csa_tree_add_51_79_groupi_n_7058 ,csa_tree_add_51_79_groupi_n_7057);
  and csa_tree_add_51_79_groupi_g38498(csa_tree_add_51_79_groupi_n_7553 ,csa_tree_add_51_79_groupi_n_7058 ,csa_tree_add_51_79_groupi_n_7057);
  or csa_tree_add_51_79_groupi_g38499(csa_tree_add_51_79_groupi_n_7552 ,csa_tree_add_51_79_groupi_n_7050 ,csa_tree_add_51_79_groupi_n_7049);
  and csa_tree_add_51_79_groupi_g38500(csa_tree_add_51_79_groupi_n_7551 ,csa_tree_add_51_79_groupi_n_7050 ,csa_tree_add_51_79_groupi_n_7049);
  nor csa_tree_add_51_79_groupi_g38501(csa_tree_add_51_79_groupi_n_7550 ,csa_tree_add_51_79_groupi_n_6745 ,csa_tree_add_51_79_groupi_n_7055);
  or csa_tree_add_51_79_groupi_g38502(csa_tree_add_51_79_groupi_n_7549 ,csa_tree_add_51_79_groupi_n_7033 ,csa_tree_add_51_79_groupi_n_7021);
  or csa_tree_add_51_79_groupi_g38503(csa_tree_add_51_79_groupi_n_7548 ,csa_tree_add_51_79_groupi_n_7002 ,csa_tree_add_51_79_groupi_n_7036);
  or csa_tree_add_51_79_groupi_g38504(csa_tree_add_51_79_groupi_n_7547 ,csa_tree_add_51_79_groupi_n_7032 ,csa_tree_add_51_79_groupi_n_7028);
  or csa_tree_add_51_79_groupi_g38505(csa_tree_add_51_79_groupi_n_7546 ,csa_tree_add_51_79_groupi_n_6135 ,csa_tree_add_51_79_groupi_n_6985);
  nor csa_tree_add_51_79_groupi_g38506(csa_tree_add_51_79_groupi_n_7545 ,csa_tree_add_51_79_groupi_n_6739 ,csa_tree_add_51_79_groupi_n_6981);
  and csa_tree_add_51_79_groupi_g38507(csa_tree_add_51_79_groupi_n_7544 ,csa_tree_add_51_79_groupi_n_7032 ,csa_tree_add_51_79_groupi_n_7028);
  or csa_tree_add_51_79_groupi_g38508(csa_tree_add_51_79_groupi_n_7543 ,csa_tree_add_51_79_groupi_n_7018 ,csa_tree_add_51_79_groupi_n_7006);
  or csa_tree_add_51_79_groupi_g38509(csa_tree_add_51_79_groupi_n_7542 ,csa_tree_add_51_79_groupi_n_7115 ,csa_tree_add_51_79_groupi_n_6943);
  or csa_tree_add_51_79_groupi_g38510(csa_tree_add_51_79_groupi_n_7541 ,csa_tree_add_51_79_groupi_n_7004 ,csa_tree_add_51_79_groupi_n_6994);
  and csa_tree_add_51_79_groupi_g38511(csa_tree_add_51_79_groupi_n_7540 ,csa_tree_add_51_79_groupi_n_7018 ,csa_tree_add_51_79_groupi_n_7006);
  and csa_tree_add_51_79_groupi_g38512(csa_tree_add_51_79_groupi_n_7539 ,csa_tree_add_51_79_groupi_n_7004 ,csa_tree_add_51_79_groupi_n_6994);
  or csa_tree_add_51_79_groupi_g38513(csa_tree_add_51_79_groupi_n_7538 ,csa_tree_add_51_79_groupi_n_6990 ,csa_tree_add_51_79_groupi_n_6975);
  or csa_tree_add_51_79_groupi_g38514(csa_tree_add_51_79_groupi_n_7537 ,csa_tree_add_51_79_groupi_n_6989 ,csa_tree_add_51_79_groupi_n_6986);
  and csa_tree_add_51_79_groupi_g38515(csa_tree_add_51_79_groupi_n_7536 ,csa_tree_add_51_79_groupi_n_7033 ,csa_tree_add_51_79_groupi_n_7021);
  and csa_tree_add_51_79_groupi_g38516(csa_tree_add_51_79_groupi_n_7535 ,csa_tree_add_51_79_groupi_n_6989 ,csa_tree_add_51_79_groupi_n_6986);
  or csa_tree_add_51_79_groupi_g38517(csa_tree_add_51_79_groupi_n_7534 ,csa_tree_add_51_79_groupi_n_6972 ,csa_tree_add_51_79_groupi_n_6967);
  and csa_tree_add_51_79_groupi_g38518(csa_tree_add_51_79_groupi_n_7533 ,csa_tree_add_51_79_groupi_n_6990 ,csa_tree_add_51_79_groupi_n_6975);
  and csa_tree_add_51_79_groupi_g38519(csa_tree_add_51_79_groupi_n_7532 ,csa_tree_add_51_79_groupi_n_6972 ,csa_tree_add_51_79_groupi_n_6967);
  or csa_tree_add_51_79_groupi_g38520(csa_tree_add_51_79_groupi_n_7531 ,csa_tree_add_51_79_groupi_n_6965 ,csa_tree_add_51_79_groupi_n_6964);
  and csa_tree_add_51_79_groupi_g38521(csa_tree_add_51_79_groupi_n_7530 ,csa_tree_add_51_79_groupi_n_6965 ,csa_tree_add_51_79_groupi_n_6964);
  or csa_tree_add_51_79_groupi_g38522(csa_tree_add_51_79_groupi_n_7529 ,csa_tree_add_51_79_groupi_n_6735 ,csa_tree_add_51_79_groupi_n_6834);
  or csa_tree_add_51_79_groupi_g38523(csa_tree_add_51_79_groupi_n_7528 ,csa_tree_add_51_79_groupi_n_6740 ,csa_tree_add_51_79_groupi_n_6980);
  or csa_tree_add_51_79_groupi_g38524(csa_tree_add_51_79_groupi_n_7527 ,csa_tree_add_51_79_groupi_n_7060 ,csa_tree_add_51_79_groupi_n_7059);
  and csa_tree_add_51_79_groupi_g38525(csa_tree_add_51_79_groupi_n_7526 ,csa_tree_add_51_79_groupi_n_7060 ,csa_tree_add_51_79_groupi_n_7059);
  or csa_tree_add_51_79_groupi_g38526(csa_tree_add_51_79_groupi_n_7525 ,csa_tree_add_51_79_groupi_n_6999 ,csa_tree_add_51_79_groupi_n_6995);
  nor csa_tree_add_51_79_groupi_g38527(csa_tree_add_51_79_groupi_n_7524 ,csa_tree_add_51_79_groupi_n_6848 ,csa_tree_add_51_79_groupi_n_6835);
  nor csa_tree_add_51_79_groupi_g38528(csa_tree_add_51_79_groupi_n_7523 ,csa_tree_add_51_79_groupi_n_6136 ,csa_tree_add_51_79_groupi_n_6984);
  or csa_tree_add_51_79_groupi_g38529(csa_tree_add_51_79_groupi_n_7522 ,csa_tree_add_51_79_groupi_n_7052 ,csa_tree_add_51_79_groupi_n_7051);
  or csa_tree_add_51_79_groupi_g38530(csa_tree_add_51_79_groupi_n_7521 ,csa_tree_add_51_79_groupi_n_6743 ,csa_tree_add_51_79_groupi_n_7040);
  and csa_tree_add_51_79_groupi_g38531(csa_tree_add_51_79_groupi_n_7520 ,csa_tree_add_51_79_groupi_n_7052 ,csa_tree_add_51_79_groupi_n_7051);
  or csa_tree_add_51_79_groupi_g38532(csa_tree_add_51_79_groupi_n_7519 ,csa_tree_add_51_79_groupi_n_7046 ,csa_tree_add_51_79_groupi_n_7041);
  or csa_tree_add_51_79_groupi_g38533(csa_tree_add_51_79_groupi_n_7518 ,csa_tree_add_51_79_groupi_n_7044 ,csa_tree_add_51_79_groupi_n_7043);
  or csa_tree_add_51_79_groupi_g38534(csa_tree_add_51_79_groupi_n_7517 ,csa_tree_add_51_79_groupi_n_7038 ,csa_tree_add_51_79_groupi_n_7023);
  and csa_tree_add_51_79_groupi_g38535(csa_tree_add_51_79_groupi_n_7516 ,csa_tree_add_51_79_groupi_n_7044 ,csa_tree_add_51_79_groupi_n_7043);
  or csa_tree_add_51_79_groupi_g38536(csa_tree_add_51_79_groupi_n_7515 ,csa_tree_add_51_79_groupi_n_7037 ,csa_tree_add_51_79_groupi_n_7034);
  nor csa_tree_add_51_79_groupi_g38537(csa_tree_add_51_79_groupi_n_7514 ,csa_tree_add_51_79_groupi_n_7045 ,csa_tree_add_51_79_groupi_n_7042);
  or csa_tree_add_51_79_groupi_g38538(csa_tree_add_51_79_groupi_n_7513 ,csa_tree_add_51_79_groupi_n_7031 ,csa_tree_add_51_79_groupi_n_7030);
  and csa_tree_add_51_79_groupi_g38539(csa_tree_add_51_79_groupi_n_7512 ,csa_tree_add_51_79_groupi_n_7037 ,csa_tree_add_51_79_groupi_n_7034);
  and csa_tree_add_51_79_groupi_g38540(csa_tree_add_51_79_groupi_n_7511 ,csa_tree_add_51_79_groupi_n_6746 ,csa_tree_add_51_79_groupi_n_6979);
  and csa_tree_add_51_79_groupi_g38541(csa_tree_add_51_79_groupi_n_7510 ,csa_tree_add_51_79_groupi_n_6743 ,csa_tree_add_51_79_groupi_n_7040);
  or csa_tree_add_51_79_groupi_g38542(csa_tree_add_51_79_groupi_n_7509 ,csa_tree_add_51_79_groupi_n_7027 ,csa_tree_add_51_79_groupi_n_7026);
  and csa_tree_add_51_79_groupi_g38543(csa_tree_add_51_79_groupi_n_7508 ,csa_tree_add_51_79_groupi_n_7031 ,csa_tree_add_51_79_groupi_n_7030);
  nor csa_tree_add_51_79_groupi_g38544(csa_tree_add_51_79_groupi_n_7507 ,csa_tree_add_51_79_groupi_n_5851 ,csa_tree_add_51_79_groupi_n_6820);
  nor csa_tree_add_51_79_groupi_g38545(csa_tree_add_51_79_groupi_n_7506 ,csa_tree_add_51_79_groupi_n_6870 ,csa_tree_add_51_79_groupi_n_7025);
  and csa_tree_add_51_79_groupi_g38546(csa_tree_add_51_79_groupi_n_7505 ,csa_tree_add_51_79_groupi_n_6128 ,csa_tree_add_51_79_groupi_n_7000);
  or csa_tree_add_51_79_groupi_g38547(csa_tree_add_51_79_groupi_n_7504 ,csa_tree_add_51_79_groupi_n_6871 ,csa_tree_add_51_79_groupi_n_7024);
  or csa_tree_add_51_79_groupi_g38548(csa_tree_add_51_79_groupi_n_7503 ,csa_tree_add_51_79_groupi_n_23 ,csa_tree_add_51_79_groupi_n_14);
  and csa_tree_add_51_79_groupi_g38549(csa_tree_add_51_79_groupi_n_7502 ,csa_tree_add_51_79_groupi_n_7027 ,csa_tree_add_51_79_groupi_n_7026);
  or csa_tree_add_51_79_groupi_g38550(csa_tree_add_51_79_groupi_n_7501 ,csa_tree_add_51_79_groupi_n_7001 ,csa_tree_add_51_79_groupi_n_6825);
  or csa_tree_add_51_79_groupi_g38551(csa_tree_add_51_79_groupi_n_7500 ,csa_tree_add_51_79_groupi_n_7016 ,csa_tree_add_51_79_groupi_n_7014);
  and csa_tree_add_51_79_groupi_g38552(csa_tree_add_51_79_groupi_n_7499 ,csa_tree_add_51_79_groupi_n_7016 ,csa_tree_add_51_79_groupi_n_7014);
  or csa_tree_add_51_79_groupi_g38553(csa_tree_add_51_79_groupi_n_7498 ,csa_tree_add_51_79_groupi_n_7039 ,csa_tree_add_51_79_groupi_n_6992);
  or csa_tree_add_51_79_groupi_g38554(csa_tree_add_51_79_groupi_n_7497 ,csa_tree_add_51_79_groupi_n_6133 ,csa_tree_add_51_79_groupi_n_7010);
  or csa_tree_add_51_79_groupi_g38555(csa_tree_add_51_79_groupi_n_7496 ,csa_tree_add_51_79_groupi_n_5308 ,csa_tree_add_51_79_groupi_n_7008);
  nor csa_tree_add_51_79_groupi_g38556(csa_tree_add_51_79_groupi_n_7495 ,csa_tree_add_51_79_groupi_n_6843 ,csa_tree_add_51_79_groupi_n_6836);
  nor csa_tree_add_51_79_groupi_g38557(csa_tree_add_51_79_groupi_n_7494 ,csa_tree_add_51_79_groupi_n_5309 ,csa_tree_add_51_79_groupi_n_7007);
  or csa_tree_add_51_79_groupi_g38558(csa_tree_add_51_79_groupi_n_7493 ,csa_tree_add_51_79_groupi_n_6868 ,csa_tree_add_51_79_groupi_n_6997);
  or csa_tree_add_51_79_groupi_g38559(csa_tree_add_51_79_groupi_n_7492 ,csa_tree_add_51_79_groupi_n_6998 ,csa_tree_add_51_79_groupi_n_6991);
  or csa_tree_add_51_79_groupi_g38560(csa_tree_add_51_79_groupi_n_7491 ,csa_tree_add_51_79_groupi_n_5865 ,csa_tree_add_51_79_groupi_n_6952);
  and csa_tree_add_51_79_groupi_g38561(csa_tree_add_51_79_groupi_n_7490 ,csa_tree_add_51_79_groupi_n_6999 ,csa_tree_add_51_79_groupi_n_6995);
  nor csa_tree_add_51_79_groupi_g38562(csa_tree_add_51_79_groupi_n_7489 ,csa_tree_add_51_79_groupi_n_6134 ,csa_tree_add_51_79_groupi_n_7009);
  nor csa_tree_add_51_79_groupi_g38563(csa_tree_add_51_79_groupi_n_7488 ,csa_tree_add_51_79_groupi_n_6869 ,csa_tree_add_51_79_groupi_n_6996);
  or csa_tree_add_51_79_groupi_g38564(csa_tree_add_51_79_groupi_n_7487 ,csa_tree_add_51_79_groupi_n_6866 ,csa_tree_add_51_79_groupi_n_6988);
  or csa_tree_add_51_79_groupi_g38565(csa_tree_add_51_79_groupi_n_7486 ,csa_tree_add_51_79_groupi_n_6453 ,csa_tree_add_51_79_groupi_n_6814);
  or csa_tree_add_51_79_groupi_g38566(csa_tree_add_51_79_groupi_n_7485 ,csa_tree_add_51_79_groupi_n_6746 ,csa_tree_add_51_79_groupi_n_6979);
  and csa_tree_add_51_79_groupi_g38567(csa_tree_add_51_79_groupi_n_7484 ,csa_tree_add_51_79_groupi_n_7038 ,csa_tree_add_51_79_groupi_n_7023);
  or csa_tree_add_51_79_groupi_g38568(csa_tree_add_51_79_groupi_n_7483 ,csa_tree_add_51_79_groupi_n_6983 ,csa_tree_add_51_79_groupi_n_6982);
  and csa_tree_add_51_79_groupi_g38569(csa_tree_add_51_79_groupi_n_7482 ,csa_tree_add_51_79_groupi_n_6983 ,csa_tree_add_51_79_groupi_n_6982);
  and csa_tree_add_51_79_groupi_g38570(csa_tree_add_51_79_groupi_n_7481 ,csa_tree_add_51_79_groupi_n_6998 ,csa_tree_add_51_79_groupi_n_6991);
  or csa_tree_add_51_79_groupi_g38571(csa_tree_add_51_79_groupi_n_7480 ,csa_tree_add_51_79_groupi_n_6978 ,csa_tree_add_51_79_groupi_n_6970);
  or csa_tree_add_51_79_groupi_g38572(csa_tree_add_51_79_groupi_n_7479 ,csa_tree_add_51_79_groupi_n_6890 ,csa_tree_add_51_79_groupi_n_6977);
  or csa_tree_add_51_79_groupi_g38573(csa_tree_add_51_79_groupi_n_7478 ,csa_tree_add_51_79_groupi_n_6976 ,csa_tree_add_51_79_groupi_n_6974);
  and csa_tree_add_51_79_groupi_g38574(csa_tree_add_51_79_groupi_n_7477 ,csa_tree_add_51_79_groupi_n_6890 ,csa_tree_add_51_79_groupi_n_6977);
  or csa_tree_add_51_79_groupi_g38575(csa_tree_add_51_79_groupi_n_7476 ,csa_tree_add_51_79_groupi_n_7070 ,csa_tree_add_51_79_groupi_n_6956);
  and csa_tree_add_51_79_groupi_g38576(csa_tree_add_51_79_groupi_n_7475 ,csa_tree_add_51_79_groupi_n_6976 ,csa_tree_add_51_79_groupi_n_6974);
  and csa_tree_add_51_79_groupi_g38577(csa_tree_add_51_79_groupi_n_7474 ,csa_tree_add_51_79_groupi_n_6978 ,csa_tree_add_51_79_groupi_n_6970);
  or csa_tree_add_51_79_groupi_g38578(csa_tree_add_51_79_groupi_n_7473 ,csa_tree_add_51_79_groupi_n_6962 ,csa_tree_add_51_79_groupi_n_6817);
  or csa_tree_add_51_79_groupi_g38579(csa_tree_add_51_79_groupi_n_7472 ,csa_tree_add_51_79_groupi_n_7054 ,csa_tree_add_51_79_groupi_n_7013);
  and csa_tree_add_51_79_groupi_g38580(csa_tree_add_51_79_groupi_n_7471 ,csa_tree_add_51_79_groupi_n_6962 ,csa_tree_add_51_79_groupi_n_6817);
  or csa_tree_add_51_79_groupi_g38581(csa_tree_add_51_79_groupi_n_7470 ,csa_tree_add_51_79_groupi_n_6865 ,csa_tree_add_51_79_groupi_n_6821);
  and csa_tree_add_51_79_groupi_g38582(csa_tree_add_51_79_groupi_n_7469 ,csa_tree_add_51_79_groupi_n_6865 ,csa_tree_add_51_79_groupi_n_6821);
  or csa_tree_add_51_79_groupi_g38583(csa_tree_add_51_79_groupi_n_7468 ,csa_tree_add_51_79_groupi_n_6904 ,csa_tree_add_51_79_groupi_n_6946);
  and csa_tree_add_51_79_groupi_g38584(csa_tree_add_51_79_groupi_n_7467 ,csa_tree_add_51_79_groupi_n_7039 ,csa_tree_add_51_79_groupi_n_6992);
  and csa_tree_add_51_79_groupi_g38585(csa_tree_add_51_79_groupi_n_7466 ,csa_tree_add_51_79_groupi_n_6879 ,csa_tree_add_51_79_groupi_n_6878);
  or csa_tree_add_51_79_groupi_g38586(csa_tree_add_51_79_groupi_n_7465 ,csa_tree_add_51_79_groupi_n_6758 ,csa_tree_add_51_79_groupi_n_6811);
  nor csa_tree_add_51_79_groupi_g38587(csa_tree_add_51_79_groupi_n_7464 ,csa_tree_add_51_79_groupi_n_6841 ,csa_tree_add_51_79_groupi_n_6837);
  or csa_tree_add_51_79_groupi_g38588(csa_tree_add_51_79_groupi_n_7463 ,csa_tree_add_51_79_groupi_n_6840 ,csa_tree_add_51_79_groupi_n_6851);
  or csa_tree_add_51_79_groupi_g38589(csa_tree_add_51_79_groupi_n_7462 ,csa_tree_add_51_79_groupi_n_6856 ,csa_tree_add_51_79_groupi_n_6858);
  and csa_tree_add_51_79_groupi_g38590(csa_tree_add_51_79_groupi_n_7461 ,csa_tree_add_51_79_groupi_n_6862 ,csa_tree_add_51_79_groupi_n_6873);
  and csa_tree_add_51_79_groupi_g38591(csa_tree_add_51_79_groupi_n_7460 ,csa_tree_add_51_79_groupi_n_7054 ,csa_tree_add_51_79_groupi_n_7013);
  nor csa_tree_add_51_79_groupi_g38592(csa_tree_add_51_79_groupi_n_7459 ,csa_tree_add_51_79_groupi_n_6722 ,csa_tree_add_51_79_groupi_n_6853);
  or csa_tree_add_51_79_groupi_g38593(csa_tree_add_51_79_groupi_n_7458 ,csa_tree_add_51_79_groupi_n_6862 ,csa_tree_add_51_79_groupi_n_6873);
  and csa_tree_add_51_79_groupi_g38594(csa_tree_add_51_79_groupi_n_7457 ,csa_tree_add_51_79_groupi_n_6856 ,csa_tree_add_51_79_groupi_n_6858);
  or csa_tree_add_51_79_groupi_g38595(csa_tree_add_51_79_groupi_n_7456 ,csa_tree_add_51_79_groupi_n_6863 ,csa_tree_add_51_79_groupi_n_6864);
  or csa_tree_add_51_79_groupi_g38596(csa_tree_add_51_79_groupi_n_7455 ,csa_tree_add_51_79_groupi_n_7029 ,csa_tree_add_51_79_groupi_n_6827);
  and csa_tree_add_51_79_groupi_g38597(csa_tree_add_51_79_groupi_n_7454 ,csa_tree_add_51_79_groupi_n_6863 ,csa_tree_add_51_79_groupi_n_6864);
  or csa_tree_add_51_79_groupi_g38598(csa_tree_add_51_79_groupi_n_7453 ,csa_tree_add_51_79_groupi_n_6457 ,csa_tree_add_51_79_groupi_n_6796);
  or csa_tree_add_51_79_groupi_g38599(csa_tree_add_51_79_groupi_n_7452 ,csa_tree_add_51_79_groupi_n_6458 ,csa_tree_add_51_79_groupi_n_6792);
  or csa_tree_add_51_79_groupi_g38600(csa_tree_add_51_79_groupi_n_7451 ,csa_tree_add_51_79_groupi_n_6912 ,csa_tree_add_51_79_groupi_n_6810);
  or csa_tree_add_51_79_groupi_g38601(csa_tree_add_51_79_groupi_n_7450 ,csa_tree_add_51_79_groupi_n_6879 ,csa_tree_add_51_79_groupi_n_6878);
  nor csa_tree_add_51_79_groupi_g38602(csa_tree_add_51_79_groupi_n_7449 ,csa_tree_add_51_79_groupi_n_6867 ,csa_tree_add_51_79_groupi_n_6987);
  and csa_tree_add_51_79_groupi_g38603(csa_tree_add_51_79_groupi_n_7448 ,csa_tree_add_51_79_groupi_n_7001 ,csa_tree_add_51_79_groupi_n_6825);
  or csa_tree_add_51_79_groupi_g38604(csa_tree_add_51_79_groupi_n_7447 ,csa_tree_add_51_79_groupi_n_6721 ,csa_tree_add_51_79_groupi_n_6852);
  or csa_tree_add_51_79_groupi_g38605(csa_tree_add_51_79_groupi_n_7446 ,csa_tree_add_51_79_groupi_n_18 ,csa_tree_add_51_79_groupi_n_17);
  or csa_tree_add_51_79_groupi_g38606(csa_tree_add_51_79_groupi_n_7445 ,csa_tree_add_51_79_groupi_n_6876 ,csa_tree_add_51_79_groupi_n_6885);
  and csa_tree_add_51_79_groupi_g38607(csa_tree_add_51_79_groupi_n_7444 ,csa_tree_add_51_79_groupi_n_6891 ,csa_tree_add_51_79_groupi_n_6882);
  or csa_tree_add_51_79_groupi_g38608(csa_tree_add_51_79_groupi_n_7443 ,csa_tree_add_51_79_groupi_n_6519 ,csa_tree_add_51_79_groupi_n_6913);
  nor csa_tree_add_51_79_groupi_g38609(csa_tree_add_51_79_groupi_n_7442 ,csa_tree_add_51_79_groupi_n_6839 ,csa_tree_add_51_79_groupi_n_6838);
  nor csa_tree_add_51_79_groupi_g38610(csa_tree_add_51_79_groupi_n_7441 ,csa_tree_add_51_79_groupi_n_6877 ,csa_tree_add_51_79_groupi_n_6884);
  and csa_tree_add_51_79_groupi_g38611(csa_tree_add_51_79_groupi_n_7440 ,csa_tree_add_51_79_groupi_n_7082 ,csa_tree_add_51_79_groupi_n_6789);
  or csa_tree_add_51_79_groupi_g38612(csa_tree_add_51_79_groupi_n_7439 ,csa_tree_add_51_79_groupi_n_6938 ,csa_tree_add_51_79_groupi_n_6784);
  or csa_tree_add_51_79_groupi_g38613(csa_tree_add_51_79_groupi_n_7438 ,csa_tree_add_51_79_groupi_n_6894 ,csa_tree_add_51_79_groupi_n_6893);
  or csa_tree_add_51_79_groupi_g38614(csa_tree_add_51_79_groupi_n_7437 ,csa_tree_add_51_79_groupi_n_6935 ,csa_tree_add_51_79_groupi_n_6787);
  and csa_tree_add_51_79_groupi_g38615(csa_tree_add_51_79_groupi_n_7436 ,csa_tree_add_51_79_groupi_n_6894 ,csa_tree_add_51_79_groupi_n_6893);
  and csa_tree_add_51_79_groupi_g38616(csa_tree_add_51_79_groupi_n_7435 ,csa_tree_add_51_79_groupi_n_7029 ,csa_tree_add_51_79_groupi_n_6827);
  or csa_tree_add_51_79_groupi_g38617(csa_tree_add_51_79_groupi_n_7434 ,csa_tree_add_51_79_groupi_n_6872 ,csa_tree_add_51_79_groupi_n_6898);
  or csa_tree_add_51_79_groupi_g38618(csa_tree_add_51_79_groupi_n_7433 ,csa_tree_add_51_79_groupi_n_6824 ,csa_tree_add_51_79_groupi_n_6895);
  nor csa_tree_add_51_79_groupi_g38619(csa_tree_add_51_79_groupi_n_7432 ,csa_tree_add_51_79_groupi_n_5852 ,csa_tree_add_51_79_groupi_n_6888);
  and csa_tree_add_51_79_groupi_g38620(csa_tree_add_51_79_groupi_n_7431 ,csa_tree_add_51_79_groupi_n_6824 ,csa_tree_add_51_79_groupi_n_6895);
  or csa_tree_add_51_79_groupi_g38621(csa_tree_add_51_79_groupi_n_7430 ,csa_tree_add_51_79_groupi_n_6892 ,csa_tree_add_51_79_groupi_n_6889);
  and csa_tree_add_51_79_groupi_g38622(csa_tree_add_51_79_groupi_n_7429 ,csa_tree_add_51_79_groupi_n_6872 ,csa_tree_add_51_79_groupi_n_6898);
  and csa_tree_add_51_79_groupi_g38623(csa_tree_add_51_79_groupi_n_7428 ,csa_tree_add_51_79_groupi_n_5851 ,csa_tree_add_51_79_groupi_n_6820);
  and csa_tree_add_51_79_groupi_g38624(csa_tree_add_51_79_groupi_n_7427 ,csa_tree_add_51_79_groupi_n_6892 ,csa_tree_add_51_79_groupi_n_6889);
  or csa_tree_add_51_79_groupi_g38625(csa_tree_add_51_79_groupi_n_7426 ,csa_tree_add_51_79_groupi_n_15 ,csa_tree_add_51_79_groupi_n_16);
  or csa_tree_add_51_79_groupi_g38626(csa_tree_add_51_79_groupi_n_7425 ,csa_tree_add_51_79_groupi_n_12 ,csa_tree_add_51_79_groupi_n_19);
  or csa_tree_add_51_79_groupi_g38627(csa_tree_add_51_79_groupi_n_7424 ,csa_tree_add_51_79_groupi_n_6875 ,csa_tree_add_51_79_groupi_n_6874);
  or csa_tree_add_51_79_groupi_g38628(csa_tree_add_51_79_groupi_n_7423 ,csa_tree_add_51_79_groupi_n_5840 ,csa_tree_add_51_79_groupi_n_6860);
  and csa_tree_add_51_79_groupi_g38629(csa_tree_add_51_79_groupi_n_7422 ,csa_tree_add_51_79_groupi_n_6875 ,csa_tree_add_51_79_groupi_n_6874);
  or csa_tree_add_51_79_groupi_g38630(csa_tree_add_51_79_groupi_n_7421 ,csa_tree_add_51_79_groupi_n_6859 ,csa_tree_add_51_79_groupi_n_6828);
  or csa_tree_add_51_79_groupi_g38631(csa_tree_add_51_79_groupi_n_7420 ,csa_tree_add_51_79_groupi_n_5853 ,csa_tree_add_51_79_groupi_n_6887);
  or csa_tree_add_51_79_groupi_g38632(csa_tree_add_51_79_groupi_n_7419 ,csa_tree_add_51_79_groupi_n_6822 ,csa_tree_add_51_79_groupi_n_6896);
  and csa_tree_add_51_79_groupi_g38633(csa_tree_add_51_79_groupi_n_7418 ,csa_tree_add_51_79_groupi_n_6859 ,csa_tree_add_51_79_groupi_n_6828);
  nor csa_tree_add_51_79_groupi_g38634(csa_tree_add_51_79_groupi_n_7417 ,csa_tree_add_51_79_groupi_n_5841 ,csa_tree_add_51_79_groupi_n_6861);
  or csa_tree_add_51_79_groupi_g38635(csa_tree_add_51_79_groupi_n_7416 ,csa_tree_add_51_79_groupi_n_6819 ,csa_tree_add_51_79_groupi_n_6816);
  and csa_tree_add_51_79_groupi_g38636(csa_tree_add_51_79_groupi_n_7415 ,csa_tree_add_51_79_groupi_n_6819 ,csa_tree_add_51_79_groupi_n_6816);
  or csa_tree_add_51_79_groupi_g38637(csa_tree_add_51_79_groupi_n_7414 ,csa_tree_add_51_79_groupi_n_6891 ,csa_tree_add_51_79_groupi_n_6882);
  or csa_tree_add_51_79_groupi_g38638(csa_tree_add_51_79_groupi_n_7413 ,csa_tree_add_51_79_groupi_n_6759 ,csa_tree_add_51_79_groupi_n_6807);
  or csa_tree_add_51_79_groupi_g38639(csa_tree_add_51_79_groupi_n_7412 ,csa_tree_add_51_79_groupi_n_6969 ,csa_tree_add_51_79_groupi_n_6968);
  and csa_tree_add_51_79_groupi_g38640(csa_tree_add_51_79_groupi_n_7411 ,csa_tree_add_51_79_groupi_n_6969 ,csa_tree_add_51_79_groupi_n_6968);
  or csa_tree_add_51_79_groupi_g38641(csa_tree_add_51_79_groupi_n_7410 ,csa_tree_add_51_79_groupi_n_6880 ,csa_tree_add_51_79_groupi_n_6826);
  or csa_tree_add_51_79_groupi_g38642(csa_tree_add_51_79_groupi_n_7409 ,csa_tree_add_51_79_groupi_n_6842 ,csa_tree_add_51_79_groupi_n_6886);
  and csa_tree_add_51_79_groupi_g38643(csa_tree_add_51_79_groupi_n_7408 ,csa_tree_add_51_79_groupi_n_6842 ,csa_tree_add_51_79_groupi_n_6886);
  and csa_tree_add_51_79_groupi_g38644(csa_tree_add_51_79_groupi_n_7407 ,csa_tree_add_51_79_groupi_n_6880 ,csa_tree_add_51_79_groupi_n_6826);
  or csa_tree_add_51_79_groupi_g38645(csa_tree_add_51_79_groupi_n_7406 ,csa_tree_add_51_79_groupi_n_6881 ,csa_tree_add_51_79_groupi_n_6883);
  and csa_tree_add_51_79_groupi_g38646(csa_tree_add_51_79_groupi_n_7405 ,csa_tree_add_51_79_groupi_n_6881 ,csa_tree_add_51_79_groupi_n_6883);
  or csa_tree_add_51_79_groupi_g38647(csa_tree_add_51_79_groupi_n_7404 ,csa_tree_add_51_79_groupi_n_6459 ,csa_tree_add_51_79_groupi_n_6793);
  or csa_tree_add_51_79_groupi_g38648(csa_tree_add_51_79_groupi_n_7403 ,csa_tree_add_51_79_groupi_n_6454 ,csa_tree_add_51_79_groupi_n_6800);
  or csa_tree_add_51_79_groupi_g38649(csa_tree_add_51_79_groupi_n_7402 ,csa_tree_add_51_79_groupi_n_6456 ,csa_tree_add_51_79_groupi_n_6797);
  or csa_tree_add_51_79_groupi_g38650(csa_tree_add_51_79_groupi_n_7401 ,csa_tree_add_51_79_groupi_n_6460 ,csa_tree_add_51_79_groupi_n_6798);
  or csa_tree_add_51_79_groupi_g38651(csa_tree_add_51_79_groupi_n_7400 ,csa_tree_add_51_79_groupi_n_6761 ,csa_tree_add_51_79_groupi_n_6803);
  or csa_tree_add_51_79_groupi_g38652(csa_tree_add_51_79_groupi_n_7399 ,csa_tree_add_51_79_groupi_n_6832 ,csa_tree_add_51_79_groupi_n_6831);
  and csa_tree_add_51_79_groupi_g38653(csa_tree_add_51_79_groupi_n_7398 ,csa_tree_add_51_79_groupi_n_6832 ,csa_tree_add_51_79_groupi_n_6831);
  or csa_tree_add_51_79_groupi_g38654(csa_tree_add_51_79_groupi_n_7397 ,csa_tree_add_51_79_groupi_n_6830 ,csa_tree_add_51_79_groupi_n_6829);
  and csa_tree_add_51_79_groupi_g38655(csa_tree_add_51_79_groupi_n_7396 ,csa_tree_add_51_79_groupi_n_6830 ,csa_tree_add_51_79_groupi_n_6829);
  nor csa_tree_add_51_79_groupi_g38656(csa_tree_add_51_79_groupi_n_7395 ,csa_tree_add_51_79_groupi_n_6736 ,csa_tree_add_51_79_groupi_n_6833);
  nor csa_tree_add_51_79_groupi_g38657(csa_tree_add_51_79_groupi_n_7394 ,csa_tree_add_51_79_groupi_n_6150 ,csa_tree_add_51_79_groupi_n_6941);
  or csa_tree_add_51_79_groupi_g38658(csa_tree_add_51_79_groupi_n_7393 ,csa_tree_add_51_79_groupi_n_6762 ,csa_tree_add_51_79_groupi_n_6805);
  or csa_tree_add_51_79_groupi_g38659(csa_tree_add_51_79_groupi_n_7392 ,csa_tree_add_51_79_groupi_n_22 ,csa_tree_add_51_79_groupi_n_21);
  nor csa_tree_add_51_79_groupi_g38660(csa_tree_add_51_79_groupi_n_7391 ,csa_tree_add_51_79_groupi_n_6847 ,csa_tree_add_51_79_groupi_n_6846);
  or csa_tree_add_51_79_groupi_g38661(csa_tree_add_51_79_groupi_n_7390 ,csa_tree_add_51_79_groupi_n_20 ,csa_tree_add_51_79_groupi_n_13);
  nor csa_tree_add_51_79_groupi_g38662(csa_tree_add_51_79_groupi_n_7389 ,csa_tree_add_51_79_groupi_n_6845 ,csa_tree_add_51_79_groupi_n_6844);
  xnor csa_tree_add_51_79_groupi_g38663(csa_tree_add_51_79_groupi_n_7635 ,csa_tree_add_51_79_groupi_n_5541 ,csa_tree_add_51_79_groupi_n_6366);
  and csa_tree_add_51_79_groupi_g38664(csa_tree_add_51_79_groupi_n_7634 ,csa_tree_add_51_79_groupi_n_6599 ,csa_tree_add_51_79_groupi_n_6947);
  or csa_tree_add_51_79_groupi_g38665(csa_tree_add_51_79_groupi_n_7633 ,csa_tree_add_51_79_groupi_n_6634 ,csa_tree_add_51_79_groupi_n_6959);
  xnor csa_tree_add_51_79_groupi_g38666(csa_tree_add_51_79_groupi_n_7631 ,csa_tree_add_51_79_groupi_n_4904 ,csa_tree_add_51_79_groupi_n_6251);
  xnor csa_tree_add_51_79_groupi_g38667(csa_tree_add_51_79_groupi_n_7630 ,csa_tree_add_51_79_groupi_n_4864 ,csa_tree_add_51_79_groupi_n_6219);
  xnor csa_tree_add_51_79_groupi_g38668(csa_tree_add_51_79_groupi_n_7629 ,csa_tree_add_51_79_groupi_n_4874 ,csa_tree_add_51_79_groupi_n_6214);
  xnor csa_tree_add_51_79_groupi_g38669(csa_tree_add_51_79_groupi_n_7628 ,csa_tree_add_51_79_groupi_n_5520 ,csa_tree_add_51_79_groupi_n_6388);
  xor csa_tree_add_51_79_groupi_g38670(csa_tree_add_51_79_groupi_n_7627 ,csa_tree_add_51_79_groupi_n_3817 ,csa_tree_add_51_79_groupi_n_6224);
  xnor csa_tree_add_51_79_groupi_g38671(csa_tree_add_51_79_groupi_n_7626 ,csa_tree_add_51_79_groupi_n_3227 ,csa_tree_add_51_79_groupi_n_6201);
  xor csa_tree_add_51_79_groupi_g38672(csa_tree_add_51_79_groupi_n_7625 ,csa_tree_add_51_79_groupi_n_4858 ,csa_tree_add_51_79_groupi_n_6194);
  xnor csa_tree_add_51_79_groupi_g38673(csa_tree_add_51_79_groupi_n_7624 ,csa_tree_add_51_79_groupi_n_5112 ,csa_tree_add_51_79_groupi_n_6377);
  xor csa_tree_add_51_79_groupi_g38674(csa_tree_add_51_79_groupi_n_7623 ,csa_tree_add_51_79_groupi_n_3229 ,csa_tree_add_51_79_groupi_n_6188);
  xnor csa_tree_add_51_79_groupi_g38675(csa_tree_add_51_79_groupi_n_7621 ,csa_tree_add_51_79_groupi_n_3812 ,csa_tree_add_51_79_groupi_n_6179);
  xnor csa_tree_add_51_79_groupi_g38676(csa_tree_add_51_79_groupi_n_7619 ,csa_tree_add_51_79_groupi_n_3233 ,csa_tree_add_51_79_groupi_n_6237);
  xnor csa_tree_add_51_79_groupi_g38677(csa_tree_add_51_79_groupi_n_7618 ,csa_tree_add_51_79_groupi_n_3792 ,csa_tree_add_51_79_groupi_n_6235);
  and csa_tree_add_51_79_groupi_g38678(csa_tree_add_51_79_groupi_n_7617 ,csa_tree_add_51_79_groupi_n_6586 ,csa_tree_add_51_79_groupi_n_6950);
  xnor csa_tree_add_51_79_groupi_g38679(csa_tree_add_51_79_groupi_n_7616 ,csa_tree_add_51_79_groupi_n_4849 ,csa_tree_add_51_79_groupi_n_6383);
  xnor csa_tree_add_51_79_groupi_g38680(csa_tree_add_51_79_groupi_n_7614 ,csa_tree_add_51_79_groupi_n_5104 ,csa_tree_add_51_79_groupi_n_6370);
  and csa_tree_add_51_79_groupi_g38681(csa_tree_add_51_79_groupi_n_7611 ,csa_tree_add_51_79_groupi_n_6538 ,csa_tree_add_51_79_groupi_n_6783);
  and csa_tree_add_51_79_groupi_g38682(csa_tree_add_51_79_groupi_n_7610 ,csa_tree_add_51_79_groupi_n_6540 ,csa_tree_add_51_79_groupi_n_6813);
  or csa_tree_add_51_79_groupi_g38683(csa_tree_add_51_79_groupi_n_7609 ,csa_tree_add_51_79_groupi_n_6509 ,csa_tree_add_51_79_groupi_n_6790);
  or csa_tree_add_51_79_groupi_g38684(csa_tree_add_51_79_groupi_n_7607 ,csa_tree_add_51_79_groupi_n_6592 ,csa_tree_add_51_79_groupi_n_6954);
  xnor csa_tree_add_51_79_groupi_g38685(csa_tree_add_51_79_groupi_n_7605 ,csa_tree_add_51_79_groupi_n_5452 ,csa_tree_add_51_79_groupi_n_6382);
  xnor csa_tree_add_51_79_groupi_g38686(csa_tree_add_51_79_groupi_n_7603 ,csa_tree_add_51_79_groupi_n_4843 ,csa_tree_add_51_79_groupi_n_6386);
  xnor csa_tree_add_51_79_groupi_g38687(csa_tree_add_51_79_groupi_n_7601 ,csa_tree_add_51_79_groupi_n_3197 ,csa_tree_add_51_79_groupi_n_6195);
  xnor csa_tree_add_51_79_groupi_g38688(csa_tree_add_51_79_groupi_n_7600 ,csa_tree_add_51_79_groupi_n_5093 ,csa_tree_add_51_79_groupi_n_6379);
  xnor csa_tree_add_51_79_groupi_g38689(csa_tree_add_51_79_groupi_n_7599 ,csa_tree_add_51_79_groupi_n_5459 ,csa_tree_add_51_79_groupi_n_6378);
  and csa_tree_add_51_79_groupi_g38690(csa_tree_add_51_79_groupi_n_7598 ,csa_tree_add_51_79_groupi_n_5654 ,csa_tree_add_51_79_groupi_n_6788);
  and csa_tree_add_51_79_groupi_g38691(csa_tree_add_51_79_groupi_n_7596 ,csa_tree_add_51_79_groupi_n_6482 ,csa_tree_add_51_79_groupi_n_6786);
  xnor csa_tree_add_51_79_groupi_g38692(csa_tree_add_51_79_groupi_n_7595 ,csa_tree_add_51_79_groupi_n_3813 ,csa_tree_add_51_79_groupi_n_6191);
  xnor csa_tree_add_51_79_groupi_g38693(csa_tree_add_51_79_groupi_n_7593 ,csa_tree_add_51_79_groupi_n_5435 ,csa_tree_add_51_79_groupi_n_6350);
  and csa_tree_add_51_79_groupi_g38694(csa_tree_add_51_79_groupi_n_7592 ,csa_tree_add_51_79_groupi_n_5749 ,csa_tree_add_51_79_groupi_n_6778);
  xnor csa_tree_add_51_79_groupi_g38696(csa_tree_add_51_79_groupi_n_7589 ,csa_tree_add_51_79_groupi_n_3762 ,csa_tree_add_51_79_groupi_n_6180);
  xnor csa_tree_add_51_79_groupi_g38697(csa_tree_add_51_79_groupi_n_7587 ,csa_tree_add_51_79_groupi_n_5503 ,csa_tree_add_51_79_groupi_n_6337);
  xnor csa_tree_add_51_79_groupi_g38698(csa_tree_add_51_79_groupi_n_7585 ,csa_tree_add_51_79_groupi_n_5268 ,csa_tree_add_51_79_groupi_n_6389);
  and csa_tree_add_51_79_groupi_g38699(csa_tree_add_51_79_groupi_n_7583 ,csa_tree_add_51_79_groupi_n_6508 ,csa_tree_add_51_79_groupi_n_6785);
  xnor csa_tree_add_51_79_groupi_g38700(csa_tree_add_51_79_groupi_n_7582 ,csa_tree_add_51_79_groupi_n_5375 ,csa_tree_add_51_79_groupi_n_6367);
  xnor csa_tree_add_51_79_groupi_g38701(csa_tree_add_51_79_groupi_n_7580 ,csa_tree_add_51_79_groupi_n_4962 ,csa_tree_add_51_79_groupi_n_6384);
  xnor csa_tree_add_51_79_groupi_g38702(csa_tree_add_51_79_groupi_n_7578 ,csa_tree_add_51_79_groupi_n_5250 ,csa_tree_add_51_79_groupi_n_6244);
  and csa_tree_add_51_79_groupi_g38703(csa_tree_add_51_79_groupi_n_7576 ,csa_tree_add_51_79_groupi_n_6649 ,csa_tree_add_51_79_groupi_n_6944);
  not csa_tree_add_51_79_groupi_g38704(csa_tree_add_51_79_groupi_n_7351 ,csa_tree_add_51_79_groupi_n_7350);
  not csa_tree_add_51_79_groupi_g38705(csa_tree_add_51_79_groupi_n_7346 ,csa_tree_add_51_79_groupi_n_7345);
  not csa_tree_add_51_79_groupi_g38706(csa_tree_add_51_79_groupi_n_7315 ,csa_tree_add_51_79_groupi_n_7316);
  not csa_tree_add_51_79_groupi_g38707(csa_tree_add_51_79_groupi_n_7312 ,csa_tree_add_51_79_groupi_n_7313);
  not csa_tree_add_51_79_groupi_g38709(csa_tree_add_51_79_groupi_n_7306 ,csa_tree_add_51_79_groupi_n_7307);
  not csa_tree_add_51_79_groupi_g38710(csa_tree_add_51_79_groupi_n_7303 ,csa_tree_add_51_79_groupi_n_7304);
  not csa_tree_add_51_79_groupi_g38711(csa_tree_add_51_79_groupi_n_7301 ,csa_tree_add_51_79_groupi_n_7300);
  not csa_tree_add_51_79_groupi_g38712(csa_tree_add_51_79_groupi_n_7292 ,csa_tree_add_51_79_groupi_n_7293);
  not csa_tree_add_51_79_groupi_g38713(csa_tree_add_51_79_groupi_n_7291 ,csa_tree_add_51_79_groupi_n_7290);
  not csa_tree_add_51_79_groupi_g38714(csa_tree_add_51_79_groupi_n_7288 ,csa_tree_add_51_79_groupi_n_7289);
  not csa_tree_add_51_79_groupi_g38715(csa_tree_add_51_79_groupi_n_7286 ,csa_tree_add_51_79_groupi_n_7287);
  not csa_tree_add_51_79_groupi_g38716(csa_tree_add_51_79_groupi_n_7274 ,csa_tree_add_51_79_groupi_n_7275);
  not csa_tree_add_51_79_groupi_g38717(csa_tree_add_51_79_groupi_n_7267 ,csa_tree_add_51_79_groupi_n_7268);
  not csa_tree_add_51_79_groupi_g38718(csa_tree_add_51_79_groupi_n_7261 ,csa_tree_add_51_79_groupi_n_7262);
  not csa_tree_add_51_79_groupi_g38719(csa_tree_add_51_79_groupi_n_7255 ,csa_tree_add_51_79_groupi_n_7256);
  not csa_tree_add_51_79_groupi_g38720(csa_tree_add_51_79_groupi_n_7250 ,csa_tree_add_51_79_groupi_n_7251);
  not csa_tree_add_51_79_groupi_g38721(csa_tree_add_51_79_groupi_n_7246 ,csa_tree_add_51_79_groupi_n_7247);
  not csa_tree_add_51_79_groupi_g38722(csa_tree_add_51_79_groupi_n_7243 ,csa_tree_add_51_79_groupi_n_7244);
  not csa_tree_add_51_79_groupi_g38723(csa_tree_add_51_79_groupi_n_7239 ,csa_tree_add_51_79_groupi_n_7240);
  not csa_tree_add_51_79_groupi_g38724(csa_tree_add_51_79_groupi_n_7234 ,csa_tree_add_51_79_groupi_n_7235);
  not csa_tree_add_51_79_groupi_g38725(csa_tree_add_51_79_groupi_n_7231 ,csa_tree_add_51_79_groupi_n_7232);
  not csa_tree_add_51_79_groupi_g38726(csa_tree_add_51_79_groupi_n_7218 ,csa_tree_add_51_79_groupi_n_7219);
  not csa_tree_add_51_79_groupi_g38727(csa_tree_add_51_79_groupi_n_7216 ,csa_tree_add_51_79_groupi_n_7217);
  not csa_tree_add_51_79_groupi_g38728(csa_tree_add_51_79_groupi_n_7214 ,csa_tree_add_51_79_groupi_n_7215);
  not csa_tree_add_51_79_groupi_g38730(csa_tree_add_51_79_groupi_n_7208 ,csa_tree_add_51_79_groupi_n_7209);
  not csa_tree_add_51_79_groupi_g38731(csa_tree_add_51_79_groupi_n_7206 ,csa_tree_add_51_79_groupi_n_0);
  not csa_tree_add_51_79_groupi_g38732(csa_tree_add_51_79_groupi_n_7197 ,csa_tree_add_51_79_groupi_n_7198);
  not csa_tree_add_51_79_groupi_g38733(csa_tree_add_51_79_groupi_n_7195 ,csa_tree_add_51_79_groupi_n_7196);
  not csa_tree_add_51_79_groupi_g38734(csa_tree_add_51_79_groupi_n_7193 ,csa_tree_add_51_79_groupi_n_7194);
  not csa_tree_add_51_79_groupi_g38735(csa_tree_add_51_79_groupi_n_7188 ,csa_tree_add_51_79_groupi_n_7189);
  not csa_tree_add_51_79_groupi_g38736(csa_tree_add_51_79_groupi_n_7186 ,csa_tree_add_51_79_groupi_n_7187);
  not csa_tree_add_51_79_groupi_g38737(csa_tree_add_51_79_groupi_n_7184 ,csa_tree_add_51_79_groupi_n_7185);
  not csa_tree_add_51_79_groupi_g38738(csa_tree_add_51_79_groupi_n_7180 ,csa_tree_add_51_79_groupi_n_7181);
  not csa_tree_add_51_79_groupi_g38739(csa_tree_add_51_79_groupi_n_7178 ,csa_tree_add_51_79_groupi_n_7179);
  not csa_tree_add_51_79_groupi_g38740(csa_tree_add_51_79_groupi_n_7174 ,csa_tree_add_51_79_groupi_n_7175);
  not csa_tree_add_51_79_groupi_g38741(csa_tree_add_51_79_groupi_n_7169 ,csa_tree_add_51_79_groupi_n_7170);
  not csa_tree_add_51_79_groupi_g38742(csa_tree_add_51_79_groupi_n_7163 ,csa_tree_add_51_79_groupi_n_7164);
  not csa_tree_add_51_79_groupi_g38743(csa_tree_add_51_79_groupi_n_7160 ,csa_tree_add_51_79_groupi_n_7161);
  not csa_tree_add_51_79_groupi_g38744(csa_tree_add_51_79_groupi_n_7158 ,csa_tree_add_51_79_groupi_n_7159);
  not csa_tree_add_51_79_groupi_g38745(csa_tree_add_51_79_groupi_n_7156 ,csa_tree_add_51_79_groupi_n_7157);
  not csa_tree_add_51_79_groupi_g38746(csa_tree_add_51_79_groupi_n_7154 ,csa_tree_add_51_79_groupi_n_7155);
  not csa_tree_add_51_79_groupi_g38747(csa_tree_add_51_79_groupi_n_7146 ,csa_tree_add_51_79_groupi_n_7147);
  not csa_tree_add_51_79_groupi_g38748(csa_tree_add_51_79_groupi_n_7144 ,csa_tree_add_51_79_groupi_n_7145);
  not csa_tree_add_51_79_groupi_g38749(csa_tree_add_51_79_groupi_n_7138 ,csa_tree_add_51_79_groupi_n_7139);
  not csa_tree_add_51_79_groupi_g38750(csa_tree_add_51_79_groupi_n_7136 ,csa_tree_add_51_79_groupi_n_7137);
  xnor csa_tree_add_51_79_groupi_g38751(csa_tree_add_51_79_groupi_n_7135 ,csa_tree_add_51_79_groupi_n_6439 ,csa_tree_add_51_79_groupi_n_6438);
  xnor csa_tree_add_51_79_groupi_g38752(csa_tree_add_51_79_groupi_n_7134 ,csa_tree_add_51_79_groupi_n_6762 ,csa_tree_add_51_79_groupi_n_6730);
  xnor csa_tree_add_51_79_groupi_g38753(csa_tree_add_51_79_groupi_n_7133 ,csa_tree_add_51_79_groupi_n_6440 ,csa_tree_add_51_79_groupi_n_6727);
  xnor csa_tree_add_51_79_groupi_g38754(csa_tree_add_51_79_groupi_n_7132 ,csa_tree_add_51_79_groupi_n_6460 ,csa_tree_add_51_79_groupi_n_6400);
  xnor csa_tree_add_51_79_groupi_g38755(csa_tree_add_51_79_groupi_n_7131 ,csa_tree_add_51_79_groupi_n_6759 ,csa_tree_add_51_79_groupi_n_6726);
  xnor csa_tree_add_51_79_groupi_g38756(csa_tree_add_51_79_groupi_n_7130 ,csa_tree_add_51_79_groupi_n_6758 ,csa_tree_add_51_79_groupi_n_6395);
  xnor csa_tree_add_51_79_groupi_g38757(csa_tree_add_51_79_groupi_n_7129 ,csa_tree_add_51_79_groupi_n_6448 ,csa_tree_add_51_79_groupi_n_6733);
  xnor csa_tree_add_51_79_groupi_g38758(csa_tree_add_51_79_groupi_n_7128 ,csa_tree_add_51_79_groupi_n_6737 ,csa_tree_add_51_79_groupi_n_6738);
  xnor csa_tree_add_51_79_groupi_g38759(csa_tree_add_51_79_groupi_n_7127 ,csa_tree_add_51_79_groupi_n_6435 ,csa_tree_add_51_79_groupi_n_6734);
  xnor csa_tree_add_51_79_groupi_g38760(csa_tree_add_51_79_groupi_n_7126 ,csa_tree_add_51_79_groupi_n_6748 ,csa_tree_add_51_79_groupi_n_6750);
  xnor csa_tree_add_51_79_groupi_g38761(csa_tree_add_51_79_groupi_n_7125 ,csa_tree_add_51_79_groupi_n_6444 ,csa_tree_add_51_79_groupi_n_6443);
  xnor csa_tree_add_51_79_groupi_g38762(csa_tree_add_51_79_groupi_n_7124 ,csa_tree_add_51_79_groupi_n_6447 ,csa_tree_add_51_79_groupi_n_6446);
  xnor csa_tree_add_51_79_groupi_g38763(csa_tree_add_51_79_groupi_n_7123 ,csa_tree_add_51_79_groupi_n_6457 ,csa_tree_add_51_79_groupi_n_6449);
  xnor csa_tree_add_51_79_groupi_g38764(csa_tree_add_51_79_groupi_n_7122 ,csa_tree_add_51_79_groupi_n_6450 ,csa_tree_add_51_79_groupi_n_4821);
  xnor csa_tree_add_51_79_groupi_g38765(csa_tree_add_51_79_groupi_n_7121 ,csa_tree_add_51_79_groupi_n_6416 ,csa_tree_add_51_79_groupi_n_6410);
  xnor csa_tree_add_51_79_groupi_g38766(csa_tree_add_51_79_groupi_n_7120 ,csa_tree_add_51_79_groupi_n_6434 ,csa_tree_add_51_79_groupi_n_6433);
  xnor csa_tree_add_51_79_groupi_g38767(csa_tree_add_51_79_groupi_n_7119 ,csa_tree_add_51_79_groupi_n_6127 ,csa_tree_add_51_79_groupi_n_6413);
  xnor csa_tree_add_51_79_groupi_g38768(csa_tree_add_51_79_groupi_n_7118 ,csa_tree_add_51_79_groupi_n_6455 ,csa_tree_add_51_79_groupi_n_6);
  xor csa_tree_add_51_79_groupi_g38769(csa_tree_add_51_79_groupi_n_7388 ,csa_tree_add_51_79_groupi_n_3808 ,csa_tree_add_51_79_groupi_n_6359);
  xnor csa_tree_add_51_79_groupi_g38770(csa_tree_add_51_79_groupi_n_7387 ,csa_tree_add_51_79_groupi_n_3780 ,csa_tree_add_51_79_groupi_n_6392);
  xnor csa_tree_add_51_79_groupi_g38771(csa_tree_add_51_79_groupi_n_7386 ,csa_tree_add_51_79_groupi_n_5049 ,csa_tree_add_51_79_groupi_n_6318);
  xnor csa_tree_add_51_79_groupi_g38772(csa_tree_add_51_79_groupi_n_7385 ,csa_tree_add_51_79_groupi_n_4920 ,csa_tree_add_51_79_groupi_n_6285);
  xnor csa_tree_add_51_79_groupi_g38773(csa_tree_add_51_79_groupi_n_7384 ,csa_tree_add_51_79_groupi_n_4854 ,csa_tree_add_51_79_groupi_n_6315);
  xnor csa_tree_add_51_79_groupi_g38774(csa_tree_add_51_79_groupi_n_7383 ,csa_tree_add_51_79_groupi_n_5450 ,csa_tree_add_51_79_groupi_n_6311);
  xnor csa_tree_add_51_79_groupi_g38775(csa_tree_add_51_79_groupi_n_7382 ,csa_tree_add_51_79_groupi_n_5475 ,csa_tree_add_51_79_groupi_n_6309);
  xnor csa_tree_add_51_79_groupi_g38776(csa_tree_add_51_79_groupi_n_7381 ,csa_tree_add_51_79_groupi_n_5542 ,csa_tree_add_51_79_groupi_n_6301);
  xnor csa_tree_add_51_79_groupi_g38777(csa_tree_add_51_79_groupi_n_7380 ,csa_tree_add_51_79_groupi_n_5533 ,csa_tree_add_51_79_groupi_n_6300);
  xnor csa_tree_add_51_79_groupi_g38778(csa_tree_add_51_79_groupi_n_7379 ,csa_tree_add_51_79_groupi_n_5526 ,csa_tree_add_51_79_groupi_n_6310);
  xnor csa_tree_add_51_79_groupi_g38779(csa_tree_add_51_79_groupi_n_7378 ,csa_tree_add_51_79_groupi_n_5536 ,csa_tree_add_51_79_groupi_n_6297);
  xnor csa_tree_add_51_79_groupi_g38780(csa_tree_add_51_79_groupi_n_7377 ,csa_tree_add_51_79_groupi_n_5491 ,csa_tree_add_51_79_groupi_n_6295);
  xnor csa_tree_add_51_79_groupi_g38781(csa_tree_add_51_79_groupi_n_7376 ,csa_tree_add_51_79_groupi_n_5065 ,csa_tree_add_51_79_groupi_n_6290);
  xnor csa_tree_add_51_79_groupi_g38782(csa_tree_add_51_79_groupi_n_7375 ,csa_tree_add_51_79_groupi_n_5457 ,csa_tree_add_51_79_groupi_n_6287);
  xnor csa_tree_add_51_79_groupi_g38783(csa_tree_add_51_79_groupi_n_7374 ,csa_tree_add_51_79_groupi_n_5469 ,csa_tree_add_51_79_groupi_n_6279);
  xnor csa_tree_add_51_79_groupi_g38784(csa_tree_add_51_79_groupi_n_7373 ,csa_tree_add_51_79_groupi_n_5500 ,csa_tree_add_51_79_groupi_n_6286);
  xnor csa_tree_add_51_79_groupi_g38785(csa_tree_add_51_79_groupi_n_7372 ,csa_tree_add_51_79_groupi_n_5078 ,csa_tree_add_51_79_groupi_n_6282);
  xnor csa_tree_add_51_79_groupi_g38786(csa_tree_add_51_79_groupi_n_7371 ,csa_tree_add_51_79_groupi_n_5460 ,csa_tree_add_51_79_groupi_n_6273);
  xnor csa_tree_add_51_79_groupi_g38787(csa_tree_add_51_79_groupi_n_7370 ,csa_tree_add_51_79_groupi_n_5458 ,csa_tree_add_51_79_groupi_n_6271);
  xnor csa_tree_add_51_79_groupi_g38788(csa_tree_add_51_79_groupi_n_7369 ,csa_tree_add_51_79_groupi_n_5438 ,csa_tree_add_51_79_groupi_n_6269);
  xnor csa_tree_add_51_79_groupi_g38789(csa_tree_add_51_79_groupi_n_7368 ,csa_tree_add_51_79_groupi_n_5092 ,csa_tree_add_51_79_groupi_n_6292);
  xnor csa_tree_add_51_79_groupi_g38790(csa_tree_add_51_79_groupi_n_7367 ,csa_tree_add_51_79_groupi_n_5021 ,csa_tree_add_51_79_groupi_n_6321);
  xnor csa_tree_add_51_79_groupi_g38791(csa_tree_add_51_79_groupi_n_7366 ,csa_tree_add_51_79_groupi_n_5073 ,csa_tree_add_51_79_groupi_n_6296);
  xnor csa_tree_add_51_79_groupi_g38792(csa_tree_add_51_79_groupi_n_7365 ,csa_tree_add_51_79_groupi_n_5067 ,csa_tree_add_51_79_groupi_n_6261);
  xnor csa_tree_add_51_79_groupi_g38793(csa_tree_add_51_79_groupi_n_7364 ,csa_tree_add_51_79_groupi_n_5068 ,csa_tree_add_51_79_groupi_n_6259);
  xnor csa_tree_add_51_79_groupi_g38794(csa_tree_add_51_79_groupi_n_7363 ,csa_tree_add_51_79_groupi_n_5047 ,csa_tree_add_51_79_groupi_n_6307);
  xnor csa_tree_add_51_79_groupi_g38795(csa_tree_add_51_79_groupi_n_7362 ,csa_tree_add_51_79_groupi_n_4973 ,csa_tree_add_51_79_groupi_n_6258);
  xnor csa_tree_add_51_79_groupi_g38796(csa_tree_add_51_79_groupi_n_7361 ,csa_tree_add_51_79_groupi_n_4794 ,csa_tree_add_51_79_groupi_n_6257);
  xnor csa_tree_add_51_79_groupi_g38797(csa_tree_add_51_79_groupi_n_7360 ,csa_tree_add_51_79_groupi_n_4835 ,csa_tree_add_51_79_groupi_n_6255);
  xnor csa_tree_add_51_79_groupi_g38798(csa_tree_add_51_79_groupi_n_7359 ,csa_tree_add_51_79_groupi_n_3794 ,csa_tree_add_51_79_groupi_n_6192);
  xnor csa_tree_add_51_79_groupi_g38799(csa_tree_add_51_79_groupi_n_7358 ,csa_tree_add_51_79_groupi_n_4805 ,csa_tree_add_51_79_groupi_n_6252);
  xnor csa_tree_add_51_79_groupi_g38800(csa_tree_add_51_79_groupi_n_7357 ,csa_tree_add_51_79_groupi_n_5087 ,csa_tree_add_51_79_groupi_n_6206);
  xnor csa_tree_add_51_79_groupi_g38801(csa_tree_add_51_79_groupi_n_7356 ,csa_tree_add_51_79_groupi_n_5012 ,csa_tree_add_51_79_groupi_n_6182);
  xnor csa_tree_add_51_79_groupi_g38802(csa_tree_add_51_79_groupi_n_7355 ,csa_tree_add_51_79_groupi_n_5025 ,csa_tree_add_51_79_groupi_n_6165);
  xnor csa_tree_add_51_79_groupi_g38803(csa_tree_add_51_79_groupi_n_7354 ,csa_tree_add_51_79_groupi_n_5023 ,csa_tree_add_51_79_groupi_n_6357);
  xnor csa_tree_add_51_79_groupi_g38804(csa_tree_add_51_79_groupi_n_7353 ,csa_tree_add_51_79_groupi_n_5014 ,csa_tree_add_51_79_groupi_n_6374);
  xnor csa_tree_add_51_79_groupi_g38805(csa_tree_add_51_79_groupi_n_7352 ,csa_tree_add_51_79_groupi_n_5079 ,csa_tree_add_51_79_groupi_n_6380);
  xnor csa_tree_add_51_79_groupi_g38806(csa_tree_add_51_79_groupi_n_7350 ,csa_tree_add_51_79_groupi_n_4946 ,csa_tree_add_51_79_groupi_n_6243);
  xnor csa_tree_add_51_79_groupi_g38807(csa_tree_add_51_79_groupi_n_7349 ,csa_tree_add_51_79_groupi_n_3269 ,csa_tree_add_51_79_groupi_n_6159);
  xnor csa_tree_add_51_79_groupi_g38808(csa_tree_add_51_79_groupi_n_7348 ,csa_tree_add_51_79_groupi_n_5554 ,csa_tree_add_51_79_groupi_n_6364);
  xnor csa_tree_add_51_79_groupi_g38809(csa_tree_add_51_79_groupi_n_7347 ,csa_tree_add_51_79_groupi_n_3765 ,csa_tree_add_51_79_groupi_n_6217);
  xnor csa_tree_add_51_79_groupi_g38810(csa_tree_add_51_79_groupi_n_7345 ,csa_tree_add_51_79_groupi_n_4942 ,csa_tree_add_51_79_groupi_n_6229);
  xnor csa_tree_add_51_79_groupi_g38811(csa_tree_add_51_79_groupi_n_7344 ,csa_tree_add_51_79_groupi_n_5432 ,csa_tree_add_51_79_groupi_n_6239);
  xnor csa_tree_add_51_79_groupi_g38812(csa_tree_add_51_79_groupi_n_7343 ,csa_tree_add_51_79_groupi_n_3783 ,csa_tree_add_51_79_groupi_n_6204);
  xnor csa_tree_add_51_79_groupi_g38813(csa_tree_add_51_79_groupi_n_7342 ,csa_tree_add_51_79_groupi_n_5350 ,csa_tree_add_51_79_groupi_n_6230);
  xnor csa_tree_add_51_79_groupi_g38814(csa_tree_add_51_79_groupi_n_7341 ,csa_tree_add_51_79_groupi_n_5411 ,csa_tree_add_51_79_groupi_n_6227);
  xnor csa_tree_add_51_79_groupi_g38815(csa_tree_add_51_79_groupi_n_7340 ,csa_tree_add_51_79_groupi_n_4815 ,csa_tree_add_51_79_groupi_n_6226);
  xnor csa_tree_add_51_79_groupi_g38816(csa_tree_add_51_79_groupi_n_7339 ,csa_tree_add_51_79_groupi_n_5066 ,csa_tree_add_51_79_groupi_n_6222);
  xnor csa_tree_add_51_79_groupi_g38817(csa_tree_add_51_79_groupi_n_7338 ,csa_tree_add_51_79_groupi_n_5052 ,csa_tree_add_51_79_groupi_n_6218);
  xnor csa_tree_add_51_79_groupi_g38818(csa_tree_add_51_79_groupi_n_7337 ,csa_tree_add_51_79_groupi_n_4949 ,csa_tree_add_51_79_groupi_n_6210);
  xnor csa_tree_add_51_79_groupi_g38819(csa_tree_add_51_79_groupi_n_7336 ,csa_tree_add_51_79_groupi_n_3778 ,csa_tree_add_51_79_groupi_n_6381);
  xnor csa_tree_add_51_79_groupi_g38820(csa_tree_add_51_79_groupi_n_7335 ,csa_tree_add_51_79_groupi_n_5572 ,csa_tree_add_51_79_groupi_n_6249);
  xnor csa_tree_add_51_79_groupi_g38821(csa_tree_add_51_79_groupi_n_7334 ,csa_tree_add_51_79_groupi_n_5480 ,csa_tree_add_51_79_groupi_n_6238);
  xnor csa_tree_add_51_79_groupi_g38822(csa_tree_add_51_79_groupi_n_7333 ,csa_tree_add_51_79_groupi_n_4939 ,csa_tree_add_51_79_groupi_n_6168);
  xnor csa_tree_add_51_79_groupi_g38823(csa_tree_add_51_79_groupi_n_7332 ,csa_tree_add_51_79_groupi_n_3827 ,csa_tree_add_51_79_groupi_n_6376);
  xnor csa_tree_add_51_79_groupi_g38824(csa_tree_add_51_79_groupi_n_7331 ,csa_tree_add_51_79_groupi_n_5576 ,csa_tree_add_51_79_groupi_n_6183);
  xnor csa_tree_add_51_79_groupi_g38825(csa_tree_add_51_79_groupi_n_7330 ,csa_tree_add_51_79_groupi_n_3775 ,csa_tree_add_51_79_groupi_n_6393);
  xnor csa_tree_add_51_79_groupi_g38826(csa_tree_add_51_79_groupi_n_7329 ,csa_tree_add_51_79_groupi_n_3742 ,csa_tree_add_51_79_groupi_n_6354);
  xnor csa_tree_add_51_79_groupi_g38827(csa_tree_add_51_79_groupi_n_7328 ,csa_tree_add_51_79_groupi_n_5324 ,csa_tree_add_51_79_groupi_n_6169);
  xnor csa_tree_add_51_79_groupi_g38828(csa_tree_add_51_79_groupi_n_7327 ,csa_tree_add_51_79_groupi_n_5505 ,csa_tree_add_51_79_groupi_n_6163);
  xnor csa_tree_add_51_79_groupi_g38829(csa_tree_add_51_79_groupi_n_7326 ,csa_tree_add_51_79_groupi_n_5386 ,csa_tree_add_51_79_groupi_n_6171);
  xnor csa_tree_add_51_79_groupi_g38830(csa_tree_add_51_79_groupi_n_7325 ,csa_tree_add_51_79_groupi_n_3246 ,csa_tree_add_51_79_groupi_n_6361);
  xnor csa_tree_add_51_79_groupi_g38831(csa_tree_add_51_79_groupi_n_7324 ,csa_tree_add_51_79_groupi_n_5396 ,csa_tree_add_51_79_groupi_n_6343);
  xnor csa_tree_add_51_79_groupi_g38832(csa_tree_add_51_79_groupi_n_7323 ,csa_tree_add_51_79_groupi_n_5471 ,csa_tree_add_51_79_groupi_n_6233);
  xnor csa_tree_add_51_79_groupi_g38833(csa_tree_add_51_79_groupi_n_7322 ,csa_tree_add_51_79_groupi_n_5385 ,csa_tree_add_51_79_groupi_n_6187);
  xnor csa_tree_add_51_79_groupi_g38834(csa_tree_add_51_79_groupi_n_7321 ,csa_tree_add_51_79_groupi_n_5289 ,csa_tree_add_51_79_groupi_n_6342);
  xnor csa_tree_add_51_79_groupi_g38835(csa_tree_add_51_79_groupi_n_7320 ,csa_tree_add_51_79_groupi_n_5273 ,csa_tree_add_51_79_groupi_n_6323);
  xnor csa_tree_add_51_79_groupi_g38836(csa_tree_add_51_79_groupi_n_7319 ,csa_tree_add_51_79_groupi_n_4711 ,csa_tree_add_51_79_groupi_n_1);
  xnor csa_tree_add_51_79_groupi_g38837(csa_tree_add_51_79_groupi_n_7318 ,csa_tree_add_51_79_groupi_n_5272 ,csa_tree_add_51_79_groupi_n_6368);
  xnor csa_tree_add_51_79_groupi_g38838(csa_tree_add_51_79_groupi_n_7317 ,csa_tree_add_51_79_groupi_n_5482 ,csa_tree_add_51_79_groupi_n_6278);
  xnor csa_tree_add_51_79_groupi_g38839(csa_tree_add_51_79_groupi_n_7316 ,csa_tree_add_51_79_groupi_n_5281 ,csa_tree_add_51_79_groupi_n_6332);
  xnor csa_tree_add_51_79_groupi_g38840(csa_tree_add_51_79_groupi_n_7314 ,csa_tree_add_51_79_groupi_n_5473 ,csa_tree_add_51_79_groupi_n_6281);
  xnor csa_tree_add_51_79_groupi_g38841(csa_tree_add_51_79_groupi_n_7313 ,csa_tree_add_51_79_groupi_n_5456 ,csa_tree_add_51_79_groupi_n_6275);
  xnor csa_tree_add_51_79_groupi_g38842(csa_tree_add_51_79_groupi_n_7311 ,csa_tree_add_51_79_groupi_n_5018 ,csa_tree_add_51_79_groupi_n_6274);
  xnor csa_tree_add_51_79_groupi_g38843(csa_tree_add_51_79_groupi_n_7310 ,csa_tree_add_51_79_groupi_n_5381 ,csa_tree_add_51_79_groupi_n_6358);
  xnor csa_tree_add_51_79_groupi_g38844(csa_tree_add_51_79_groupi_n_7309 ,csa_tree_add_51_79_groupi_n_5070 ,csa_tree_add_51_79_groupi_n_6272);
  xnor csa_tree_add_51_79_groupi_g38845(csa_tree_add_51_79_groupi_n_7308 ,csa_tree_add_51_79_groupi_n_5011 ,csa_tree_add_51_79_groupi_n_6304);
  xnor csa_tree_add_51_79_groupi_g38846(csa_tree_add_51_79_groupi_n_7307 ,csa_tree_add_51_79_groupi_n_5388 ,csa_tree_add_51_79_groupi_n_6344);
  xnor csa_tree_add_51_79_groupi_g38847(csa_tree_add_51_79_groupi_n_7305 ,csa_tree_add_51_79_groupi_n_5436 ,csa_tree_add_51_79_groupi_n_6303);
  xnor csa_tree_add_51_79_groupi_g38848(csa_tree_add_51_79_groupi_n_7304 ,csa_tree_add_51_79_groupi_n_5490 ,csa_tree_add_51_79_groupi_n_6355);
  xnor csa_tree_add_51_79_groupi_g38849(csa_tree_add_51_79_groupi_n_7302 ,csa_tree_add_51_79_groupi_n_5053 ,csa_tree_add_51_79_groupi_n_6268);
  xnor csa_tree_add_51_79_groupi_g38850(csa_tree_add_51_79_groupi_n_7300 ,csa_tree_add_51_79_groupi_n_6151 ,csa_tree_add_51_79_groupi_n_1);
  xnor csa_tree_add_51_79_groupi_g38851(csa_tree_add_51_79_groupi_n_7299 ,csa_tree_add_51_79_groupi_n_5050 ,csa_tree_add_51_79_groupi_n_6267);
  xnor csa_tree_add_51_79_groupi_g38852(csa_tree_add_51_79_groupi_n_7298 ,csa_tree_add_51_79_groupi_n_5048 ,csa_tree_add_51_79_groupi_n_6266);
  xnor csa_tree_add_51_79_groupi_g38854(csa_tree_add_51_79_groupi_n_7297 ,csa_tree_add_51_79_groupi_n_5056 ,csa_tree_add_51_79_groupi_n_6314);
  xnor csa_tree_add_51_79_groupi_g38855(csa_tree_add_51_79_groupi_n_7296 ,csa_tree_add_51_79_groupi_n_5543 ,csa_tree_add_51_79_groupi_n_6353);
  xnor csa_tree_add_51_79_groupi_g38856(csa_tree_add_51_79_groupi_n_7295 ,csa_tree_add_51_79_groupi_n_5064 ,csa_tree_add_51_79_groupi_n_6263);
  xnor csa_tree_add_51_79_groupi_g38857(csa_tree_add_51_79_groupi_n_7294 ,csa_tree_add_51_79_groupi_n_5082 ,csa_tree_add_51_79_groupi_n_6262);
  xnor csa_tree_add_51_79_groupi_g38858(csa_tree_add_51_79_groupi_n_7293 ,csa_tree_add_51_79_groupi_n_5030 ,csa_tree_add_51_79_groupi_n_6362);
  xnor csa_tree_add_51_79_groupi_g38859(csa_tree_add_51_79_groupi_n_7290 ,csa_tree_add_51_79_groupi_n_5466 ,csa_tree_add_51_79_groupi_n_6352);
  xnor csa_tree_add_51_79_groupi_g38860(csa_tree_add_51_79_groupi_n_7289 ,csa_tree_add_51_79_groupi_n_5564 ,csa_tree_add_51_79_groupi_n_6346);
  xnor csa_tree_add_51_79_groupi_g38861(csa_tree_add_51_79_groupi_n_7287 ,csa_tree_add_51_79_groupi_n_3769 ,csa_tree_add_51_79_groupi_n_6202);
  xnor csa_tree_add_51_79_groupi_g38862(csa_tree_add_51_79_groupi_n_7285 ,csa_tree_add_51_79_groupi_n_4978 ,csa_tree_add_51_79_groupi_n_6254);
  xnor csa_tree_add_51_79_groupi_g38863(csa_tree_add_51_79_groupi_n_7284 ,csa_tree_add_51_79_groupi_n_4842 ,csa_tree_add_51_79_groupi_n_6256);
  xnor csa_tree_add_51_79_groupi_g38864(csa_tree_add_51_79_groupi_n_7283 ,csa_tree_add_51_79_groupi_n_5106 ,csa_tree_add_51_79_groupi_n_6322);
  xnor csa_tree_add_51_79_groupi_g38865(csa_tree_add_51_79_groupi_n_7282 ,csa_tree_add_51_79_groupi_n_4921 ,csa_tree_add_51_79_groupi_n_6328);
  xnor csa_tree_add_51_79_groupi_g38866(csa_tree_add_51_79_groupi_n_7281 ,csa_tree_add_51_79_groupi_n_4817 ,csa_tree_add_51_79_groupi_n_6253);
  xnor csa_tree_add_51_79_groupi_g38867(csa_tree_add_51_79_groupi_n_7280 ,csa_tree_add_51_79_groupi_n_4846 ,csa_tree_add_51_79_groupi_n_6320);
  xnor csa_tree_add_51_79_groupi_g38868(csa_tree_add_51_79_groupi_n_7279 ,csa_tree_add_51_79_groupi_n_5039 ,csa_tree_add_51_79_groupi_n_6260);
  xnor csa_tree_add_51_79_groupi_g38869(csa_tree_add_51_79_groupi_n_7278 ,csa_tree_add_51_79_groupi_n_5004 ,csa_tree_add_51_79_groupi_n_6228);
  xnor csa_tree_add_51_79_groupi_g38870(csa_tree_add_51_79_groupi_n_7277 ,csa_tree_add_51_79_groupi_n_5083 ,csa_tree_add_51_79_groupi_n_6213);
  xnor csa_tree_add_51_79_groupi_g38871(csa_tree_add_51_79_groupi_n_7276 ,csa_tree_add_51_79_groupi_n_5037 ,csa_tree_add_51_79_groupi_n_6236);
  xnor csa_tree_add_51_79_groupi_g38872(csa_tree_add_51_79_groupi_n_7275 ,csa_tree_add_51_79_groupi_n_5179 ,csa_tree_add_51_79_groupi_n_6189);
  xnor csa_tree_add_51_79_groupi_g38873(csa_tree_add_51_79_groupi_n_7273 ,csa_tree_add_51_79_groupi_n_5072 ,csa_tree_add_51_79_groupi_n_6198);
  xnor csa_tree_add_51_79_groupi_g38874(csa_tree_add_51_79_groupi_n_7272 ,csa_tree_add_51_79_groupi_n_5088 ,csa_tree_add_51_79_groupi_n_6280);
  xnor csa_tree_add_51_79_groupi_g38875(csa_tree_add_51_79_groupi_n_7271 ,csa_tree_add_51_79_groupi_n_5016 ,csa_tree_add_51_79_groupi_n_6177);
  xnor csa_tree_add_51_79_groupi_g38876(csa_tree_add_51_79_groupi_n_7270 ,csa_tree_add_51_79_groupi_n_5015 ,csa_tree_add_51_79_groupi_n_6167);
  xnor csa_tree_add_51_79_groupi_g38877(csa_tree_add_51_79_groupi_n_7269 ,csa_tree_add_51_79_groupi_n_5019 ,csa_tree_add_51_79_groupi_n_6166);
  xnor csa_tree_add_51_79_groupi_g38878(csa_tree_add_51_79_groupi_n_7268 ,csa_tree_add_51_79_groupi_n_5306 ,csa_tree_add_51_79_groupi_n_6340);
  xnor csa_tree_add_51_79_groupi_g38879(csa_tree_add_51_79_groupi_n_7266 ,csa_tree_add_51_79_groupi_n_5020 ,csa_tree_add_51_79_groupi_n_6164);
  xnor csa_tree_add_51_79_groupi_g38880(csa_tree_add_51_79_groupi_n_7265 ,csa_tree_add_51_79_groupi_n_5041 ,csa_tree_add_51_79_groupi_n_6334);
  xnor csa_tree_add_51_79_groupi_g38881(csa_tree_add_51_79_groupi_n_7264 ,csa_tree_add_51_79_groupi_n_5036 ,csa_tree_add_51_79_groupi_n_6325);
  xnor csa_tree_add_51_79_groupi_g38882(csa_tree_add_51_79_groupi_n_7263 ,csa_tree_add_51_79_groupi_n_5090 ,csa_tree_add_51_79_groupi_n_6317);
  xnor csa_tree_add_51_79_groupi_g38883(csa_tree_add_51_79_groupi_n_7262 ,csa_tree_add_51_79_groupi_n_5031 ,csa_tree_add_51_79_groupi_n_6369);
  xnor csa_tree_add_51_79_groupi_g38884(csa_tree_add_51_79_groupi_n_7260 ,csa_tree_add_51_79_groupi_n_5069 ,csa_tree_add_51_79_groupi_n_6241);
  xnor csa_tree_add_51_79_groupi_g38885(csa_tree_add_51_79_groupi_n_7259 ,csa_tree_add_51_79_groupi_n_5032 ,csa_tree_add_51_79_groupi_n_6246);
  xnor csa_tree_add_51_79_groupi_g38886(csa_tree_add_51_79_groupi_n_7258 ,csa_tree_add_51_79_groupi_n_5081 ,csa_tree_add_51_79_groupi_n_6277);
  xnor csa_tree_add_51_79_groupi_g38887(csa_tree_add_51_79_groupi_n_7257 ,csa_tree_add_51_79_groupi_n_4966 ,csa_tree_add_51_79_groupi_n_6316);
  xnor csa_tree_add_51_79_groupi_g38888(csa_tree_add_51_79_groupi_n_7256 ,csa_tree_add_51_79_groupi_n_5476 ,csa_tree_add_51_79_groupi_n_6338);
  xnor csa_tree_add_51_79_groupi_g38889(csa_tree_add_51_79_groupi_n_7254 ,csa_tree_add_51_79_groupi_n_5111 ,csa_tree_add_51_79_groupi_n_6313);
  xnor csa_tree_add_51_79_groupi_g38890(csa_tree_add_51_79_groupi_n_7253 ,csa_tree_add_51_79_groupi_n_5570 ,csa_tree_add_51_79_groupi_n_6312);
  xnor csa_tree_add_51_79_groupi_g38891(csa_tree_add_51_79_groupi_n_7252 ,csa_tree_add_51_79_groupi_n_5488 ,csa_tree_add_51_79_groupi_n_6305);
  xnor csa_tree_add_51_79_groupi_g38892(csa_tree_add_51_79_groupi_n_7251 ,csa_tree_add_51_79_groupi_n_3740 ,csa_tree_add_51_79_groupi_n_6385);
  xnor csa_tree_add_51_79_groupi_g38893(csa_tree_add_51_79_groupi_n_7249 ,csa_tree_add_51_79_groupi_n_24 ,csa_tree_add_51_79_groupi_n_6326);
  xnor csa_tree_add_51_79_groupi_g38894(csa_tree_add_51_79_groupi_n_7248 ,csa_tree_add_51_79_groupi_n_5574 ,csa_tree_add_51_79_groupi_n_6293);
  xnor csa_tree_add_51_79_groupi_g38895(csa_tree_add_51_79_groupi_n_7247 ,csa_tree_add_51_79_groupi_n_3810 ,csa_tree_add_51_79_groupi_n_6184);
  xnor csa_tree_add_51_79_groupi_g38896(csa_tree_add_51_79_groupi_n_7245 ,csa_tree_add_51_79_groupi_n_5013 ,csa_tree_add_51_79_groupi_n_6299);
  xnor csa_tree_add_51_79_groupi_g38897(csa_tree_add_51_79_groupi_n_7244 ,csa_tree_add_51_79_groupi_n_3300 ,csa_tree_add_51_79_groupi_n_6341);
  xnor csa_tree_add_51_79_groupi_g38898(csa_tree_add_51_79_groupi_n_7242 ,csa_tree_add_51_79_groupi_n_5442 ,csa_tree_add_51_79_groupi_n_6308);
  xnor csa_tree_add_51_79_groupi_g38899(csa_tree_add_51_79_groupi_n_7241 ,csa_tree_add_51_79_groupi_n_5060 ,csa_tree_add_51_79_groupi_n_6264);
  xnor csa_tree_add_51_79_groupi_g38900(csa_tree_add_51_79_groupi_n_7240 ,csa_tree_add_51_79_groupi_n_5317 ,csa_tree_add_51_79_groupi_n_6390);
  xnor csa_tree_add_51_79_groupi_g38901(csa_tree_add_51_79_groupi_n_7238 ,csa_tree_add_51_79_groupi_n_4912 ,csa_tree_add_51_79_groupi_n_6223);
  xnor csa_tree_add_51_79_groupi_g38902(csa_tree_add_51_79_groupi_n_7237 ,csa_tree_add_51_79_groupi_n_5492 ,csa_tree_add_51_79_groupi_n_6283);
  xnor csa_tree_add_51_79_groupi_g38903(csa_tree_add_51_79_groupi_n_7236 ,csa_tree_add_51_79_groupi_n_3750 ,csa_tree_add_51_79_groupi_n_6387);
  xnor csa_tree_add_51_79_groupi_g38904(csa_tree_add_51_79_groupi_n_7235 ,csa_tree_add_51_79_groupi_n_4820 ,csa_tree_add_51_79_groupi_n_6220);
  xnor csa_tree_add_51_79_groupi_g38905(csa_tree_add_51_79_groupi_n_7233 ,csa_tree_add_51_79_groupi_n_5512 ,csa_tree_add_51_79_groupi_n_6291);
  xnor csa_tree_add_51_79_groupi_g38906(csa_tree_add_51_79_groupi_n_7232 ,csa_tree_add_51_79_groupi_n_4878 ,csa_tree_add_51_79_groupi_n_6216);
  xnor csa_tree_add_51_79_groupi_g38907(csa_tree_add_51_79_groupi_n_7230 ,csa_tree_add_51_79_groupi_n_4875 ,csa_tree_add_51_79_groupi_n_6212);
  xnor csa_tree_add_51_79_groupi_g38908(csa_tree_add_51_79_groupi_n_7229 ,csa_tree_add_51_79_groupi_n_4954 ,csa_tree_add_51_79_groupi_n_6205);
  xnor csa_tree_add_51_79_groupi_g38909(csa_tree_add_51_79_groupi_n_7228 ,csa_tree_add_51_79_groupi_n_4950 ,csa_tree_add_51_79_groupi_n_6211);
  xnor csa_tree_add_51_79_groupi_g38910(csa_tree_add_51_79_groupi_n_7227 ,csa_tree_add_51_79_groupi_n_5470 ,csa_tree_add_51_79_groupi_n_6294);
  xnor csa_tree_add_51_79_groupi_g38911(csa_tree_add_51_79_groupi_n_7226 ,csa_tree_add_51_79_groupi_n_5118 ,csa_tree_add_51_79_groupi_n_6215);
  xnor csa_tree_add_51_79_groupi_g38912(csa_tree_add_51_79_groupi_n_7225 ,csa_tree_add_51_79_groupi_n_4871 ,csa_tree_add_51_79_groupi_n_6209);
  xnor csa_tree_add_51_79_groupi_g38913(csa_tree_add_51_79_groupi_n_7224 ,csa_tree_add_51_79_groupi_n_4930 ,csa_tree_add_51_79_groupi_n_6208);
  xnor csa_tree_add_51_79_groupi_g38914(csa_tree_add_51_79_groupi_n_7223 ,csa_tree_add_51_79_groupi_n_5084 ,csa_tree_add_51_79_groupi_n_6207);
  xnor csa_tree_add_51_79_groupi_g38915(csa_tree_add_51_79_groupi_n_7222 ,csa_tree_add_51_79_groupi_n_5449 ,csa_tree_add_51_79_groupi_n_6200);
  xnor csa_tree_add_51_79_groupi_g38916(csa_tree_add_51_79_groupi_n_7221 ,csa_tree_add_51_79_groupi_n_5468 ,csa_tree_add_51_79_groupi_n_6199);
  xnor csa_tree_add_51_79_groupi_g38917(csa_tree_add_51_79_groupi_n_7220 ,csa_tree_add_51_79_groupi_n_5502 ,csa_tree_add_51_79_groupi_n_6302);
  xnor csa_tree_add_51_79_groupi_g38918(csa_tree_add_51_79_groupi_n_7219 ,csa_tree_add_51_79_groupi_n_5229 ,csa_tree_add_51_79_groupi_n_6336);
  xnor csa_tree_add_51_79_groupi_g38919(csa_tree_add_51_79_groupi_n_7217 ,csa_tree_add_51_79_groupi_n_5098 ,csa_tree_add_51_79_groupi_n_6197);
  xnor csa_tree_add_51_79_groupi_g38920(csa_tree_add_51_79_groupi_n_7215 ,csa_tree_add_51_79_groupi_n_5417 ,csa_tree_add_51_79_groupi_n_6231);
  xnor csa_tree_add_51_79_groupi_g38921(csa_tree_add_51_79_groupi_n_7213 ,csa_tree_add_51_79_groupi_n_5017 ,csa_tree_add_51_79_groupi_n_6298);
  xnor csa_tree_add_51_79_groupi_g38922(csa_tree_add_51_79_groupi_n_7212 ,csa_tree_add_51_79_groupi_n_5514 ,csa_tree_add_51_79_groupi_n_6196);
  xnor csa_tree_add_51_79_groupi_g38923(csa_tree_add_51_79_groupi_n_7211 ,csa_tree_add_51_79_groupi_n_5465 ,csa_tree_add_51_79_groupi_n_6193);
  xnor csa_tree_add_51_79_groupi_g38924(csa_tree_add_51_79_groupi_n_7210 ,csa_tree_add_51_79_groupi_n_5550 ,csa_tree_add_51_79_groupi_n_6276);
  xnor csa_tree_add_51_79_groupi_g38925(csa_tree_add_51_79_groupi_n_7209 ,csa_tree_add_51_79_groupi_n_4844 ,csa_tree_add_51_79_groupi_n_6190);
  xnor csa_tree_add_51_79_groupi_g38926(csa_tree_add_51_79_groupi_n_7207 ,csa_tree_add_51_79_groupi_n_5568 ,csa_tree_add_51_79_groupi_n_6185);
  xnor csa_tree_add_51_79_groupi_g38928(csa_tree_add_51_79_groupi_n_7205 ,csa_tree_add_51_79_groupi_n_5540 ,csa_tree_add_51_79_groupi_n_6176);
  xnor csa_tree_add_51_79_groupi_g38929(csa_tree_add_51_79_groupi_n_7204 ,csa_tree_add_51_79_groupi_n_5548 ,csa_tree_add_51_79_groupi_n_6175);
  xnor csa_tree_add_51_79_groupi_g38930(csa_tree_add_51_79_groupi_n_7203 ,csa_tree_add_51_79_groupi_n_5527 ,csa_tree_add_51_79_groupi_n_6270);
  xnor csa_tree_add_51_79_groupi_g38931(csa_tree_add_51_79_groupi_n_7202 ,csa_tree_add_51_79_groupi_n_5535 ,csa_tree_add_51_79_groupi_n_6174);
  xnor csa_tree_add_51_79_groupi_g38932(csa_tree_add_51_79_groupi_n_7201 ,csa_tree_add_51_79_groupi_n_5547 ,csa_tree_add_51_79_groupi_n_6247);
  xnor csa_tree_add_51_79_groupi_g38933(csa_tree_add_51_79_groupi_n_7200 ,csa_tree_add_51_79_groupi_n_5215 ,csa_tree_add_51_79_groupi_n_6173);
  xnor csa_tree_add_51_79_groupi_g38934(csa_tree_add_51_79_groupi_n_7199 ,csa_tree_add_51_79_groupi_n_5537 ,csa_tree_add_51_79_groupi_n_6172);
  xnor csa_tree_add_51_79_groupi_g38935(csa_tree_add_51_79_groupi_n_7198 ,csa_tree_add_51_79_groupi_n_5372 ,csa_tree_add_51_79_groupi_n_6330);
  xnor csa_tree_add_51_79_groupi_g38936(csa_tree_add_51_79_groupi_n_7196 ,csa_tree_add_51_79_groupi_n_5251 ,csa_tree_add_51_79_groupi_n_6240);
  xnor csa_tree_add_51_79_groupi_g38937(csa_tree_add_51_79_groupi_n_7194 ,csa_tree_add_51_79_groupi_n_5325 ,csa_tree_add_51_79_groupi_n_6162);
  xnor csa_tree_add_51_79_groupi_g38938(csa_tree_add_51_79_groupi_n_7192 ,csa_tree_add_51_79_groupi_n_4861 ,csa_tree_add_51_79_groupi_n_6170);
  xnor csa_tree_add_51_79_groupi_g38939(csa_tree_add_51_79_groupi_n_7191 ,csa_tree_add_51_79_groupi_n_5552 ,csa_tree_add_51_79_groupi_n_6306);
  xnor csa_tree_add_51_79_groupi_g38940(csa_tree_add_51_79_groupi_n_7190 ,csa_tree_add_51_79_groupi_n_5486 ,csa_tree_add_51_79_groupi_n_6356);
  xnor csa_tree_add_51_79_groupi_g38941(csa_tree_add_51_79_groupi_n_7189 ,csa_tree_add_51_79_groupi_n_3306 ,csa_tree_add_51_79_groupi_n_6234);
  xnor csa_tree_add_51_79_groupi_g38942(csa_tree_add_51_79_groupi_n_7187 ,csa_tree_add_51_79_groupi_n_5413 ,csa_tree_add_51_79_groupi_n_6160);
  xnor csa_tree_add_51_79_groupi_g38943(csa_tree_add_51_79_groupi_n_7185 ,csa_tree_add_51_79_groupi_n_5489 ,csa_tree_add_51_79_groupi_n_6157);
  xnor csa_tree_add_51_79_groupi_g38944(csa_tree_add_51_79_groupi_n_7183 ,csa_tree_add_51_79_groupi_n_5344 ,csa_tree_add_51_79_groupi_n_6245);
  xnor csa_tree_add_51_79_groupi_g38945(csa_tree_add_51_79_groupi_n_7182 ,csa_tree_add_51_79_groupi_n_5507 ,csa_tree_add_51_79_groupi_n_6284);
  xnor csa_tree_add_51_79_groupi_g38946(csa_tree_add_51_79_groupi_n_7181 ,csa_tree_add_51_79_groupi_n_5529 ,csa_tree_add_51_79_groupi_n_6158);
  xnor csa_tree_add_51_79_groupi_g38947(csa_tree_add_51_79_groupi_n_7179 ,csa_tree_add_51_79_groupi_n_5282 ,csa_tree_add_51_79_groupi_n_6186);
  xnor csa_tree_add_51_79_groupi_g38948(csa_tree_add_51_79_groupi_n_7177 ,csa_tree_add_51_79_groupi_n_5027 ,csa_tree_add_51_79_groupi_n_6363);
  xnor csa_tree_add_51_79_groupi_g38949(csa_tree_add_51_79_groupi_n_7176 ,csa_tree_add_51_79_groupi_n_4976 ,csa_tree_add_51_79_groupi_n_6221);
  xnor csa_tree_add_51_79_groupi_g38950(csa_tree_add_51_79_groupi_n_7175 ,csa_tree_add_51_79_groupi_n_5116 ,csa_tree_add_51_79_groupi_n_6329);
  xnor csa_tree_add_51_79_groupi_g38951(csa_tree_add_51_79_groupi_n_7173 ,csa_tree_add_51_79_groupi_n_5024 ,csa_tree_add_51_79_groupi_n_6289);
  xnor csa_tree_add_51_79_groupi_g38952(csa_tree_add_51_79_groupi_n_7172 ,csa_tree_add_51_79_groupi_n_5028 ,csa_tree_add_51_79_groupi_n_6319);
  xnor csa_tree_add_51_79_groupi_g38953(csa_tree_add_51_79_groupi_n_7171 ,csa_tree_add_51_79_groupi_n_5481 ,csa_tree_add_51_79_groupi_n_6232);
  xnor csa_tree_add_51_79_groupi_g38954(csa_tree_add_51_79_groupi_n_7170 ,csa_tree_add_51_79_groupi_n_5504 ,csa_tree_add_51_79_groupi_n_6250);
  xnor csa_tree_add_51_79_groupi_g38955(csa_tree_add_51_79_groupi_n_7168 ,csa_tree_add_51_79_groupi_n_4863 ,csa_tree_add_51_79_groupi_n_6351);
  xnor csa_tree_add_51_79_groupi_g38956(csa_tree_add_51_79_groupi_n_7167 ,csa_tree_add_51_79_groupi_n_5464 ,csa_tree_add_51_79_groupi_n_6242);
  xnor csa_tree_add_51_79_groupi_g38957(csa_tree_add_51_79_groupi_n_7166 ,csa_tree_add_51_79_groupi_n_5440 ,csa_tree_add_51_79_groupi_n_6288);
  xnor csa_tree_add_51_79_groupi_g38958(csa_tree_add_51_79_groupi_n_7165 ,csa_tree_add_51_79_groupi_n_5198 ,csa_tree_add_51_79_groupi_n_6324);
  xnor csa_tree_add_51_79_groupi_g38959(csa_tree_add_51_79_groupi_n_7164 ,csa_tree_add_51_79_groupi_n_5054 ,csa_tree_add_51_79_groupi_n_6331);
  xnor csa_tree_add_51_79_groupi_g38960(csa_tree_add_51_79_groupi_n_7162 ,csa_tree_add_51_79_groupi_n_5043 ,csa_tree_add_51_79_groupi_n_6265);
  xnor csa_tree_add_51_79_groupi_g38961(csa_tree_add_51_79_groupi_n_7161 ,csa_tree_add_51_79_groupi_n_5307 ,csa_tree_add_51_79_groupi_n_6203);
  xnor csa_tree_add_51_79_groupi_g38962(csa_tree_add_51_79_groupi_n_7159 ,csa_tree_add_51_79_groupi_n_5231 ,csa_tree_add_51_79_groupi_n_6178);
  xnor csa_tree_add_51_79_groupi_g38963(csa_tree_add_51_79_groupi_n_7157 ,csa_tree_add_51_79_groupi_n_4968 ,csa_tree_add_51_79_groupi_n_6225);
  xnor csa_tree_add_51_79_groupi_g38964(csa_tree_add_51_79_groupi_n_7155 ,csa_tree_add_51_79_groupi_n_5394 ,csa_tree_add_51_79_groupi_n_6248);
  xnor csa_tree_add_51_79_groupi_g38965(csa_tree_add_51_79_groupi_n_7153 ,csa_tree_add_51_79_groupi_n_5563 ,csa_tree_add_51_79_groupi_n_6335);
  xnor csa_tree_add_51_79_groupi_g38966(csa_tree_add_51_79_groupi_n_7152 ,csa_tree_add_51_79_groupi_n_5462 ,csa_tree_add_51_79_groupi_n_6339);
  xnor csa_tree_add_51_79_groupi_g38967(csa_tree_add_51_79_groupi_n_7151 ,csa_tree_add_51_79_groupi_n_5493 ,csa_tree_add_51_79_groupi_n_6348);
  xnor csa_tree_add_51_79_groupi_g38968(csa_tree_add_51_79_groupi_n_7150 ,csa_tree_add_51_79_groupi_n_4801 ,csa_tree_add_51_79_groupi_n_6347);
  xnor csa_tree_add_51_79_groupi_g38969(csa_tree_add_51_79_groupi_n_7149 ,csa_tree_add_51_79_groupi_n_5545 ,csa_tree_add_51_79_groupi_n_6349);
  xnor csa_tree_add_51_79_groupi_g38970(csa_tree_add_51_79_groupi_n_7148 ,csa_tree_add_51_79_groupi_n_5329 ,csa_tree_add_51_79_groupi_n_6360);
  xnor csa_tree_add_51_79_groupi_g38971(csa_tree_add_51_79_groupi_n_7147 ,csa_tree_add_51_79_groupi_n_5252 ,csa_tree_add_51_79_groupi_n_6365);
  xnor csa_tree_add_51_79_groupi_g38972(csa_tree_add_51_79_groupi_n_7145 ,csa_tree_add_51_79_groupi_n_5258 ,csa_tree_add_51_79_groupi_n_6327);
  xnor csa_tree_add_51_79_groupi_g38973(csa_tree_add_51_79_groupi_n_7143 ,csa_tree_add_51_79_groupi_n_4830 ,csa_tree_add_51_79_groupi_n_6371);
  xnor csa_tree_add_51_79_groupi_g38974(csa_tree_add_51_79_groupi_n_7142 ,csa_tree_add_51_79_groupi_n_5123 ,csa_tree_add_51_79_groupi_n_6372);
  xnor csa_tree_add_51_79_groupi_g38975(csa_tree_add_51_79_groupi_n_7141 ,csa_tree_add_51_79_groupi_n_4831 ,csa_tree_add_51_79_groupi_n_6373);
  xnor csa_tree_add_51_79_groupi_g38976(csa_tree_add_51_79_groupi_n_7140 ,csa_tree_add_51_79_groupi_n_5298 ,csa_tree_add_51_79_groupi_n_6375);
  xnor csa_tree_add_51_79_groupi_g38977(csa_tree_add_51_79_groupi_n_7139 ,csa_tree_add_51_79_groupi_n_5295 ,csa_tree_add_51_79_groupi_n_6391);
  xnor csa_tree_add_51_79_groupi_g38978(csa_tree_add_51_79_groupi_n_7137 ,csa_tree_add_51_79_groupi_n_3281 ,csa_tree_add_51_79_groupi_n_6345);
  not csa_tree_add_51_79_groupi_g38979(csa_tree_add_51_79_groupi_n_7103 ,csa_tree_add_51_79_groupi_n_7102);
  not csa_tree_add_51_79_groupi_g38980(csa_tree_add_51_79_groupi_n_7075 ,csa_tree_add_51_79_groupi_n_7074);
  not csa_tree_add_51_79_groupi_g38981(csa_tree_add_51_79_groupi_n_7055 ,csa_tree_add_51_79_groupi_n_7056);
  not csa_tree_add_51_79_groupi_g38982(csa_tree_add_51_79_groupi_n_7045 ,csa_tree_add_51_79_groupi_n_7046);
  not csa_tree_add_51_79_groupi_g38983(csa_tree_add_51_79_groupi_n_7041 ,csa_tree_add_51_79_groupi_n_7042);
  not csa_tree_add_51_79_groupi_g38984(csa_tree_add_51_79_groupi_n_7036 ,csa_tree_add_51_79_groupi_n_7035);
  not csa_tree_add_51_79_groupi_g38985(csa_tree_add_51_79_groupi_n_7024 ,csa_tree_add_51_79_groupi_n_7025);
  not csa_tree_add_51_79_groupi_g38986(csa_tree_add_51_79_groupi_n_7011 ,csa_tree_add_51_79_groupi_n_7012);
  not csa_tree_add_51_79_groupi_g38987(csa_tree_add_51_79_groupi_n_7009 ,csa_tree_add_51_79_groupi_n_7010);
  not csa_tree_add_51_79_groupi_g38988(csa_tree_add_51_79_groupi_n_7007 ,csa_tree_add_51_79_groupi_n_7008);
  not csa_tree_add_51_79_groupi_g38989(csa_tree_add_51_79_groupi_n_7002 ,csa_tree_add_51_79_groupi_n_7003);
  not csa_tree_add_51_79_groupi_g38990(csa_tree_add_51_79_groupi_n_6996 ,csa_tree_add_51_79_groupi_n_6997);
  not csa_tree_add_51_79_groupi_g38991(csa_tree_add_51_79_groupi_n_6987 ,csa_tree_add_51_79_groupi_n_6988);
  not csa_tree_add_51_79_groupi_g38992(csa_tree_add_51_79_groupi_n_6984 ,csa_tree_add_51_79_groupi_n_6985);
  not csa_tree_add_51_79_groupi_g38993(csa_tree_add_51_79_groupi_n_6980 ,csa_tree_add_51_79_groupi_n_6981);
  not csa_tree_add_51_79_groupi_g38994(csa_tree_add_51_79_groupi_n_6960 ,csa_tree_add_51_79_groupi_n_6961);
  and csa_tree_add_51_79_groupi_g38995(csa_tree_add_51_79_groupi_n_6959 ,csa_tree_add_51_79_groupi_n_6631 ,csa_tree_add_51_79_groupi_n_6452);
  or csa_tree_add_51_79_groupi_g38996(csa_tree_add_51_79_groupi_n_6958 ,csa_tree_add_51_79_groupi_n_6753 ,csa_tree_add_51_79_groupi_n_6449);
  or csa_tree_add_51_79_groupi_g38997(csa_tree_add_51_79_groupi_n_6957 ,csa_tree_add_51_79_groupi_n_6127 ,csa_tree_add_51_79_groupi_n_6413);
  and csa_tree_add_51_79_groupi_g38998(csa_tree_add_51_79_groupi_n_6956 ,csa_tree_add_51_79_groupi_n_6443 ,csa_tree_add_51_79_groupi_n_6444);
  or csa_tree_add_51_79_groupi_g38999(csa_tree_add_51_79_groupi_n_6955 ,csa_tree_add_51_79_groupi_n_6443 ,csa_tree_add_51_79_groupi_n_6444);
  and csa_tree_add_51_79_groupi_g39000(csa_tree_add_51_79_groupi_n_6954 ,csa_tree_add_51_79_groupi_n_6608 ,csa_tree_add_51_79_groupi_n_6451);
  and csa_tree_add_51_79_groupi_g39001(csa_tree_add_51_79_groupi_n_6953 ,csa_tree_add_51_79_groupi_n_6127 ,csa_tree_add_51_79_groupi_n_6413);
  nor csa_tree_add_51_79_groupi_g39002(csa_tree_add_51_79_groupi_n_6952 ,csa_tree_add_51_79_groupi_n_4804 ,csa_tree_add_51_79_groupi_n_6422);
  or csa_tree_add_51_79_groupi_g39003(csa_tree_add_51_79_groupi_n_6951 ,csa_tree_add_51_79_groupi_n_5335 ,csa_tree_add_51_79_groupi_n_6445);
  or csa_tree_add_51_79_groupi_g39004(csa_tree_add_51_79_groupi_n_6950 ,csa_tree_add_51_79_groupi_n_6149 ,csa_tree_add_51_79_groupi_n_6584);
  or csa_tree_add_51_79_groupi_g39005(csa_tree_add_51_79_groupi_n_6949 ,csa_tree_add_51_79_groupi_n_6433 ,csa_tree_add_51_79_groupi_n_6434);
  and csa_tree_add_51_79_groupi_g39006(csa_tree_add_51_79_groupi_n_6948 ,csa_tree_add_51_79_groupi_n_5335 ,csa_tree_add_51_79_groupi_n_6445);
  or csa_tree_add_51_79_groupi_g39007(csa_tree_add_51_79_groupi_n_6947 ,csa_tree_add_51_79_groupi_n_6147 ,csa_tree_add_51_79_groupi_n_6598);
  and csa_tree_add_51_79_groupi_g39008(csa_tree_add_51_79_groupi_n_6946 ,csa_tree_add_51_79_groupi_n_6446 ,csa_tree_add_51_79_groupi_n_6447);
  or csa_tree_add_51_79_groupi_g39009(csa_tree_add_51_79_groupi_n_6945 ,csa_tree_add_51_79_groupi_n_6756 ,csa_tree_add_51_79_groupi_n_6751);
  or csa_tree_add_51_79_groupi_g39010(csa_tree_add_51_79_groupi_n_6944 ,csa_tree_add_51_79_groupi_n_6155 ,csa_tree_add_51_79_groupi_n_6647);
  and csa_tree_add_51_79_groupi_g39011(csa_tree_add_51_79_groupi_n_6943 ,csa_tree_add_51_79_groupi_n_6438 ,csa_tree_add_51_79_groupi_n_6439);
  nor csa_tree_add_51_79_groupi_g39012(csa_tree_add_51_79_groupi_n_6942 ,csa_tree_add_51_79_groupi_n_5279 ,csa_tree_add_51_79_groupi_n_25);
  and csa_tree_add_51_79_groupi_g39013(csa_tree_add_51_79_groupi_n_6941 ,csa_tree_add_51_79_groupi_n_5279 ,csa_tree_add_51_79_groupi_n_25);
  or csa_tree_add_51_79_groupi_g39014(csa_tree_add_51_79_groupi_n_6940 ,csa_tree_add_51_79_groupi_n_6438 ,csa_tree_add_51_79_groupi_n_6439);
  and csa_tree_add_51_79_groupi_g39015(csa_tree_add_51_79_groupi_n_7117 ,csa_tree_add_51_79_groupi_n_5901 ,csa_tree_add_51_79_groupi_n_6600);
  and csa_tree_add_51_79_groupi_g39016(csa_tree_add_51_79_groupi_n_7116 ,csa_tree_add_51_79_groupi_n_6031 ,csa_tree_add_51_79_groupi_n_6675);
  and csa_tree_add_51_79_groupi_g39017(csa_tree_add_51_79_groupi_n_7115 ,csa_tree_add_51_79_groupi_n_6026 ,csa_tree_add_51_79_groupi_n_6671);
  and csa_tree_add_51_79_groupi_g39018(csa_tree_add_51_79_groupi_n_7114 ,csa_tree_add_51_79_groupi_n_6017 ,csa_tree_add_51_79_groupi_n_6636);
  and csa_tree_add_51_79_groupi_g39019(csa_tree_add_51_79_groupi_n_7113 ,csa_tree_add_51_79_groupi_n_6015 ,csa_tree_add_51_79_groupi_n_6664);
  and csa_tree_add_51_79_groupi_g39020(csa_tree_add_51_79_groupi_n_7112 ,csa_tree_add_51_79_groupi_n_6013 ,csa_tree_add_51_79_groupi_n_6665);
  and csa_tree_add_51_79_groupi_g39021(csa_tree_add_51_79_groupi_n_7111 ,csa_tree_add_51_79_groupi_n_6002 ,csa_tree_add_51_79_groupi_n_6659);
  and csa_tree_add_51_79_groupi_g39022(csa_tree_add_51_79_groupi_n_7110 ,csa_tree_add_51_79_groupi_n_5996 ,csa_tree_add_51_79_groupi_n_6656);
  and csa_tree_add_51_79_groupi_g39023(csa_tree_add_51_79_groupi_n_7109 ,csa_tree_add_51_79_groupi_n_5962 ,csa_tree_add_51_79_groupi_n_6654);
  and csa_tree_add_51_79_groupi_g39024(csa_tree_add_51_79_groupi_n_7108 ,csa_tree_add_51_79_groupi_n_5982 ,csa_tree_add_51_79_groupi_n_6650);
  and csa_tree_add_51_79_groupi_g39025(csa_tree_add_51_79_groupi_n_7107 ,csa_tree_add_51_79_groupi_n_5980 ,csa_tree_add_51_79_groupi_n_6648);
  and csa_tree_add_51_79_groupi_g39026(csa_tree_add_51_79_groupi_n_7106 ,csa_tree_add_51_79_groupi_n_6042 ,csa_tree_add_51_79_groupi_n_6681);
  and csa_tree_add_51_79_groupi_g39027(csa_tree_add_51_79_groupi_n_7105 ,csa_tree_add_51_79_groupi_n_5816 ,csa_tree_add_51_79_groupi_n_6642);
  and csa_tree_add_51_79_groupi_g39028(csa_tree_add_51_79_groupi_n_7104 ,csa_tree_add_51_79_groupi_n_5968 ,csa_tree_add_51_79_groupi_n_6635);
  or csa_tree_add_51_79_groupi_g39029(csa_tree_add_51_79_groupi_n_7102 ,csa_tree_add_51_79_groupi_n_5967 ,csa_tree_add_51_79_groupi_n_6640);
  and csa_tree_add_51_79_groupi_g39030(csa_tree_add_51_79_groupi_n_7101 ,csa_tree_add_51_79_groupi_n_5869 ,csa_tree_add_51_79_groupi_n_6670);
  and csa_tree_add_51_79_groupi_g39031(csa_tree_add_51_79_groupi_n_7100 ,csa_tree_add_51_79_groupi_n_5965 ,csa_tree_add_51_79_groupi_n_6683);
  and csa_tree_add_51_79_groupi_g39032(csa_tree_add_51_79_groupi_n_7099 ,csa_tree_add_51_79_groupi_n_5954 ,csa_tree_add_51_79_groupi_n_6629);
  and csa_tree_add_51_79_groupi_g39033(csa_tree_add_51_79_groupi_n_7098 ,csa_tree_add_51_79_groupi_n_6053 ,csa_tree_add_51_79_groupi_n_6686);
  and csa_tree_add_51_79_groupi_g39034(csa_tree_add_51_79_groupi_n_7097 ,csa_tree_add_51_79_groupi_n_5783 ,csa_tree_add_51_79_groupi_n_6627);
  and csa_tree_add_51_79_groupi_g39035(csa_tree_add_51_79_groupi_n_7096 ,csa_tree_add_51_79_groupi_n_5940 ,csa_tree_add_51_79_groupi_n_6622);
  and csa_tree_add_51_79_groupi_g39036(csa_tree_add_51_79_groupi_n_7095 ,csa_tree_add_51_79_groupi_n_5934 ,csa_tree_add_51_79_groupi_n_6618);
  and csa_tree_add_51_79_groupi_g39037(csa_tree_add_51_79_groupi_n_7094 ,csa_tree_add_51_79_groupi_n_5930 ,csa_tree_add_51_79_groupi_n_6617);
  and csa_tree_add_51_79_groupi_g39038(csa_tree_add_51_79_groupi_n_7093 ,csa_tree_add_51_79_groupi_n_5766 ,csa_tree_add_51_79_groupi_n_6615);
  and csa_tree_add_51_79_groupi_g39039(csa_tree_add_51_79_groupi_n_7092 ,csa_tree_add_51_79_groupi_n_5972 ,csa_tree_add_51_79_groupi_n_6611);
  or csa_tree_add_51_79_groupi_g39040(csa_tree_add_51_79_groupi_n_7091 ,csa_tree_add_51_79_groupi_n_5730 ,csa_tree_add_51_79_groupi_n_6601);
  and csa_tree_add_51_79_groupi_g39041(csa_tree_add_51_79_groupi_n_7090 ,csa_tree_add_51_79_groupi_n_5906 ,csa_tree_add_51_79_groupi_n_6602);
  and csa_tree_add_51_79_groupi_g39042(csa_tree_add_51_79_groupi_n_7089 ,csa_tree_add_51_79_groupi_n_6024 ,csa_tree_add_51_79_groupi_n_6660);
  and csa_tree_add_51_79_groupi_g39043(csa_tree_add_51_79_groupi_n_7088 ,csa_tree_add_51_79_groupi_n_6061 ,csa_tree_add_51_79_groupi_n_6691);
  and csa_tree_add_51_79_groupi_g39044(csa_tree_add_51_79_groupi_n_7087 ,csa_tree_add_51_79_groupi_n_5888 ,csa_tree_add_51_79_groupi_n_6591);
  and csa_tree_add_51_79_groupi_g39045(csa_tree_add_51_79_groupi_n_7086 ,csa_tree_add_51_79_groupi_n_5891 ,csa_tree_add_51_79_groupi_n_6595);
  or csa_tree_add_51_79_groupi_g39046(csa_tree_add_51_79_groupi_n_7085 ,csa_tree_add_51_79_groupi_n_6051 ,csa_tree_add_51_79_groupi_n_6680);
  and csa_tree_add_51_79_groupi_g39047(csa_tree_add_51_79_groupi_n_7084 ,csa_tree_add_51_79_groupi_n_5687 ,csa_tree_add_51_79_groupi_n_6557);
  and csa_tree_add_51_79_groupi_g39048(csa_tree_add_51_79_groupi_n_7083 ,csa_tree_add_51_79_groupi_n_5882 ,csa_tree_add_51_79_groupi_n_6590);
  or csa_tree_add_51_79_groupi_g39049(csa_tree_add_51_79_groupi_n_7082 ,csa_tree_add_51_79_groupi_n_5710 ,csa_tree_add_51_79_groupi_n_6493);
  and csa_tree_add_51_79_groupi_g39050(csa_tree_add_51_79_groupi_n_7081 ,csa_tree_add_51_79_groupi_n_5878 ,csa_tree_add_51_79_groupi_n_6589);
  and csa_tree_add_51_79_groupi_g39051(csa_tree_add_51_79_groupi_n_7080 ,csa_tree_add_51_79_groupi_n_6068 ,csa_tree_add_51_79_groupi_n_6695);
  and csa_tree_add_51_79_groupi_g39052(csa_tree_add_51_79_groupi_n_7079 ,csa_tree_add_51_79_groupi_n_5809 ,csa_tree_add_51_79_groupi_n_6582);
  and csa_tree_add_51_79_groupi_g39053(csa_tree_add_51_79_groupi_n_7078 ,csa_tree_add_51_79_groupi_n_6072 ,csa_tree_add_51_79_groupi_n_6696);
  and csa_tree_add_51_79_groupi_g39054(csa_tree_add_51_79_groupi_n_7077 ,csa_tree_add_51_79_groupi_n_6080 ,csa_tree_add_51_79_groupi_n_6700);
  and csa_tree_add_51_79_groupi_g39055(csa_tree_add_51_79_groupi_n_7076 ,csa_tree_add_51_79_groupi_n_5976 ,csa_tree_add_51_79_groupi_n_6718);
  or csa_tree_add_51_79_groupi_g39056(csa_tree_add_51_79_groupi_n_7074 ,csa_tree_add_51_79_groupi_n_5984 ,csa_tree_add_51_79_groupi_n_6576);
  and csa_tree_add_51_79_groupi_g39057(csa_tree_add_51_79_groupi_n_7073 ,csa_tree_add_51_79_groupi_n_6078 ,csa_tree_add_51_79_groupi_n_6575);
  and csa_tree_add_51_79_groupi_g39058(csa_tree_add_51_79_groupi_n_7072 ,csa_tree_add_51_79_groupi_n_5802 ,csa_tree_add_51_79_groupi_n_6572);
  and csa_tree_add_51_79_groupi_g39059(csa_tree_add_51_79_groupi_n_7071 ,csa_tree_add_51_79_groupi_n_6087 ,csa_tree_add_51_79_groupi_n_6701);
  and csa_tree_add_51_79_groupi_g39060(csa_tree_add_51_79_groupi_n_7070 ,csa_tree_add_51_79_groupi_n_5830 ,csa_tree_add_51_79_groupi_n_6569);
  and csa_tree_add_51_79_groupi_g39061(csa_tree_add_51_79_groupi_n_7069 ,csa_tree_add_51_79_groupi_n_6097 ,csa_tree_add_51_79_groupi_n_6708);
  and csa_tree_add_51_79_groupi_g39062(csa_tree_add_51_79_groupi_n_7068 ,csa_tree_add_51_79_groupi_n_5875 ,csa_tree_add_51_79_groupi_n_6563);
  and csa_tree_add_51_79_groupi_g39063(csa_tree_add_51_79_groupi_n_7067 ,csa_tree_add_51_79_groupi_n_5822 ,csa_tree_add_51_79_groupi_n_6561);
  and csa_tree_add_51_79_groupi_g39064(csa_tree_add_51_79_groupi_n_7066 ,csa_tree_add_51_79_groupi_n_6099 ,csa_tree_add_51_79_groupi_n_6705);
  and csa_tree_add_51_79_groupi_g39065(csa_tree_add_51_79_groupi_n_7065 ,csa_tree_add_51_79_groupi_n_5819 ,csa_tree_add_51_79_groupi_n_6558);
  and csa_tree_add_51_79_groupi_g39066(csa_tree_add_51_79_groupi_n_7064 ,csa_tree_add_51_79_groupi_n_6102 ,csa_tree_add_51_79_groupi_n_6709);
  and csa_tree_add_51_79_groupi_g39067(csa_tree_add_51_79_groupi_n_7063 ,csa_tree_add_51_79_groupi_n_5900 ,csa_tree_add_51_79_groupi_n_6556);
  and csa_tree_add_51_79_groupi_g39068(csa_tree_add_51_79_groupi_n_7062 ,csa_tree_add_51_79_groupi_n_5877 ,csa_tree_add_51_79_groupi_n_6478);
  and csa_tree_add_51_79_groupi_g39069(csa_tree_add_51_79_groupi_n_7061 ,csa_tree_add_51_79_groupi_n_6095 ,csa_tree_add_51_79_groupi_n_6704);
  and csa_tree_add_51_79_groupi_g39070(csa_tree_add_51_79_groupi_n_7060 ,csa_tree_add_51_79_groupi_n_6116 ,csa_tree_add_51_79_groupi_n_6644);
  and csa_tree_add_51_79_groupi_g39071(csa_tree_add_51_79_groupi_n_7059 ,csa_tree_add_51_79_groupi_n_5974 ,csa_tree_add_51_79_groupi_n_6643);
  and csa_tree_add_51_79_groupi_g39072(csa_tree_add_51_79_groupi_n_7058 ,csa_tree_add_51_79_groupi_n_6058 ,csa_tree_add_51_79_groupi_n_6690);
  and csa_tree_add_51_79_groupi_g39073(csa_tree_add_51_79_groupi_n_7057 ,csa_tree_add_51_79_groupi_n_6056 ,csa_tree_add_51_79_groupi_n_6688);
  and csa_tree_add_51_79_groupi_g39074(csa_tree_add_51_79_groupi_n_7056 ,csa_tree_add_51_79_groupi_n_6050 ,csa_tree_add_51_79_groupi_n_6682);
  and csa_tree_add_51_79_groupi_g39075(csa_tree_add_51_79_groupi_n_7054 ,csa_tree_add_51_79_groupi_n_5990 ,csa_tree_add_51_79_groupi_n_6555);
  and csa_tree_add_51_79_groupi_g39076(csa_tree_add_51_79_groupi_n_7053 ,csa_tree_add_51_79_groupi_n_6094 ,csa_tree_add_51_79_groupi_n_6706);
  and csa_tree_add_51_79_groupi_g39077(csa_tree_add_51_79_groupi_n_7052 ,csa_tree_add_51_79_groupi_n_5959 ,csa_tree_add_51_79_groupi_n_6633);
  and csa_tree_add_51_79_groupi_g39078(csa_tree_add_51_79_groupi_n_7051 ,csa_tree_add_51_79_groupi_n_5956 ,csa_tree_add_51_79_groupi_n_6630);
  and csa_tree_add_51_79_groupi_g39079(csa_tree_add_51_79_groupi_n_7050 ,csa_tree_add_51_79_groupi_n_6049 ,csa_tree_add_51_79_groupi_n_6685);
  and csa_tree_add_51_79_groupi_g39080(csa_tree_add_51_79_groupi_n_7049 ,csa_tree_add_51_79_groupi_n_6048 ,csa_tree_add_51_79_groupi_n_6684);
  and csa_tree_add_51_79_groupi_g39081(csa_tree_add_51_79_groupi_n_7048 ,csa_tree_add_51_79_groupi_n_6092 ,csa_tree_add_51_79_groupi_n_6703);
  and csa_tree_add_51_79_groupi_g39082(csa_tree_add_51_79_groupi_n_7047 ,csa_tree_add_51_79_groupi_n_6090 ,csa_tree_add_51_79_groupi_n_6702);
  and csa_tree_add_51_79_groupi_g39083(csa_tree_add_51_79_groupi_n_7046 ,csa_tree_add_51_79_groupi_n_5951 ,csa_tree_add_51_79_groupi_n_6626);
  and csa_tree_add_51_79_groupi_g39084(csa_tree_add_51_79_groupi_n_7044 ,csa_tree_add_51_79_groupi_n_5949 ,csa_tree_add_51_79_groupi_n_6625);
  and csa_tree_add_51_79_groupi_g39085(csa_tree_add_51_79_groupi_n_7043 ,csa_tree_add_51_79_groupi_n_5945 ,csa_tree_add_51_79_groupi_n_6624);
  or csa_tree_add_51_79_groupi_g39086(csa_tree_add_51_79_groupi_n_7042 ,csa_tree_add_51_79_groupi_n_5942 ,csa_tree_add_51_79_groupi_n_6623);
  and csa_tree_add_51_79_groupi_g39087(csa_tree_add_51_79_groupi_n_7040 ,csa_tree_add_51_79_groupi_n_5939 ,csa_tree_add_51_79_groupi_n_6620);
  and csa_tree_add_51_79_groupi_g39088(csa_tree_add_51_79_groupi_n_7039 ,csa_tree_add_51_79_groupi_n_5814 ,csa_tree_add_51_79_groupi_n_6510);
  and csa_tree_add_51_79_groupi_g39089(csa_tree_add_51_79_groupi_n_7038 ,csa_tree_add_51_79_groupi_n_5936 ,csa_tree_add_51_79_groupi_n_6610);
  and csa_tree_add_51_79_groupi_g39090(csa_tree_add_51_79_groupi_n_7037 ,csa_tree_add_51_79_groupi_n_5937 ,csa_tree_add_51_79_groupi_n_6621);
  and csa_tree_add_51_79_groupi_g39091(csa_tree_add_51_79_groupi_n_7035 ,csa_tree_add_51_79_groupi_n_6084 ,csa_tree_add_51_79_groupi_n_6689);
  and csa_tree_add_51_79_groupi_g39092(csa_tree_add_51_79_groupi_n_7034 ,csa_tree_add_51_79_groupi_n_5932 ,csa_tree_add_51_79_groupi_n_6619);
  and csa_tree_add_51_79_groupi_g39093(csa_tree_add_51_79_groupi_n_7033 ,csa_tree_add_51_79_groupi_n_6038 ,csa_tree_add_51_79_groupi_n_6678);
  and csa_tree_add_51_79_groupi_g39094(csa_tree_add_51_79_groupi_n_7032 ,csa_tree_add_51_79_groupi_n_6036 ,csa_tree_add_51_79_groupi_n_6677);
  and csa_tree_add_51_79_groupi_g39095(csa_tree_add_51_79_groupi_n_7031 ,csa_tree_add_51_79_groupi_n_5927 ,csa_tree_add_51_79_groupi_n_6616);
  and csa_tree_add_51_79_groupi_g39096(csa_tree_add_51_79_groupi_n_7030 ,csa_tree_add_51_79_groupi_n_5923 ,csa_tree_add_51_79_groupi_n_6613);
  and csa_tree_add_51_79_groupi_g39097(csa_tree_add_51_79_groupi_n_7029 ,csa_tree_add_51_79_groupi_n_6105 ,csa_tree_add_51_79_groupi_n_6501);
  and csa_tree_add_51_79_groupi_g39098(csa_tree_add_51_79_groupi_n_7028 ,csa_tree_add_51_79_groupi_n_6120 ,csa_tree_add_51_79_groupi_n_6676);
  and csa_tree_add_51_79_groupi_g39099(csa_tree_add_51_79_groupi_n_7027 ,csa_tree_add_51_79_groupi_n_5963 ,csa_tree_add_51_79_groupi_n_6609);
  and csa_tree_add_51_79_groupi_g39100(csa_tree_add_51_79_groupi_n_7026 ,csa_tree_add_51_79_groupi_n_5911 ,csa_tree_add_51_79_groupi_n_6605);
  and csa_tree_add_51_79_groupi_g39101(csa_tree_add_51_79_groupi_n_7025 ,csa_tree_add_51_79_groupi_n_5685 ,csa_tree_add_51_79_groupi_n_6606);
  and csa_tree_add_51_79_groupi_g39102(csa_tree_add_51_79_groupi_n_7023 ,csa_tree_add_51_79_groupi_n_5731 ,csa_tree_add_51_79_groupi_n_6603);
  and csa_tree_add_51_79_groupi_g39103(csa_tree_add_51_79_groupi_n_7022 ,csa_tree_add_51_79_groupi_n_6045 ,csa_tree_add_51_79_groupi_n_6604);
  and csa_tree_add_51_79_groupi_g39104(csa_tree_add_51_79_groupi_n_7021 ,csa_tree_add_51_79_groupi_n_6034 ,csa_tree_add_51_79_groupi_n_6669);
  and csa_tree_add_51_79_groupi_g39105(csa_tree_add_51_79_groupi_n_7020 ,csa_tree_add_51_79_groupi_n_6112 ,csa_tree_add_51_79_groupi_n_6710);
  and csa_tree_add_51_79_groupi_g39106(csa_tree_add_51_79_groupi_n_7019 ,csa_tree_add_51_79_groupi_n_6111 ,csa_tree_add_51_79_groupi_n_6712);
  and csa_tree_add_51_79_groupi_g39107(csa_tree_add_51_79_groupi_n_7018 ,csa_tree_add_51_79_groupi_n_6029 ,csa_tree_add_51_79_groupi_n_6672);
  and csa_tree_add_51_79_groupi_g39108(csa_tree_add_51_79_groupi_n_7017 ,csa_tree_add_51_79_groupi_n_5733 ,csa_tree_add_51_79_groupi_n_6632);
  and csa_tree_add_51_79_groupi_g39109(csa_tree_add_51_79_groupi_n_7016 ,csa_tree_add_51_79_groupi_n_5777 ,csa_tree_add_51_79_groupi_n_6597);
  and csa_tree_add_51_79_groupi_g39110(csa_tree_add_51_79_groupi_n_7015 ,csa_tree_add_51_79_groupi_n_6107 ,csa_tree_add_51_79_groupi_n_6711);
  and csa_tree_add_51_79_groupi_g39111(csa_tree_add_51_79_groupi_n_7014 ,csa_tree_add_51_79_groupi_n_5894 ,csa_tree_add_51_79_groupi_n_6596);
  and csa_tree_add_51_79_groupi_g39112(csa_tree_add_51_79_groupi_n_7013 ,csa_tree_add_51_79_groupi_n_6109 ,csa_tree_add_51_79_groupi_n_6554);
  and csa_tree_add_51_79_groupi_g39113(csa_tree_add_51_79_groupi_n_7012 ,csa_tree_add_51_79_groupi_n_6075 ,csa_tree_add_51_79_groupi_n_6699);
  and csa_tree_add_51_79_groupi_g39114(csa_tree_add_51_79_groupi_n_7010 ,csa_tree_add_51_79_groupi_n_5885 ,csa_tree_add_51_79_groupi_n_6593);
  and csa_tree_add_51_79_groupi_g39115(csa_tree_add_51_79_groupi_n_7008 ,csa_tree_add_51_79_groupi_n_5884 ,csa_tree_add_51_79_groupi_n_6594);
  and csa_tree_add_51_79_groupi_g39116(csa_tree_add_51_79_groupi_n_7006 ,csa_tree_add_51_79_groupi_n_6023 ,csa_tree_add_51_79_groupi_n_6667);
  and csa_tree_add_51_79_groupi_g39117(csa_tree_add_51_79_groupi_n_7005 ,csa_tree_add_51_79_groupi_n_6074 ,csa_tree_add_51_79_groupi_n_6698);
  and csa_tree_add_51_79_groupi_g39118(csa_tree_add_51_79_groupi_n_7004 ,csa_tree_add_51_79_groupi_n_6021 ,csa_tree_add_51_79_groupi_n_6668);
  and csa_tree_add_51_79_groupi_g39119(csa_tree_add_51_79_groupi_n_7003 ,csa_tree_add_51_79_groupi_n_6106 ,csa_tree_add_51_79_groupi_n_6707);
  and csa_tree_add_51_79_groupi_g39120(csa_tree_add_51_79_groupi_n_7001 ,csa_tree_add_51_79_groupi_n_5879 ,csa_tree_add_51_79_groupi_n_6513);
  or csa_tree_add_51_79_groupi_g39121(csa_tree_add_51_79_groupi_n_7000 ,csa_tree_add_51_79_groupi_n_5905 ,csa_tree_add_51_79_groupi_n_6560);
  and csa_tree_add_51_79_groupi_g39122(csa_tree_add_51_79_groupi_n_6999 ,csa_tree_add_51_79_groupi_n_5886 ,csa_tree_add_51_79_groupi_n_6588);
  and csa_tree_add_51_79_groupi_g39123(csa_tree_add_51_79_groupi_n_6998 ,csa_tree_add_51_79_groupi_n_5895 ,csa_tree_add_51_79_groupi_n_6583);
  and csa_tree_add_51_79_groupi_g39124(csa_tree_add_51_79_groupi_n_6997 ,csa_tree_add_51_79_groupi_n_5893 ,csa_tree_add_51_79_groupi_n_6585);
  and csa_tree_add_51_79_groupi_g39125(csa_tree_add_51_79_groupi_n_6995 ,csa_tree_add_51_79_groupi_n_5630 ,csa_tree_add_51_79_groupi_n_6587);
  and csa_tree_add_51_79_groupi_g39126(csa_tree_add_51_79_groupi_n_6994 ,csa_tree_add_51_79_groupi_n_6018 ,csa_tree_add_51_79_groupi_n_6666);
  and csa_tree_add_51_79_groupi_g39127(csa_tree_add_51_79_groupi_n_6993 ,csa_tree_add_51_79_groupi_n_6070 ,csa_tree_add_51_79_groupi_n_6697);
  and csa_tree_add_51_79_groupi_g39128(csa_tree_add_51_79_groupi_n_6992 ,csa_tree_add_51_79_groupi_n_5820 ,csa_tree_add_51_79_groupi_n_6559);
  and csa_tree_add_51_79_groupi_g39129(csa_tree_add_51_79_groupi_n_6991 ,csa_tree_add_51_79_groupi_n_5913 ,csa_tree_add_51_79_groupi_n_6581);
  and csa_tree_add_51_79_groupi_g39130(csa_tree_add_51_79_groupi_n_6990 ,csa_tree_add_51_79_groupi_n_6009 ,csa_tree_add_51_79_groupi_n_6662);
  and csa_tree_add_51_79_groupi_g39131(csa_tree_add_51_79_groupi_n_6989 ,csa_tree_add_51_79_groupi_n_6008 ,csa_tree_add_51_79_groupi_n_6663);
  and csa_tree_add_51_79_groupi_g39132(csa_tree_add_51_79_groupi_n_6988 ,csa_tree_add_51_79_groupi_n_5958 ,csa_tree_add_51_79_groupi_n_6578);
  and csa_tree_add_51_79_groupi_g39133(csa_tree_add_51_79_groupi_n_6986 ,csa_tree_add_51_79_groupi_n_6006 ,csa_tree_add_51_79_groupi_n_6661);
  and csa_tree_add_51_79_groupi_g39134(csa_tree_add_51_79_groupi_n_6985 ,csa_tree_add_51_79_groupi_n_5991 ,csa_tree_add_51_79_groupi_n_6645);
  and csa_tree_add_51_79_groupi_g39135(csa_tree_add_51_79_groupi_n_6983 ,csa_tree_add_51_79_groupi_n_5979 ,csa_tree_add_51_79_groupi_n_6579);
  and csa_tree_add_51_79_groupi_g39136(csa_tree_add_51_79_groupi_n_6982 ,csa_tree_add_51_79_groupi_n_6043 ,csa_tree_add_51_79_groupi_n_6577);
  and csa_tree_add_51_79_groupi_g39137(csa_tree_add_51_79_groupi_n_6981 ,csa_tree_add_51_79_groupi_n_5998 ,csa_tree_add_51_79_groupi_n_6646);
  and csa_tree_add_51_79_groupi_g39138(csa_tree_add_51_79_groupi_n_6979 ,csa_tree_add_51_79_groupi_n_5697 ,csa_tree_add_51_79_groupi_n_6571);
  and csa_tree_add_51_79_groupi_g39139(csa_tree_add_51_79_groupi_n_6978 ,csa_tree_add_51_79_groupi_n_6119 ,csa_tree_add_51_79_groupi_n_6570);
  and csa_tree_add_51_79_groupi_g39140(csa_tree_add_51_79_groupi_n_6977 ,csa_tree_add_51_79_groupi_n_5838 ,csa_tree_add_51_79_groupi_n_6573);
  and csa_tree_add_51_79_groupi_g39141(csa_tree_add_51_79_groupi_n_6976 ,csa_tree_add_51_79_groupi_n_5837 ,csa_tree_add_51_79_groupi_n_6547);
  and csa_tree_add_51_79_groupi_g39142(csa_tree_add_51_79_groupi_n_6975 ,csa_tree_add_51_79_groupi_n_6003 ,csa_tree_add_51_79_groupi_n_6658);
  and csa_tree_add_51_79_groupi_g39143(csa_tree_add_51_79_groupi_n_6974 ,csa_tree_add_51_79_groupi_n_5833 ,csa_tree_add_51_79_groupi_n_6568);
  and csa_tree_add_51_79_groupi_g39144(csa_tree_add_51_79_groupi_n_6973 ,csa_tree_add_51_79_groupi_n_6123 ,csa_tree_add_51_79_groupi_n_6714);
  and csa_tree_add_51_79_groupi_g39145(csa_tree_add_51_79_groupi_n_6972 ,csa_tree_add_51_79_groupi_n_5999 ,csa_tree_add_51_79_groupi_n_6657);
  and csa_tree_add_51_79_groupi_g39146(csa_tree_add_51_79_groupi_n_6971 ,csa_tree_add_51_79_groupi_n_5804 ,csa_tree_add_51_79_groupi_n_6491);
  and csa_tree_add_51_79_groupi_g39147(csa_tree_add_51_79_groupi_n_6970 ,csa_tree_add_51_79_groupi_n_5831 ,csa_tree_add_51_79_groupi_n_6564);
  and csa_tree_add_51_79_groupi_g39148(csa_tree_add_51_79_groupi_n_6969 ,csa_tree_add_51_79_groupi_n_5776 ,csa_tree_add_51_79_groupi_n_6567);
  and csa_tree_add_51_79_groupi_g39149(csa_tree_add_51_79_groupi_n_6968 ,csa_tree_add_51_79_groupi_n_5825 ,csa_tree_add_51_79_groupi_n_6565);
  and csa_tree_add_51_79_groupi_g39150(csa_tree_add_51_79_groupi_n_6967 ,csa_tree_add_51_79_groupi_n_5994 ,csa_tree_add_51_79_groupi_n_6655);
  and csa_tree_add_51_79_groupi_g39151(csa_tree_add_51_79_groupi_n_6966 ,csa_tree_add_51_79_groupi_n_6065 ,csa_tree_add_51_79_groupi_n_6694);
  and csa_tree_add_51_79_groupi_g39152(csa_tree_add_51_79_groupi_n_6965 ,csa_tree_add_51_79_groupi_n_5988 ,csa_tree_add_51_79_groupi_n_6653);
  and csa_tree_add_51_79_groupi_g39153(csa_tree_add_51_79_groupi_n_6964 ,csa_tree_add_51_79_groupi_n_5985 ,csa_tree_add_51_79_groupi_n_6651);
  and csa_tree_add_51_79_groupi_g39154(csa_tree_add_51_79_groupi_n_6963 ,csa_tree_add_51_79_groupi_n_6063 ,csa_tree_add_51_79_groupi_n_6692);
  and csa_tree_add_51_79_groupi_g39155(csa_tree_add_51_79_groupi_n_6962 ,csa_tree_add_51_79_groupi_n_5703 ,csa_tree_add_51_79_groupi_n_6541);
  or csa_tree_add_51_79_groupi_g39156(csa_tree_add_51_79_groupi_n_6961 ,csa_tree_add_51_79_groupi_n_6118 ,csa_tree_add_51_79_groupi_n_6716);
  not csa_tree_add_51_79_groupi_g39158(csa_tree_add_51_79_groupi_n_6924 ,csa_tree_add_51_79_groupi_n_6923);
  not csa_tree_add_51_79_groupi_g39160(csa_tree_add_51_79_groupi_n_6896 ,csa_tree_add_51_79_groupi_n_6897);
  not csa_tree_add_51_79_groupi_g39161(csa_tree_add_51_79_groupi_n_6888 ,csa_tree_add_51_79_groupi_n_6887);
  not csa_tree_add_51_79_groupi_g39162(csa_tree_add_51_79_groupi_n_6884 ,csa_tree_add_51_79_groupi_n_6885);
  not csa_tree_add_51_79_groupi_g39163(csa_tree_add_51_79_groupi_n_6876 ,csa_tree_add_51_79_groupi_n_6877);
  not csa_tree_add_51_79_groupi_g39164(csa_tree_add_51_79_groupi_n_6870 ,csa_tree_add_51_79_groupi_n_6871);
  not csa_tree_add_51_79_groupi_g39165(csa_tree_add_51_79_groupi_n_6868 ,csa_tree_add_51_79_groupi_n_6869);
  not csa_tree_add_51_79_groupi_g39166(csa_tree_add_51_79_groupi_n_6866 ,csa_tree_add_51_79_groupi_n_6867);
  not csa_tree_add_51_79_groupi_g39167(csa_tree_add_51_79_groupi_n_6861 ,csa_tree_add_51_79_groupi_n_6860);
  not csa_tree_add_51_79_groupi_g39168(csa_tree_add_51_79_groupi_n_6854 ,csa_tree_add_51_79_groupi_n_6855);
  not csa_tree_add_51_79_groupi_g39169(csa_tree_add_51_79_groupi_n_6853 ,csa_tree_add_51_79_groupi_n_6852);
  not csa_tree_add_51_79_groupi_g39170(csa_tree_add_51_79_groupi_n_6849 ,csa_tree_add_51_79_groupi_n_6850);
  not csa_tree_add_51_79_groupi_g39171(csa_tree_add_51_79_groupi_n_6848 ,csa_tree_add_51_79_groupi_n_23);
  not csa_tree_add_51_79_groupi_g39172(csa_tree_add_51_79_groupi_n_6847 ,csa_tree_add_51_79_groupi_n_22);
  not csa_tree_add_51_79_groupi_g39173(csa_tree_add_51_79_groupi_n_6846 ,csa_tree_add_51_79_groupi_n_21);
  not csa_tree_add_51_79_groupi_g39174(csa_tree_add_51_79_groupi_n_6845 ,csa_tree_add_51_79_groupi_n_20);
  not csa_tree_add_51_79_groupi_g39175(csa_tree_add_51_79_groupi_n_6844 ,csa_tree_add_51_79_groupi_n_13);
  not csa_tree_add_51_79_groupi_g39176(csa_tree_add_51_79_groupi_n_6843 ,csa_tree_add_51_79_groupi_n_12);
  not csa_tree_add_51_79_groupi_g39177(csa_tree_add_51_79_groupi_n_6841 ,csa_tree_add_51_79_groupi_n_18);
  not csa_tree_add_51_79_groupi_g39178(csa_tree_add_51_79_groupi_n_6839 ,csa_tree_add_51_79_groupi_n_15);
  not csa_tree_add_51_79_groupi_g39179(csa_tree_add_51_79_groupi_n_6838 ,csa_tree_add_51_79_groupi_n_16);
  not csa_tree_add_51_79_groupi_g39180(csa_tree_add_51_79_groupi_n_6837 ,csa_tree_add_51_79_groupi_n_17);
  not csa_tree_add_51_79_groupi_g39181(csa_tree_add_51_79_groupi_n_6836 ,csa_tree_add_51_79_groupi_n_19);
  not csa_tree_add_51_79_groupi_g39182(csa_tree_add_51_79_groupi_n_6835 ,csa_tree_add_51_79_groupi_n_14);
  not csa_tree_add_51_79_groupi_g39183(csa_tree_add_51_79_groupi_n_6834 ,csa_tree_add_51_79_groupi_n_6833);
  not csa_tree_add_51_79_groupi_g39184(csa_tree_add_51_79_groupi_n_6822 ,csa_tree_add_51_79_groupi_n_6823);
  or csa_tree_add_51_79_groupi_g39185(csa_tree_add_51_79_groupi_n_6815 ,csa_tree_add_51_79_groupi_n_6446 ,csa_tree_add_51_79_groupi_n_6447);
  and csa_tree_add_51_79_groupi_g39186(csa_tree_add_51_79_groupi_n_6814 ,csa_tree_add_51_79_groupi_n_6433 ,csa_tree_add_51_79_groupi_n_6434);
  or csa_tree_add_51_79_groupi_g39187(csa_tree_add_51_79_groupi_n_6813 ,csa_tree_add_51_79_groupi_n_6152 ,csa_tree_add_51_79_groupi_n_6539);
  or csa_tree_add_51_79_groupi_g39188(csa_tree_add_51_79_groupi_n_6812 ,csa_tree_add_51_79_groupi_n_4803 ,csa_tree_add_51_79_groupi_n_6421);
  nor csa_tree_add_51_79_groupi_g39189(csa_tree_add_51_79_groupi_n_6811 ,csa_tree_add_51_79_groupi_n_6395 ,csa_tree_add_51_79_groupi_n_6397);
  nor csa_tree_add_51_79_groupi_g39190(csa_tree_add_51_79_groupi_n_6810 ,csa_tree_add_51_79_groupi_n_6748 ,csa_tree_add_51_79_groupi_n_6750);
  or csa_tree_add_51_79_groupi_g39191(csa_tree_add_51_79_groupi_n_6809 ,csa_tree_add_51_79_groupi_n_6747 ,csa_tree_add_51_79_groupi_n_6749);
  or csa_tree_add_51_79_groupi_g39192(csa_tree_add_51_79_groupi_n_6808 ,csa_tree_add_51_79_groupi_n_6394 ,csa_tree_add_51_79_groupi_n_6396);
  nor csa_tree_add_51_79_groupi_g39193(csa_tree_add_51_79_groupi_n_6807 ,csa_tree_add_51_79_groupi_n_6726 ,csa_tree_add_51_79_groupi_n_6724);
  or csa_tree_add_51_79_groupi_g39194(csa_tree_add_51_79_groupi_n_6806 ,csa_tree_add_51_79_groupi_n_6725 ,csa_tree_add_51_79_groupi_n_6723);
  nor csa_tree_add_51_79_groupi_g39195(csa_tree_add_51_79_groupi_n_6805 ,csa_tree_add_51_79_groupi_n_6732 ,csa_tree_add_51_79_groupi_n_6730);
  or csa_tree_add_51_79_groupi_g39196(csa_tree_add_51_79_groupi_n_6804 ,csa_tree_add_51_79_groupi_n_6731 ,csa_tree_add_51_79_groupi_n_6729);
  and csa_tree_add_51_79_groupi_g39197(csa_tree_add_51_79_groupi_n_6803 ,csa_tree_add_51_79_groupi_n_6738 ,csa_tree_add_51_79_groupi_n_6737);
  or csa_tree_add_51_79_groupi_g39198(csa_tree_add_51_79_groupi_n_6802 ,csa_tree_add_51_79_groupi_n_6738 ,csa_tree_add_51_79_groupi_n_6737);
  or csa_tree_add_51_79_groupi_g39199(csa_tree_add_51_79_groupi_n_6801 ,csa_tree_add_51_79_groupi_n_6400 ,csa_tree_add_51_79_groupi_n_6441);
  and csa_tree_add_51_79_groupi_g39200(csa_tree_add_51_79_groupi_n_6800 ,csa_tree_add_51_79_groupi_n_6733 ,csa_tree_add_51_79_groupi_n_6448);
  or csa_tree_add_51_79_groupi_g39201(csa_tree_add_51_79_groupi_n_6799 ,csa_tree_add_51_79_groupi_n_6733 ,csa_tree_add_51_79_groupi_n_6448);
  and csa_tree_add_51_79_groupi_g39202(csa_tree_add_51_79_groupi_n_6798 ,csa_tree_add_51_79_groupi_n_6400 ,csa_tree_add_51_79_groupi_n_6441);
  and csa_tree_add_51_79_groupi_g39203(csa_tree_add_51_79_groupi_n_6797 ,csa_tree_add_51_79_groupi_n_6727 ,csa_tree_add_51_79_groupi_n_6440);
  and csa_tree_add_51_79_groupi_g39204(csa_tree_add_51_79_groupi_n_6796 ,csa_tree_add_51_79_groupi_n_6753 ,csa_tree_add_51_79_groupi_n_6449);
  or csa_tree_add_51_79_groupi_g39205(csa_tree_add_51_79_groupi_n_6795 ,csa_tree_add_51_79_groupi_n_4821 ,csa_tree_add_51_79_groupi_n_6450);
  or csa_tree_add_51_79_groupi_g39206(csa_tree_add_51_79_groupi_n_6794 ,csa_tree_add_51_79_groupi_n_6727 ,csa_tree_add_51_79_groupi_n_6440);
  and csa_tree_add_51_79_groupi_g39207(csa_tree_add_51_79_groupi_n_6793 ,csa_tree_add_51_79_groupi_n_6734 ,csa_tree_add_51_79_groupi_n_6435);
  and csa_tree_add_51_79_groupi_g39208(csa_tree_add_51_79_groupi_n_6792 ,csa_tree_add_51_79_groupi_n_4821 ,csa_tree_add_51_79_groupi_n_6450);
  or csa_tree_add_51_79_groupi_g39209(csa_tree_add_51_79_groupi_n_6791 ,csa_tree_add_51_79_groupi_n_6734 ,csa_tree_add_51_79_groupi_n_6435);
  and csa_tree_add_51_79_groupi_g39210(csa_tree_add_51_79_groupi_n_6790 ,csa_tree_add_51_79_groupi_n_6156 ,csa_tree_add_51_79_groupi_n_6505);
  or csa_tree_add_51_79_groupi_g39211(csa_tree_add_51_79_groupi_n_6789 ,csa_tree_add_51_79_groupi_n_6432 ,csa_tree_add_51_79_groupi_n_6431);
  or csa_tree_add_51_79_groupi_g39212(csa_tree_add_51_79_groupi_n_6788 ,csa_tree_add_51_79_groupi_n_5652 ,csa_tree_add_51_79_groupi_n_24);
  nor csa_tree_add_51_79_groupi_g39213(csa_tree_add_51_79_groupi_n_6787 ,csa_tree_add_51_79_groupi_n_6757 ,csa_tree_add_51_79_groupi_n_6752);
  or csa_tree_add_51_79_groupi_g39214(csa_tree_add_51_79_groupi_n_6786 ,csa_tree_add_51_79_groupi_n_5863 ,csa_tree_add_51_79_groupi_n_6481);
  or csa_tree_add_51_79_groupi_g39215(csa_tree_add_51_79_groupi_n_6785 ,csa_tree_add_51_79_groupi_n_5864 ,csa_tree_add_51_79_groupi_n_6506);
  and csa_tree_add_51_79_groupi_g39216(csa_tree_add_51_79_groupi_n_6784 ,csa_tree_add_51_79_groupi_n_6410 ,csa_tree_add_51_79_groupi_n_6416);
  or csa_tree_add_51_79_groupi_g39217(csa_tree_add_51_79_groupi_n_6783 ,csa_tree_add_51_79_groupi_n_5866 ,csa_tree_add_51_79_groupi_n_6679);
  or csa_tree_add_51_79_groupi_g39218(csa_tree_add_51_79_groupi_n_6782 ,csa_tree_add_51_79_groupi_n_6720 ,csa_tree_add_51_79_groupi_n_5843);
  or csa_tree_add_51_79_groupi_g39219(csa_tree_add_51_79_groupi_n_6781 ,csa_tree_add_51_79_groupi_n_6410 ,csa_tree_add_51_79_groupi_n_6416);
  and csa_tree_add_51_79_groupi_g39220(csa_tree_add_51_79_groupi_n_6780 ,csa_tree_add_51_79_groupi_n_6432 ,csa_tree_add_51_79_groupi_n_6431);
  nor csa_tree_add_51_79_groupi_g39221(csa_tree_add_51_79_groupi_n_6779 ,csa_tree_add_51_79_groupi_n_6719 ,csa_tree_add_51_79_groupi_n_5844);
  or csa_tree_add_51_79_groupi_g39222(csa_tree_add_51_79_groupi_n_6778 ,csa_tree_add_51_79_groupi_n_6104 ,csa_tree_add_51_79_groupi_n_6455);
  xnor csa_tree_add_51_79_groupi_g39223(csa_tree_add_51_79_groupi_n_6777 ,csa_tree_add_51_79_groupi_n_5849 ,csa_tree_add_51_79_groupi_n_5850);
  xnor csa_tree_add_51_79_groupi_g39224(csa_tree_add_51_79_groupi_n_6776 ,csa_tree_add_51_79_groupi_n_6139 ,csa_tree_add_51_79_groupi_n_5301);
  xnor csa_tree_add_51_79_groupi_g39225(csa_tree_add_51_79_groupi_n_6775 ,csa_tree_add_51_79_groupi_n_6145 ,csa_tree_add_51_79_groupi_n_6146);
  xnor csa_tree_add_51_79_groupi_g39226(csa_tree_add_51_79_groupi_n_6774 ,csa_tree_add_51_79_groupi_n_5842 ,csa_tree_add_51_79_groupi_n_5859);
  xnor csa_tree_add_51_79_groupi_g39227(csa_tree_add_51_79_groupi_n_6773 ,csa_tree_add_51_79_groupi_n_4804 ,csa_tree_add_51_79_groupi_n_5865);
  xnor csa_tree_add_51_79_groupi_g39228(csa_tree_add_51_79_groupi_n_6772 ,csa_tree_add_51_79_groupi_n_5856 ,csa_tree_add_51_79_groupi_n_5858);
  xor csa_tree_add_51_79_groupi_g39229(csa_tree_add_51_79_groupi_n_6771 ,csa_tree_add_51_79_groupi_n_5279 ,csa_tree_add_51_79_groupi_n_6150);
  xnor csa_tree_add_51_79_groupi_g39230(csa_tree_add_51_79_groupi_n_6770 ,csa_tree_add_51_79_groupi_n_5335 ,csa_tree_add_51_79_groupi_n_6153);
  xnor csa_tree_add_51_79_groupi_g39231(csa_tree_add_51_79_groupi_n_6769 ,csa_tree_add_51_79_groupi_n_5866 ,csa_tree_add_51_79_groupi_n_5854);
  xnor csa_tree_add_51_79_groupi_g39232(csa_tree_add_51_79_groupi_n_6768 ,csa_tree_add_51_79_groupi_n_5401 ,csa_tree_add_51_79_groupi_n_6143);
  xnor csa_tree_add_51_79_groupi_g39233(csa_tree_add_51_79_groupi_n_6767 ,csa_tree_add_51_79_groupi_n_6147 ,csa_tree_add_51_79_groupi_n_6132);
  xnor csa_tree_add_51_79_groupi_g39234(csa_tree_add_51_79_groupi_n_6766 ,csa_tree_add_51_79_groupi_n_6152 ,csa_tree_add_51_79_groupi_n_6141);
  xnor csa_tree_add_51_79_groupi_g39235(csa_tree_add_51_79_groupi_n_6765 ,csa_tree_add_51_79_groupi_n_6140 ,csa_tree_add_51_79_groupi_n_5860);
  xnor csa_tree_add_51_79_groupi_g39236(csa_tree_add_51_79_groupi_n_6764 ,csa_tree_add_51_79_groupi_n_5845 ,csa_tree_add_51_79_groupi_n_5864);
  xnor csa_tree_add_51_79_groupi_g39237(csa_tree_add_51_79_groupi_n_6763 ,csa_tree_add_51_79_groupi_n_6138 ,csa_tree_add_51_79_groupi_n_6155);
  and csa_tree_add_51_79_groupi_g39238(csa_tree_add_51_79_groupi_n_6939 ,csa_tree_add_51_79_groupi_n_5609 ,csa_tree_add_51_79_groupi_n_6522);
  and csa_tree_add_51_79_groupi_g39239(csa_tree_add_51_79_groupi_n_6938 ,csa_tree_add_51_79_groupi_n_5702 ,csa_tree_add_51_79_groupi_n_6500);
  and csa_tree_add_51_79_groupi_g39240(csa_tree_add_51_79_groupi_n_6937 ,csa_tree_add_51_79_groupi_n_5694 ,csa_tree_add_51_79_groupi_n_6496);
  and csa_tree_add_51_79_groupi_g39241(csa_tree_add_51_79_groupi_n_6936 ,csa_tree_add_51_79_groupi_n_5692 ,csa_tree_add_51_79_groupi_n_6494);
  and csa_tree_add_51_79_groupi_g39242(csa_tree_add_51_79_groupi_n_6935 ,csa_tree_add_51_79_groupi_n_5689 ,csa_tree_add_51_79_groupi_n_6480);
  and csa_tree_add_51_79_groupi_g39243(csa_tree_add_51_79_groupi_n_6934 ,csa_tree_add_51_79_groupi_n_5751 ,csa_tree_add_51_79_groupi_n_6674);
  and csa_tree_add_51_79_groupi_g39244(csa_tree_add_51_79_groupi_n_6933 ,csa_tree_add_51_79_groupi_n_5674 ,csa_tree_add_51_79_groupi_n_6488);
  and csa_tree_add_51_79_groupi_g39245(csa_tree_add_51_79_groupi_n_6932 ,csa_tree_add_51_79_groupi_n_5669 ,csa_tree_add_51_79_groupi_n_6484);
  and csa_tree_add_51_79_groupi_g39246(csa_tree_add_51_79_groupi_n_6931 ,csa_tree_add_51_79_groupi_n_5664 ,csa_tree_add_51_79_groupi_n_6483);
  or csa_tree_add_51_79_groupi_g39247(csa_tree_add_51_79_groupi_n_6930 ,csa_tree_add_51_79_groupi_n_5656 ,csa_tree_add_51_79_groupi_n_6476);
  and csa_tree_add_51_79_groupi_g39248(csa_tree_add_51_79_groupi_n_6929 ,csa_tree_add_51_79_groupi_n_5726 ,csa_tree_add_51_79_groupi_n_6717);
  and csa_tree_add_51_79_groupi_g39249(csa_tree_add_51_79_groupi_n_6928 ,csa_tree_add_51_79_groupi_n_5647 ,csa_tree_add_51_79_groupi_n_6474);
  and csa_tree_add_51_79_groupi_g39250(csa_tree_add_51_79_groupi_n_6927 ,csa_tree_add_51_79_groupi_n_5637 ,csa_tree_add_51_79_groupi_n_6470);
  and csa_tree_add_51_79_groupi_g39251(csa_tree_add_51_79_groupi_n_6926 ,csa_tree_add_51_79_groupi_n_5636 ,csa_tree_add_51_79_groupi_n_6469);
  and csa_tree_add_51_79_groupi_g39252(csa_tree_add_51_79_groupi_n_6925 ,csa_tree_add_51_79_groupi_n_5625 ,csa_tree_add_51_79_groupi_n_6464);
  or csa_tree_add_51_79_groupi_g39253(csa_tree_add_51_79_groupi_n_6923 ,csa_tree_add_51_79_groupi_n_5622 ,csa_tree_add_51_79_groupi_n_6462);
  and csa_tree_add_51_79_groupi_g39254(csa_tree_add_51_79_groupi_n_6922 ,csa_tree_add_51_79_groupi_n_5620 ,csa_tree_add_51_79_groupi_n_6465);
  and csa_tree_add_51_79_groupi_g39255(csa_tree_add_51_79_groupi_n_6921 ,csa_tree_add_51_79_groupi_n_5915 ,csa_tree_add_51_79_groupi_n_6715);
  and csa_tree_add_51_79_groupi_g39256(csa_tree_add_51_79_groupi_n_6920 ,csa_tree_add_51_79_groupi_n_5613 ,csa_tree_add_51_79_groupi_n_6574);
  and csa_tree_add_51_79_groupi_g39257(csa_tree_add_51_79_groupi_n_6919 ,csa_tree_add_51_79_groupi_n_5599 ,csa_tree_add_51_79_groupi_n_6628);
  and csa_tree_add_51_79_groupi_g39258(csa_tree_add_51_79_groupi_n_6918 ,csa_tree_add_51_79_groupi_n_5764 ,csa_tree_add_51_79_groupi_n_6537);
  and csa_tree_add_51_79_groupi_g39259(csa_tree_add_51_79_groupi_n_6917 ,csa_tree_add_51_79_groupi_n_5607 ,csa_tree_add_51_79_groupi_n_6527);
  and csa_tree_add_51_79_groupi_g39260(csa_tree_add_51_79_groupi_n_6916 ,csa_tree_add_51_79_groupi_n_5601 ,csa_tree_add_51_79_groupi_n_6607);
  and csa_tree_add_51_79_groupi_g39261(csa_tree_add_51_79_groupi_n_6915 ,csa_tree_add_51_79_groupi_n_5922 ,csa_tree_add_51_79_groupi_n_6550);
  and csa_tree_add_51_79_groupi_g39262(csa_tree_add_51_79_groupi_n_6914 ,csa_tree_add_51_79_groupi_n_5740 ,csa_tree_add_51_79_groupi_n_6515);
  and csa_tree_add_51_79_groupi_g39263(csa_tree_add_51_79_groupi_n_6913 ,csa_tree_add_51_79_groupi_n_5741 ,csa_tree_add_51_79_groupi_n_6518);
  and csa_tree_add_51_79_groupi_g39264(csa_tree_add_51_79_groupi_n_6912 ,csa_tree_add_51_79_groupi_n_5743 ,csa_tree_add_51_79_groupi_n_6517);
  and csa_tree_add_51_79_groupi_g39265(csa_tree_add_51_79_groupi_n_6911 ,csa_tree_add_51_79_groupi_n_5964 ,csa_tree_add_51_79_groupi_n_6562);
  and csa_tree_add_51_79_groupi_g39266(csa_tree_add_51_79_groupi_n_6910 ,csa_tree_add_51_79_groupi_n_5704 ,csa_tree_add_51_79_groupi_n_6533);
  and csa_tree_add_51_79_groupi_g39267(csa_tree_add_51_79_groupi_n_6909 ,csa_tree_add_51_79_groupi_n_5827 ,csa_tree_add_51_79_groupi_n_6566);
  and csa_tree_add_51_79_groupi_g39268(csa_tree_add_51_79_groupi_n_6908 ,csa_tree_add_51_79_groupi_n_6121 ,csa_tree_add_51_79_groupi_n_6528);
  and csa_tree_add_51_79_groupi_g39269(csa_tree_add_51_79_groupi_n_6907 ,csa_tree_add_51_79_groupi_n_5775 ,csa_tree_add_51_79_groupi_n_6553);
  and csa_tree_add_51_79_groupi_g39270(csa_tree_add_51_79_groupi_n_6906 ,csa_tree_add_51_79_groupi_n_5779 ,csa_tree_add_51_79_groupi_n_6503);
  and csa_tree_add_51_79_groupi_g39271(csa_tree_add_51_79_groupi_n_6905 ,csa_tree_add_51_79_groupi_n_6122 ,csa_tree_add_51_79_groupi_n_6612);
  and csa_tree_add_51_79_groupi_g39272(csa_tree_add_51_79_groupi_n_6904 ,csa_tree_add_51_79_groupi_n_5786 ,csa_tree_add_51_79_groupi_n_6543);
  and csa_tree_add_51_79_groupi_g39273(csa_tree_add_51_79_groupi_n_6903 ,csa_tree_add_51_79_groupi_n_5785 ,csa_tree_add_51_79_groupi_n_6639);
  and csa_tree_add_51_79_groupi_g39274(csa_tree_add_51_79_groupi_n_6902 ,csa_tree_add_51_79_groupi_n_5780 ,csa_tree_add_51_79_groupi_n_6544);
  and csa_tree_add_51_79_groupi_g39275(csa_tree_add_51_79_groupi_n_6901 ,csa_tree_add_51_79_groupi_n_5881 ,csa_tree_add_51_79_groupi_n_6502);
  and csa_tree_add_51_79_groupi_g39276(csa_tree_add_51_79_groupi_n_6900 ,csa_tree_add_51_79_groupi_n_5797 ,csa_tree_add_51_79_groupi_n_6549);
  and csa_tree_add_51_79_groupi_g39277(csa_tree_add_51_79_groupi_n_6899 ,csa_tree_add_51_79_groupi_n_6125 ,csa_tree_add_51_79_groupi_n_6713);
  and csa_tree_add_51_79_groupi_g39278(csa_tree_add_51_79_groupi_n_6898 ,csa_tree_add_51_79_groupi_n_5680 ,csa_tree_add_51_79_groupi_n_6487);
  or csa_tree_add_51_79_groupi_g39279(csa_tree_add_51_79_groupi_n_6897 ,csa_tree_add_51_79_groupi_n_5798 ,csa_tree_add_51_79_groupi_n_6461);
  and csa_tree_add_51_79_groupi_g39280(csa_tree_add_51_79_groupi_n_6895 ,csa_tree_add_51_79_groupi_n_5678 ,csa_tree_add_51_79_groupi_n_6489);
  and csa_tree_add_51_79_groupi_g39281(csa_tree_add_51_79_groupi_n_6894 ,csa_tree_add_51_79_groupi_n_5698 ,csa_tree_add_51_79_groupi_n_6499);
  and csa_tree_add_51_79_groupi_g39282(csa_tree_add_51_79_groupi_n_6893 ,csa_tree_add_51_79_groupi_n_5696 ,csa_tree_add_51_79_groupi_n_6497);
  and csa_tree_add_51_79_groupi_g39283(csa_tree_add_51_79_groupi_n_6892 ,csa_tree_add_51_79_groupi_n_5670 ,csa_tree_add_51_79_groupi_n_6486);
  and csa_tree_add_51_79_groupi_g39284(csa_tree_add_51_79_groupi_n_6891 ,csa_tree_add_51_79_groupi_n_5744 ,csa_tree_add_51_79_groupi_n_6507);
  and csa_tree_add_51_79_groupi_g39285(csa_tree_add_51_79_groupi_n_6890 ,csa_tree_add_51_79_groupi_n_5732 ,csa_tree_add_51_79_groupi_n_6552);
  and csa_tree_add_51_79_groupi_g39286(csa_tree_add_51_79_groupi_n_6889 ,csa_tree_add_51_79_groupi_n_5666 ,csa_tree_add_51_79_groupi_n_6485);
  or csa_tree_add_51_79_groupi_g39287(csa_tree_add_51_79_groupi_n_6887 ,csa_tree_add_51_79_groupi_n_5668 ,csa_tree_add_51_79_groupi_n_6479);
  and csa_tree_add_51_79_groupi_g39288(csa_tree_add_51_79_groupi_n_6886 ,csa_tree_add_51_79_groupi_n_5606 ,csa_tree_add_51_79_groupi_n_6525);
  and csa_tree_add_51_79_groupi_g39289(csa_tree_add_51_79_groupi_n_6885 ,csa_tree_add_51_79_groupi_n_5713 ,csa_tree_add_51_79_groupi_n_6614);
  and csa_tree_add_51_79_groupi_g39290(csa_tree_add_51_79_groupi_n_6883 ,csa_tree_add_51_79_groupi_n_5603 ,csa_tree_add_51_79_groupi_n_6580);
  and csa_tree_add_51_79_groupi_g39291(csa_tree_add_51_79_groupi_n_6882 ,csa_tree_add_51_79_groupi_n_5801 ,csa_tree_add_51_79_groupi_n_6524);
  and csa_tree_add_51_79_groupi_g39292(csa_tree_add_51_79_groupi_n_6881 ,csa_tree_add_51_79_groupi_n_5605 ,csa_tree_add_51_79_groupi_n_6534);
  and csa_tree_add_51_79_groupi_g39293(csa_tree_add_51_79_groupi_n_6880 ,csa_tree_add_51_79_groupi_n_5723 ,csa_tree_add_51_79_groupi_n_6542);
  and csa_tree_add_51_79_groupi_g39294(csa_tree_add_51_79_groupi_n_6879 ,csa_tree_add_51_79_groupi_n_5738 ,csa_tree_add_51_79_groupi_n_6516);
  and csa_tree_add_51_79_groupi_g39295(csa_tree_add_51_79_groupi_n_6878 ,csa_tree_add_51_79_groupi_n_5611 ,csa_tree_add_51_79_groupi_n_6514);
  or csa_tree_add_51_79_groupi_g39296(csa_tree_add_51_79_groupi_n_6877 ,csa_tree_add_51_79_groupi_n_5717 ,csa_tree_add_51_79_groupi_n_6504);
  and csa_tree_add_51_79_groupi_g39297(csa_tree_add_51_79_groupi_n_6875 ,csa_tree_add_51_79_groupi_n_5653 ,csa_tree_add_51_79_groupi_n_6477);
  and csa_tree_add_51_79_groupi_g39298(csa_tree_add_51_79_groupi_n_6874 ,csa_tree_add_51_79_groupi_n_5649 ,csa_tree_add_51_79_groupi_n_6475);
  and csa_tree_add_51_79_groupi_g39299(csa_tree_add_51_79_groupi_n_6873 ,csa_tree_add_51_79_groupi_n_5746 ,csa_tree_add_51_79_groupi_n_6520);
  and csa_tree_add_51_79_groupi_g39300(csa_tree_add_51_79_groupi_n_6872 ,csa_tree_add_51_79_groupi_n_5684 ,csa_tree_add_51_79_groupi_n_6492);
  or csa_tree_add_51_79_groupi_g39301(csa_tree_add_51_79_groupi_n_6871 ,csa_tree_add_51_79_groupi_n_5914 ,csa_tree_add_51_79_groupi_n_6673);
  or csa_tree_add_51_79_groupi_g39302(csa_tree_add_51_79_groupi_n_6869 ,csa_tree_add_51_79_groupi_n_5872 ,csa_tree_add_51_79_groupi_n_6652);
  or csa_tree_add_51_79_groupi_g39303(csa_tree_add_51_79_groupi_n_6867 ,csa_tree_add_51_79_groupi_n_5948 ,csa_tree_add_51_79_groupi_n_6693);
  and csa_tree_add_51_79_groupi_g39304(csa_tree_add_51_79_groupi_n_6865 ,csa_tree_add_51_79_groupi_n_5722 ,csa_tree_add_51_79_groupi_n_6546);
  and csa_tree_add_51_79_groupi_g39305(csa_tree_add_51_79_groupi_n_6864 ,csa_tree_add_51_79_groupi_n_6001 ,csa_tree_add_51_79_groupi_n_6526);
  and csa_tree_add_51_79_groupi_g39306(csa_tree_add_51_79_groupi_n_6863 ,csa_tree_add_51_79_groupi_n_5754 ,csa_tree_add_51_79_groupi_n_6548);
  and csa_tree_add_51_79_groupi_g39307(csa_tree_add_51_79_groupi_n_6862 ,csa_tree_add_51_79_groupi_n_5729 ,csa_tree_add_51_79_groupi_n_6523);
  and csa_tree_add_51_79_groupi_g39308(csa_tree_add_51_79_groupi_n_6860 ,csa_tree_add_51_79_groupi_n_5646 ,csa_tree_add_51_79_groupi_n_6472);
  and csa_tree_add_51_79_groupi_g39309(csa_tree_add_51_79_groupi_n_6859 ,csa_tree_add_51_79_groupi_n_5644 ,csa_tree_add_51_79_groupi_n_6473);
  and csa_tree_add_51_79_groupi_g39310(csa_tree_add_51_79_groupi_n_6858 ,csa_tree_add_51_79_groupi_n_6101 ,csa_tree_add_51_79_groupi_n_6529);
  and csa_tree_add_51_79_groupi_g39311(csa_tree_add_51_79_groupi_n_6857 ,csa_tree_add_51_79_groupi_n_5760 ,csa_tree_add_51_79_groupi_n_6531);
  and csa_tree_add_51_79_groupi_g39312(csa_tree_add_51_79_groupi_n_6856 ,csa_tree_add_51_79_groupi_n_5761 ,csa_tree_add_51_79_groupi_n_6532);
  and csa_tree_add_51_79_groupi_g39313(csa_tree_add_51_79_groupi_n_6855 ,csa_tree_add_51_79_groupi_n_5753 ,csa_tree_add_51_79_groupi_n_6638);
  and csa_tree_add_51_79_groupi_g39314(csa_tree_add_51_79_groupi_n_6852 ,csa_tree_add_51_79_groupi_n_5767 ,csa_tree_add_51_79_groupi_n_6530);
  and csa_tree_add_51_79_groupi_g39315(csa_tree_add_51_79_groupi_n_6851 ,csa_tree_add_51_79_groupi_n_5768 ,csa_tree_add_51_79_groupi_n_6641);
  xnor csa_tree_add_51_79_groupi_g39316(csa_tree_add_51_79_groupi_n_6850 ,csa_tree_add_51_79_groupi_n_4284 ,csa_tree_add_51_79_groupi_n_5861);
  and csa_tree_add_51_79_groupi_g39323(csa_tree_add_51_79_groupi_n_6842 ,csa_tree_add_51_79_groupi_n_5772 ,csa_tree_add_51_79_groupi_n_6536);
  and csa_tree_add_51_79_groupi_g39325(csa_tree_add_51_79_groupi_n_6840 ,csa_tree_add_51_79_groupi_n_5747 ,csa_tree_add_51_79_groupi_n_6535);
  or csa_tree_add_51_79_groupi_g39331(csa_tree_add_51_79_groupi_n_6833 ,csa_tree_add_51_79_groupi_n_5641 ,csa_tree_add_51_79_groupi_n_6463);
  xnor csa_tree_add_51_79_groupi_g39332(csa_tree_add_51_79_groupi_n_6832 ,csa_tree_add_51_79_groupi_n_4286 ,csa_tree_add_51_79_groupi_n_5589);
  xnor csa_tree_add_51_79_groupi_g39333(csa_tree_add_51_79_groupi_n_6831 ,csa_tree_add_51_79_groupi_n_4300 ,csa_tree_add_51_79_groupi_n_5590);
  xnor csa_tree_add_51_79_groupi_g39334(csa_tree_add_51_79_groupi_n_6830 ,csa_tree_add_51_79_groupi_n_4292 ,csa_tree_add_51_79_groupi_n_5591);
  xnor csa_tree_add_51_79_groupi_g39335(csa_tree_add_51_79_groupi_n_6829 ,csa_tree_add_51_79_groupi_n_4287 ,csa_tree_add_51_79_groupi_n_5592);
  and csa_tree_add_51_79_groupi_g39336(csa_tree_add_51_79_groupi_n_6828 ,csa_tree_add_51_79_groupi_n_5642 ,csa_tree_add_51_79_groupi_n_6471);
  and csa_tree_add_51_79_groupi_g39337(csa_tree_add_51_79_groupi_n_6827 ,csa_tree_add_51_79_groupi_n_5699 ,csa_tree_add_51_79_groupi_n_6498);
  and csa_tree_add_51_79_groupi_g39338(csa_tree_add_51_79_groupi_n_6826 ,csa_tree_add_51_79_groupi_n_5918 ,csa_tree_add_51_79_groupi_n_6637);
  and csa_tree_add_51_79_groupi_g39339(csa_tree_add_51_79_groupi_n_6825 ,csa_tree_add_51_79_groupi_n_5794 ,csa_tree_add_51_79_groupi_n_6511);
  and csa_tree_add_51_79_groupi_g39340(csa_tree_add_51_79_groupi_n_6824 ,csa_tree_add_51_79_groupi_n_5682 ,csa_tree_add_51_79_groupi_n_6490);
  or csa_tree_add_51_79_groupi_g39341(csa_tree_add_51_79_groupi_n_6823 ,csa_tree_add_51_79_groupi_n_5634 ,csa_tree_add_51_79_groupi_n_6468);
  and csa_tree_add_51_79_groupi_g39342(csa_tree_add_51_79_groupi_n_6821 ,csa_tree_add_51_79_groupi_n_5790 ,csa_tree_add_51_79_groupi_n_6545);
  or csa_tree_add_51_79_groupi_g39343(csa_tree_add_51_79_groupi_n_6820 ,csa_tree_add_51_79_groupi_n_5612 ,csa_tree_add_51_79_groupi_n_6687);
  and csa_tree_add_51_79_groupi_g39344(csa_tree_add_51_79_groupi_n_6819 ,csa_tree_add_51_79_groupi_n_5629 ,csa_tree_add_51_79_groupi_n_6467);
  xnor csa_tree_add_51_79_groupi_g39345(csa_tree_add_51_79_groupi_n_6818 ,csa_tree_add_51_79_groupi_n_4285 ,csa_tree_add_51_79_groupi_n_5593);
  and csa_tree_add_51_79_groupi_g39346(csa_tree_add_51_79_groupi_n_6817 ,csa_tree_add_51_79_groupi_n_5806 ,csa_tree_add_51_79_groupi_n_6551);
  and csa_tree_add_51_79_groupi_g39347(csa_tree_add_51_79_groupi_n_6816 ,csa_tree_add_51_79_groupi_n_5627 ,csa_tree_add_51_79_groupi_n_6466);
  not csa_tree_add_51_79_groupi_g39349(csa_tree_add_51_79_groupi_n_6757 ,csa_tree_add_51_79_groupi_n_6756);
  not csa_tree_add_51_79_groupi_g39350(csa_tree_add_51_79_groupi_n_6754 ,csa_tree_add_51_79_groupi_n_6755);
  not csa_tree_add_51_79_groupi_g39351(csa_tree_add_51_79_groupi_n_6751 ,csa_tree_add_51_79_groupi_n_6752);
  not csa_tree_add_51_79_groupi_g39352(csa_tree_add_51_79_groupi_n_6750 ,csa_tree_add_51_79_groupi_n_6749);
  not csa_tree_add_51_79_groupi_g39353(csa_tree_add_51_79_groupi_n_6748 ,csa_tree_add_51_79_groupi_n_6747);
  not csa_tree_add_51_79_groupi_g39354(csa_tree_add_51_79_groupi_n_6744 ,csa_tree_add_51_79_groupi_n_6745);
  not csa_tree_add_51_79_groupi_g39355(csa_tree_add_51_79_groupi_n_6742 ,csa_tree_add_51_79_groupi_n_6741);
  not csa_tree_add_51_79_groupi_g39356(csa_tree_add_51_79_groupi_n_6739 ,csa_tree_add_51_79_groupi_n_6740);
  not csa_tree_add_51_79_groupi_g39357(csa_tree_add_51_79_groupi_n_6736 ,csa_tree_add_51_79_groupi_n_6735);
  not csa_tree_add_51_79_groupi_g39358(csa_tree_add_51_79_groupi_n_6732 ,csa_tree_add_51_79_groupi_n_6731);
  not csa_tree_add_51_79_groupi_g39359(csa_tree_add_51_79_groupi_n_6730 ,csa_tree_add_51_79_groupi_n_6729);
  not csa_tree_add_51_79_groupi_g39360(csa_tree_add_51_79_groupi_n_6726 ,csa_tree_add_51_79_groupi_n_6725);
  not csa_tree_add_51_79_groupi_g39361(csa_tree_add_51_79_groupi_n_6724 ,csa_tree_add_51_79_groupi_n_6723);
  not csa_tree_add_51_79_groupi_g39362(csa_tree_add_51_79_groupi_n_6721 ,csa_tree_add_51_79_groupi_n_6722);
  not csa_tree_add_51_79_groupi_g39363(csa_tree_add_51_79_groupi_n_6719 ,csa_tree_add_51_79_groupi_n_6720);
  or csa_tree_add_51_79_groupi_g39364(csa_tree_add_51_79_groupi_n_6718 ,csa_tree_add_51_79_groupi_n_5472 ,csa_tree_add_51_79_groupi_n_5720);
  or csa_tree_add_51_79_groupi_g39365(csa_tree_add_51_79_groupi_n_6717 ,csa_tree_add_51_79_groupi_n_5538 ,csa_tree_add_51_79_groupi_n_5711);
  nor csa_tree_add_51_79_groupi_g39366(csa_tree_add_51_79_groupi_n_6716 ,csa_tree_add_51_79_groupi_n_5555 ,csa_tree_add_51_79_groupi_n_6113);
  or csa_tree_add_51_79_groupi_g39367(csa_tree_add_51_79_groupi_n_6715 ,csa_tree_add_51_79_groupi_n_5532 ,csa_tree_add_51_79_groupi_n_6110);
  or csa_tree_add_51_79_groupi_g39368(csa_tree_add_51_79_groupi_n_6714 ,csa_tree_add_51_79_groupi_n_5565 ,csa_tree_add_51_79_groupi_n_6115);
  or csa_tree_add_51_79_groupi_g39369(csa_tree_add_51_79_groupi_n_6713 ,csa_tree_add_51_79_groupi_n_5120 ,csa_tree_add_51_79_groupi_n_5803);
  or csa_tree_add_51_79_groupi_g39370(csa_tree_add_51_79_groupi_n_6712 ,csa_tree_add_51_79_groupi_n_5531 ,csa_tree_add_51_79_groupi_n_6108);
  or csa_tree_add_51_79_groupi_g39371(csa_tree_add_51_79_groupi_n_6711 ,csa_tree_add_51_79_groupi_n_5529 ,csa_tree_add_51_79_groupi_n_6103);
  or csa_tree_add_51_79_groupi_g39372(csa_tree_add_51_79_groupi_n_6710 ,csa_tree_add_51_79_groupi_n_5515 ,csa_tree_add_51_79_groupi_n_6100);
  or csa_tree_add_51_79_groupi_g39373(csa_tree_add_51_79_groupi_n_6709 ,csa_tree_add_51_79_groupi_n_5495 ,csa_tree_add_51_79_groupi_n_6098);
  or csa_tree_add_51_79_groupi_g39374(csa_tree_add_51_79_groupi_n_6708 ,csa_tree_add_51_79_groupi_n_5492 ,csa_tree_add_51_79_groupi_n_6096);
  or csa_tree_add_51_79_groupi_g39375(csa_tree_add_51_79_groupi_n_6707 ,csa_tree_add_51_79_groupi_n_5490 ,csa_tree_add_51_79_groupi_n_6086);
  or csa_tree_add_51_79_groupi_g39376(csa_tree_add_51_79_groupi_n_6706 ,csa_tree_add_51_79_groupi_n_5488 ,csa_tree_add_51_79_groupi_n_6093);
  or csa_tree_add_51_79_groupi_g39377(csa_tree_add_51_79_groupi_n_6705 ,csa_tree_add_51_79_groupi_n_5489 ,csa_tree_add_51_79_groupi_n_6088);
  or csa_tree_add_51_79_groupi_g39378(csa_tree_add_51_79_groupi_n_6704 ,csa_tree_add_51_79_groupi_n_5030 ,csa_tree_add_51_79_groupi_n_6091);
  or csa_tree_add_51_79_groupi_g39379(csa_tree_add_51_79_groupi_n_6703 ,csa_tree_add_51_79_groupi_n_5072 ,csa_tree_add_51_79_groupi_n_6089);
  or csa_tree_add_51_79_groupi_g39380(csa_tree_add_51_79_groupi_n_6702 ,csa_tree_add_51_79_groupi_n_5479 ,csa_tree_add_51_79_groupi_n_6081);
  or csa_tree_add_51_79_groupi_g39381(csa_tree_add_51_79_groupi_n_6701 ,csa_tree_add_51_79_groupi_n_5480 ,csa_tree_add_51_79_groupi_n_6083);
  or csa_tree_add_51_79_groupi_g39382(csa_tree_add_51_79_groupi_n_6700 ,csa_tree_add_51_79_groupi_n_5477 ,csa_tree_add_51_79_groupi_n_6079);
  or csa_tree_add_51_79_groupi_g39383(csa_tree_add_51_79_groupi_n_6699 ,csa_tree_add_51_79_groupi_n_5447 ,csa_tree_add_51_79_groupi_n_6073);
  or csa_tree_add_51_79_groupi_g39384(csa_tree_add_51_79_groupi_n_6698 ,csa_tree_add_51_79_groupi_n_5442 ,csa_tree_add_51_79_groupi_n_6071);
  or csa_tree_add_51_79_groupi_g39385(csa_tree_add_51_79_groupi_n_6697 ,csa_tree_add_51_79_groupi_n_5576 ,csa_tree_add_51_79_groupi_n_6069);
  or csa_tree_add_51_79_groupi_g39386(csa_tree_add_51_79_groupi_n_6696 ,csa_tree_add_51_79_groupi_n_5575 ,csa_tree_add_51_79_groupi_n_6067);
  or csa_tree_add_51_79_groupi_g39387(csa_tree_add_51_79_groupi_n_6695 ,csa_tree_add_51_79_groupi_n_5574 ,csa_tree_add_51_79_groupi_n_6066);
  or csa_tree_add_51_79_groupi_g39388(csa_tree_add_51_79_groupi_n_6694 ,csa_tree_add_51_79_groupi_n_5012 ,csa_tree_add_51_79_groupi_n_6064);
  and csa_tree_add_51_79_groupi_g39389(csa_tree_add_51_79_groupi_n_6693 ,csa_tree_add_51_79_groupi_n_5014 ,csa_tree_add_51_79_groupi_n_5953);
  or csa_tree_add_51_79_groupi_g39390(csa_tree_add_51_79_groupi_n_6692 ,csa_tree_add_51_79_groupi_n_5572 ,csa_tree_add_51_79_groupi_n_6062);
  or csa_tree_add_51_79_groupi_g39391(csa_tree_add_51_79_groupi_n_6691 ,csa_tree_add_51_79_groupi_n_5111 ,csa_tree_add_51_79_groupi_n_6060);
  or csa_tree_add_51_79_groupi_g39392(csa_tree_add_51_79_groupi_n_6690 ,csa_tree_add_51_79_groupi_n_5570 ,csa_tree_add_51_79_groupi_n_6057);
  or csa_tree_add_51_79_groupi_g39393(csa_tree_add_51_79_groupi_n_6689 ,csa_tree_add_51_79_groupi_n_5573 ,csa_tree_add_51_79_groupi_n_6054);
  or csa_tree_add_51_79_groupi_g39394(csa_tree_add_51_79_groupi_n_6688 ,csa_tree_add_51_79_groupi_n_5450 ,csa_tree_add_51_79_groupi_n_6055);
  nor csa_tree_add_51_79_groupi_g39395(csa_tree_add_51_79_groupi_n_6687 ,csa_tree_add_51_79_groupi_n_5577 ,csa_tree_add_51_79_groupi_n_6028);
  or csa_tree_add_51_79_groupi_g39396(csa_tree_add_51_79_groupi_n_6686 ,csa_tree_add_51_79_groupi_n_5475 ,csa_tree_add_51_79_groupi_n_6052);
  or csa_tree_add_51_79_groupi_g39397(csa_tree_add_51_79_groupi_n_6685 ,csa_tree_add_51_79_groupi_n_5013 ,csa_tree_add_51_79_groupi_n_5916);
  or csa_tree_add_51_79_groupi_g39398(csa_tree_add_51_79_groupi_n_6684 ,csa_tree_add_51_79_groupi_n_5514 ,csa_tree_add_51_79_groupi_n_6047);
  or csa_tree_add_51_79_groupi_g39399(csa_tree_add_51_79_groupi_n_6683 ,csa_tree_add_51_79_groupi_n_5568 ,csa_tree_add_51_79_groupi_n_6046);
  or csa_tree_add_51_79_groupi_g39400(csa_tree_add_51_79_groupi_n_6682 ,csa_tree_add_51_79_groupi_n_5569 ,csa_tree_add_51_79_groupi_n_6044);
  or csa_tree_add_51_79_groupi_g39401(csa_tree_add_51_79_groupi_n_6681 ,csa_tree_add_51_79_groupi_n_5566 ,csa_tree_add_51_79_groupi_n_6039);
  nor csa_tree_add_51_79_groupi_g39402(csa_tree_add_51_79_groupi_n_6680 ,csa_tree_add_51_79_groupi_n_5567 ,csa_tree_add_51_79_groupi_n_6037);
  nor csa_tree_add_51_79_groupi_g39403(csa_tree_add_51_79_groupi_n_6679 ,csa_tree_add_51_79_groupi_n_1069 ,csa_tree_add_51_79_groupi_n_5848);
  or csa_tree_add_51_79_groupi_g39404(csa_tree_add_51_79_groupi_n_6678 ,csa_tree_add_51_79_groupi_n_5561 ,csa_tree_add_51_79_groupi_n_5812);
  or csa_tree_add_51_79_groupi_g39405(csa_tree_add_51_79_groupi_n_6677 ,csa_tree_add_51_79_groupi_n_5560 ,csa_tree_add_51_79_groupi_n_6035);
  or csa_tree_add_51_79_groupi_g39406(csa_tree_add_51_79_groupi_n_6676 ,csa_tree_add_51_79_groupi_n_5439 ,csa_tree_add_51_79_groupi_n_6032);
  or csa_tree_add_51_79_groupi_g39407(csa_tree_add_51_79_groupi_n_6675 ,csa_tree_add_51_79_groupi_n_5557 ,csa_tree_add_51_79_groupi_n_6030);
  or csa_tree_add_51_79_groupi_g39408(csa_tree_add_51_79_groupi_n_6674 ,csa_tree_add_51_79_groupi_n_5523 ,csa_tree_add_51_79_groupi_n_5718);
  and csa_tree_add_51_79_groupi_g39409(csa_tree_add_51_79_groupi_n_6673 ,csa_tree_add_51_79_groupi_n_5023 ,csa_tree_add_51_79_groupi_n_5910);
  or csa_tree_add_51_79_groupi_g39410(csa_tree_add_51_79_groupi_n_6672 ,csa_tree_add_51_79_groupi_n_5553 ,csa_tree_add_51_79_groupi_n_6025);
  or csa_tree_add_51_79_groupi_g39411(csa_tree_add_51_79_groupi_n_6671 ,csa_tree_add_51_79_groupi_n_5552 ,csa_tree_add_51_79_groupi_n_6022);
  or csa_tree_add_51_79_groupi_g39412(csa_tree_add_51_79_groupi_n_6670 ,csa_tree_add_51_79_groupi_n_4711 ,csa_tree_add_51_79_groupi_n_5870);
  or csa_tree_add_51_79_groupi_g39413(csa_tree_add_51_79_groupi_n_6669 ,csa_tree_add_51_79_groupi_n_5554 ,csa_tree_add_51_79_groupi_n_6027);
  or csa_tree_add_51_79_groupi_g39414(csa_tree_add_51_79_groupi_n_6668 ,csa_tree_add_51_79_groupi_n_5550 ,csa_tree_add_51_79_groupi_n_6019);
  or csa_tree_add_51_79_groupi_g39415(csa_tree_add_51_79_groupi_n_6667 ,csa_tree_add_51_79_groupi_n_5551 ,csa_tree_add_51_79_groupi_n_6016);
  or csa_tree_add_51_79_groupi_g39416(csa_tree_add_51_79_groupi_n_6666 ,csa_tree_add_51_79_groupi_n_5548 ,csa_tree_add_51_79_groupi_n_6014);
  or csa_tree_add_51_79_groupi_g39417(csa_tree_add_51_79_groupi_n_6665 ,csa_tree_add_51_79_groupi_n_5547 ,csa_tree_add_51_79_groupi_n_6011);
  or csa_tree_add_51_79_groupi_g39418(csa_tree_add_51_79_groupi_n_6664 ,csa_tree_add_51_79_groupi_n_5546 ,csa_tree_add_51_79_groupi_n_6012);
  or csa_tree_add_51_79_groupi_g39419(csa_tree_add_51_79_groupi_n_6663 ,csa_tree_add_51_79_groupi_n_5542 ,csa_tree_add_51_79_groupi_n_6007);
  or csa_tree_add_51_79_groupi_g39420(csa_tree_add_51_79_groupi_n_6662 ,csa_tree_add_51_79_groupi_n_5541 ,csa_tree_add_51_79_groupi_n_6005);
  or csa_tree_add_51_79_groupi_g39421(csa_tree_add_51_79_groupi_n_6661 ,csa_tree_add_51_79_groupi_n_5015 ,csa_tree_add_51_79_groupi_n_6004);
  or csa_tree_add_51_79_groupi_g39422(csa_tree_add_51_79_groupi_n_6660 ,csa_tree_add_51_79_groupi_n_5543 ,csa_tree_add_51_79_groupi_n_6010);
  or csa_tree_add_51_79_groupi_g39423(csa_tree_add_51_79_groupi_n_6659 ,csa_tree_add_51_79_groupi_n_5540 ,csa_tree_add_51_79_groupi_n_6000);
  or csa_tree_add_51_79_groupi_g39424(csa_tree_add_51_79_groupi_n_6658 ,csa_tree_add_51_79_groupi_n_5539 ,csa_tree_add_51_79_groupi_n_5997);
  or csa_tree_add_51_79_groupi_g39425(csa_tree_add_51_79_groupi_n_6657 ,csa_tree_add_51_79_groupi_n_5491 ,csa_tree_add_51_79_groupi_n_5995);
  or csa_tree_add_51_79_groupi_g39426(csa_tree_add_51_79_groupi_n_6656 ,csa_tree_add_51_79_groupi_n_5519 ,csa_tree_add_51_79_groupi_n_5992);
  or csa_tree_add_51_79_groupi_g39427(csa_tree_add_51_79_groupi_n_6655 ,csa_tree_add_51_79_groupi_n_5537 ,csa_tree_add_51_79_groupi_n_5993);
  or csa_tree_add_51_79_groupi_g39428(csa_tree_add_51_79_groupi_n_6654 ,csa_tree_add_51_79_groupi_n_5016 ,csa_tree_add_51_79_groupi_n_5989);
  or csa_tree_add_51_79_groupi_g39429(csa_tree_add_51_79_groupi_n_6653 ,csa_tree_add_51_79_groupi_n_5536 ,csa_tree_add_51_79_groupi_n_5986);
  and csa_tree_add_51_79_groupi_g39430(csa_tree_add_51_79_groupi_n_6652 ,csa_tree_add_51_79_groupi_n_5031 ,csa_tree_add_51_79_groupi_n_5621);
  or csa_tree_add_51_79_groupi_g39431(csa_tree_add_51_79_groupi_n_6651 ,csa_tree_add_51_79_groupi_n_5535 ,csa_tree_add_51_79_groupi_n_5983);
  or csa_tree_add_51_79_groupi_g39432(csa_tree_add_51_79_groupi_n_6650 ,csa_tree_add_51_79_groupi_n_5533 ,csa_tree_add_51_79_groupi_n_5981);
  or csa_tree_add_51_79_groupi_g39433(csa_tree_add_51_79_groupi_n_6649 ,csa_tree_add_51_79_groupi_n_6144 ,csa_tree_add_51_79_groupi_n_6138);
  or csa_tree_add_51_79_groupi_g39434(csa_tree_add_51_79_groupi_n_6648 ,csa_tree_add_51_79_groupi_n_5530 ,csa_tree_add_51_79_groupi_n_5977);
  and csa_tree_add_51_79_groupi_g39435(csa_tree_add_51_79_groupi_n_6647 ,csa_tree_add_51_79_groupi_n_6144 ,csa_tree_add_51_79_groupi_n_6138);
  or csa_tree_add_51_79_groupi_g39436(csa_tree_add_51_79_groupi_n_6646 ,csa_tree_add_51_79_groupi_n_5564 ,csa_tree_add_51_79_groupi_n_5813);
  or csa_tree_add_51_79_groupi_g39437(csa_tree_add_51_79_groupi_n_6645 ,csa_tree_add_51_79_groupi_n_5528 ,csa_tree_add_51_79_groupi_n_5970);
  or csa_tree_add_51_79_groupi_g39438(csa_tree_add_51_79_groupi_n_6644 ,csa_tree_add_51_79_groupi_n_5017 ,csa_tree_add_51_79_groupi_n_5975);
  or csa_tree_add_51_79_groupi_g39439(csa_tree_add_51_79_groupi_n_6643 ,csa_tree_add_51_79_groupi_n_5527 ,csa_tree_add_51_79_groupi_n_5792);
  or csa_tree_add_51_79_groupi_g39440(csa_tree_add_51_79_groupi_n_6642 ,csa_tree_add_51_79_groupi_n_5526 ,csa_tree_add_51_79_groupi_n_5971);
  or csa_tree_add_51_79_groupi_g39441(csa_tree_add_51_79_groupi_n_6641 ,csa_tree_add_51_79_groupi_n_5524 ,csa_tree_add_51_79_groupi_n_5920);
  nor csa_tree_add_51_79_groupi_g39442(csa_tree_add_51_79_groupi_n_6640 ,csa_tree_add_51_79_groupi_n_5510 ,csa_tree_add_51_79_groupi_n_5966);
  or csa_tree_add_51_79_groupi_g39443(csa_tree_add_51_79_groupi_n_6639 ,csa_tree_add_51_79_groupi_n_5461 ,csa_tree_add_51_79_groupi_n_5791);
  or csa_tree_add_51_79_groupi_g39444(csa_tree_add_51_79_groupi_n_6638 ,csa_tree_add_51_79_groupi_n_6151 ,csa_tree_add_51_79_groupi_n_5676);
  or csa_tree_add_51_79_groupi_g39445(csa_tree_add_51_79_groupi_n_6637 ,csa_tree_add_51_79_groupi_n_5053 ,csa_tree_add_51_79_groupi_n_6040);
  or csa_tree_add_51_79_groupi_g39446(csa_tree_add_51_79_groupi_n_6636 ,csa_tree_add_51_79_groupi_n_5522 ,csa_tree_add_51_79_groupi_n_5926);
  or csa_tree_add_51_79_groupi_g39447(csa_tree_add_51_79_groupi_n_6635 ,csa_tree_add_51_79_groupi_n_5521 ,csa_tree_add_51_79_groupi_n_5961);
  nor csa_tree_add_51_79_groupi_g39448(csa_tree_add_51_79_groupi_n_6634 ,csa_tree_add_51_79_groupi_n_5401 ,csa_tree_add_51_79_groupi_n_6142);
  or csa_tree_add_51_79_groupi_g39449(csa_tree_add_51_79_groupi_n_6633 ,csa_tree_add_51_79_groupi_n_5520 ,csa_tree_add_51_79_groupi_n_5957);
  or csa_tree_add_51_79_groupi_g39450(csa_tree_add_51_79_groupi_n_6632 ,csa_tree_add_51_79_groupi_n_5032 ,csa_tree_add_51_79_groupi_n_5778);
  or csa_tree_add_51_79_groupi_g39451(csa_tree_add_51_79_groupi_n_6631 ,csa_tree_add_51_79_groupi_n_5400 ,csa_tree_add_51_79_groupi_n_6143);
  or csa_tree_add_51_79_groupi_g39452(csa_tree_add_51_79_groupi_n_6630 ,csa_tree_add_51_79_groupi_n_5062 ,csa_tree_add_51_79_groupi_n_5955);
  or csa_tree_add_51_79_groupi_g39453(csa_tree_add_51_79_groupi_n_6629 ,csa_tree_add_51_79_groupi_n_5116 ,csa_tree_add_51_79_groupi_n_5952);
  or csa_tree_add_51_79_groupi_g39454(csa_tree_add_51_79_groupi_n_6628 ,csa_tree_add_51_79_groupi_n_5082 ,csa_tree_add_51_79_groupi_n_5598);
  or csa_tree_add_51_79_groupi_g39455(csa_tree_add_51_79_groupi_n_6627 ,csa_tree_add_51_79_groupi_n_5028 ,csa_tree_add_51_79_groupi_n_5950);
  or csa_tree_add_51_79_groupi_g39456(csa_tree_add_51_79_groupi_n_6626 ,csa_tree_add_51_79_groupi_n_5511 ,csa_tree_add_51_79_groupi_n_5943);
  or csa_tree_add_51_79_groupi_g39457(csa_tree_add_51_79_groupi_n_6625 ,csa_tree_add_51_79_groupi_n_5512 ,csa_tree_add_51_79_groupi_n_5946);
  or csa_tree_add_51_79_groupi_g39458(csa_tree_add_51_79_groupi_n_6624 ,csa_tree_add_51_79_groupi_n_5019 ,csa_tree_add_51_79_groupi_n_5941);
  and csa_tree_add_51_79_groupi_g39459(csa_tree_add_51_79_groupi_n_6623 ,csa_tree_add_51_79_groupi_n_5022 ,csa_tree_add_51_79_groupi_n_5935);
  or csa_tree_add_51_79_groupi_g39460(csa_tree_add_51_79_groupi_n_6622 ,csa_tree_add_51_79_groupi_n_5020 ,csa_tree_add_51_79_groupi_n_5938);
  or csa_tree_add_51_79_groupi_g39461(csa_tree_add_51_79_groupi_n_6621 ,csa_tree_add_51_79_groupi_n_5507 ,csa_tree_add_51_79_groupi_n_5933);
  or csa_tree_add_51_79_groupi_g39462(csa_tree_add_51_79_groupi_n_6620 ,csa_tree_add_51_79_groupi_n_5506 ,csa_tree_add_51_79_groupi_n_5929);
  or csa_tree_add_51_79_groupi_g39463(csa_tree_add_51_79_groupi_n_6619 ,csa_tree_add_51_79_groupi_n_5505 ,csa_tree_add_51_79_groupi_n_5931);
  or csa_tree_add_51_79_groupi_g39464(csa_tree_add_51_79_groupi_n_6618 ,csa_tree_add_51_79_groupi_n_5504 ,csa_tree_add_51_79_groupi_n_5928);
  or csa_tree_add_51_79_groupi_g39465(csa_tree_add_51_79_groupi_n_6617 ,csa_tree_add_51_79_groupi_n_5065 ,csa_tree_add_51_79_groupi_n_5763);
  or csa_tree_add_51_79_groupi_g39466(csa_tree_add_51_79_groupi_n_6616 ,csa_tree_add_51_79_groupi_n_5503 ,csa_tree_add_51_79_groupi_n_5924);
  or csa_tree_add_51_79_groupi_g39467(csa_tree_add_51_79_groupi_n_6615 ,csa_tree_add_51_79_groupi_n_5501 ,csa_tree_add_51_79_groupi_n_5921);
  or csa_tree_add_51_79_groupi_g39468(csa_tree_add_51_79_groupi_n_6614 ,csa_tree_add_51_79_groupi_n_5089 ,csa_tree_add_51_79_groupi_n_5709);
  or csa_tree_add_51_79_groupi_g39469(csa_tree_add_51_79_groupi_n_6613 ,csa_tree_add_51_79_groupi_n_5498 ,csa_tree_add_51_79_groupi_n_5919);
  or csa_tree_add_51_79_groupi_g39470(csa_tree_add_51_79_groupi_n_6612 ,csa_tree_add_51_79_groupi_n_5021 ,csa_tree_add_51_79_groupi_n_5705);
  or csa_tree_add_51_79_groupi_g39471(csa_tree_add_51_79_groupi_n_6611 ,csa_tree_add_51_79_groupi_n_5525 ,csa_tree_add_51_79_groupi_n_5987);
  or csa_tree_add_51_79_groupi_g39472(csa_tree_add_51_79_groupi_n_6610 ,csa_tree_add_51_79_groupi_n_5544 ,csa_tree_add_51_79_groupi_n_5909);
  or csa_tree_add_51_79_groupi_g39473(csa_tree_add_51_79_groupi_n_6609 ,csa_tree_add_51_79_groupi_n_5496 ,csa_tree_add_51_79_groupi_n_5912);
  or csa_tree_add_51_79_groupi_g39474(csa_tree_add_51_79_groupi_n_6608 ,csa_tree_add_51_79_groupi_n_5301 ,csa_tree_add_51_79_groupi_n_6139);
  or csa_tree_add_51_79_groupi_g39475(csa_tree_add_51_79_groupi_n_6607 ,csa_tree_add_51_79_groupi_n_5068 ,csa_tree_add_51_79_groupi_n_5608);
  or csa_tree_add_51_79_groupi_g39476(csa_tree_add_51_79_groupi_n_6606 ,csa_tree_add_51_79_groupi_n_5494 ,csa_tree_add_51_79_groupi_n_5908);
  or csa_tree_add_51_79_groupi_g39477(csa_tree_add_51_79_groupi_n_6605 ,csa_tree_add_51_79_groupi_n_5493 ,csa_tree_add_51_79_groupi_n_5903);
  or csa_tree_add_51_79_groupi_g39478(csa_tree_add_51_79_groupi_n_6604 ,csa_tree_add_51_79_groupi_n_5024 ,csa_tree_add_51_79_groupi_n_5907);
  or csa_tree_add_51_79_groupi_g39479(csa_tree_add_51_79_groupi_n_6603 ,csa_tree_add_51_79_groupi_n_5112 ,csa_tree_add_51_79_groupi_n_5889);
  or csa_tree_add_51_79_groupi_g39480(csa_tree_add_51_79_groupi_n_6602 ,csa_tree_add_51_79_groupi_n_5025 ,csa_tree_add_51_79_groupi_n_5904);
  and csa_tree_add_51_79_groupi_g39481(csa_tree_add_51_79_groupi_n_6601 ,csa_tree_add_51_79_groupi_n_5063 ,csa_tree_add_51_79_groupi_n_5969);
  or csa_tree_add_51_79_groupi_g39482(csa_tree_add_51_79_groupi_n_6600 ,csa_tree_add_51_79_groupi_n_5100 ,csa_tree_add_51_79_groupi_n_5899);
  or csa_tree_add_51_79_groupi_g39483(csa_tree_add_51_79_groupi_n_6599 ,csa_tree_add_51_79_groupi_n_6132 ,csa_tree_add_51_79_groupi_n_6137);
  and csa_tree_add_51_79_groupi_g39484(csa_tree_add_51_79_groupi_n_6598 ,csa_tree_add_51_79_groupi_n_6132 ,csa_tree_add_51_79_groupi_n_6137);
  or csa_tree_add_51_79_groupi_g39485(csa_tree_add_51_79_groupi_n_6597 ,csa_tree_add_51_79_groupi_n_5440 ,csa_tree_add_51_79_groupi_n_5805);
  or csa_tree_add_51_79_groupi_g39486(csa_tree_add_51_79_groupi_n_6596 ,csa_tree_add_51_79_groupi_n_5457 ,csa_tree_add_51_79_groupi_n_5892);
  or csa_tree_add_51_79_groupi_g39487(csa_tree_add_51_79_groupi_n_6595 ,csa_tree_add_51_79_groupi_n_5486 ,csa_tree_add_51_79_groupi_n_5890);
  or csa_tree_add_51_79_groupi_g39488(csa_tree_add_51_79_groupi_n_6594 ,csa_tree_add_51_79_groupi_n_5485 ,csa_tree_add_51_79_groupi_n_5883);
  or csa_tree_add_51_79_groupi_g39489(csa_tree_add_51_79_groupi_n_6593 ,csa_tree_add_51_79_groupi_n_5484 ,csa_tree_add_51_79_groupi_n_5880);
  and csa_tree_add_51_79_groupi_g39490(csa_tree_add_51_79_groupi_n_6592 ,csa_tree_add_51_79_groupi_n_5301 ,csa_tree_add_51_79_groupi_n_6139);
  or csa_tree_add_51_79_groupi_g39491(csa_tree_add_51_79_groupi_n_6591 ,csa_tree_add_51_79_groupi_n_5435 ,csa_tree_add_51_79_groupi_n_5898);
  or csa_tree_add_51_79_groupi_g39492(csa_tree_add_51_79_groupi_n_6590 ,csa_tree_add_51_79_groupi_n_5516 ,csa_tree_add_51_79_groupi_n_5874);
  or csa_tree_add_51_79_groupi_g39493(csa_tree_add_51_79_groupi_n_6589 ,csa_tree_add_51_79_groupi_n_5483 ,csa_tree_add_51_79_groupi_n_5871);
  or csa_tree_add_51_79_groupi_g39494(csa_tree_add_51_79_groupi_n_6588 ,csa_tree_add_51_79_groupi_n_5482 ,csa_tree_add_51_79_groupi_n_5887);
  or csa_tree_add_51_79_groupi_g39495(csa_tree_add_51_79_groupi_n_6587 ,csa_tree_add_51_79_groupi_n_5481 ,csa_tree_add_51_79_groupi_n_5897);
  or csa_tree_add_51_79_groupi_g39496(csa_tree_add_51_79_groupi_n_6586 ,csa_tree_add_51_79_groupi_n_5860 ,csa_tree_add_51_79_groupi_n_6140);
  or csa_tree_add_51_79_groupi_g39497(csa_tree_add_51_79_groupi_n_6585 ,csa_tree_add_51_79_groupi_n_5478 ,csa_tree_add_51_79_groupi_n_5902);
  and csa_tree_add_51_79_groupi_g39498(csa_tree_add_51_79_groupi_n_6584 ,csa_tree_add_51_79_groupi_n_5860 ,csa_tree_add_51_79_groupi_n_6140);
  or csa_tree_add_51_79_groupi_g39499(csa_tree_add_51_79_groupi_n_6583 ,csa_tree_add_51_79_groupi_n_5476 ,csa_tree_add_51_79_groupi_n_5873);
  or csa_tree_add_51_79_groupi_g39500(csa_tree_add_51_79_groupi_n_6582 ,csa_tree_add_51_79_groupi_n_5044 ,csa_tree_add_51_79_groupi_n_6114);
  or csa_tree_add_51_79_groupi_g39501(csa_tree_add_51_79_groupi_n_6581 ,csa_tree_add_51_79_groupi_n_5562 ,csa_tree_add_51_79_groupi_n_5973);
  or csa_tree_add_51_79_groupi_g39502(csa_tree_add_51_79_groupi_n_6580 ,csa_tree_add_51_79_groupi_n_5067 ,csa_tree_add_51_79_groupi_n_5602);
  or csa_tree_add_51_79_groupi_g39503(csa_tree_add_51_79_groupi_n_6579 ,csa_tree_add_51_79_groupi_n_5473 ,csa_tree_add_51_79_groupi_n_6033);
  or csa_tree_add_51_79_groupi_g39504(csa_tree_add_51_79_groupi_n_6578 ,csa_tree_add_51_79_groupi_n_5474 ,csa_tree_add_51_79_groupi_n_5978);
  or csa_tree_add_51_79_groupi_g39505(csa_tree_add_51_79_groupi_n_6577 ,csa_tree_add_51_79_groupi_n_5471 ,csa_tree_add_51_79_groupi_n_6076);
  and csa_tree_add_51_79_groupi_g39506(csa_tree_add_51_79_groupi_n_6576 ,csa_tree_add_51_79_groupi_n_5033 ,csa_tree_add_51_79_groupi_n_6085);
  or csa_tree_add_51_79_groupi_g39507(csa_tree_add_51_79_groupi_n_6575 ,csa_tree_add_51_79_groupi_n_5470 ,csa_tree_add_51_79_groupi_n_6117);
  or csa_tree_add_51_79_groupi_g39508(csa_tree_add_51_79_groupi_n_6574 ,csa_tree_add_51_79_groupi_n_5508 ,csa_tree_add_51_79_groupi_n_6124);
  or csa_tree_add_51_79_groupi_g39509(csa_tree_add_51_79_groupi_n_6573 ,csa_tree_add_51_79_groupi_n_5036 ,csa_tree_add_51_79_groupi_n_5836);
  or csa_tree_add_51_79_groupi_g39510(csa_tree_add_51_79_groupi_n_6572 ,csa_tree_add_51_79_groupi_n_5078 ,csa_tree_add_51_79_groupi_n_5835);
  or csa_tree_add_51_79_groupi_g39511(csa_tree_add_51_79_groupi_n_6571 ,csa_tree_add_51_79_groupi_n_5465 ,csa_tree_add_51_79_groupi_n_5917);
  or csa_tree_add_51_79_groupi_g39512(csa_tree_add_51_79_groupi_n_6570 ,csa_tree_add_51_79_groupi_n_5467 ,csa_tree_add_51_79_groupi_n_5832);
  or csa_tree_add_51_79_groupi_g39513(csa_tree_add_51_79_groupi_n_6569 ,csa_tree_add_51_79_groupi_n_5037 ,csa_tree_add_51_79_groupi_n_5829);
  or csa_tree_add_51_79_groupi_g39514(csa_tree_add_51_79_groupi_n_6568 ,csa_tree_add_51_79_groupi_n_5102 ,csa_tree_add_51_79_groupi_n_5828);
  or csa_tree_add_51_79_groupi_g39515(csa_tree_add_51_79_groupi_n_6567 ,csa_tree_add_51_79_groupi_n_5039 ,csa_tree_add_51_79_groupi_n_5826);
  or csa_tree_add_51_79_groupi_g39516(csa_tree_add_51_79_groupi_n_6566 ,csa_tree_add_51_79_groupi_n_5464 ,csa_tree_add_51_79_groupi_n_5823);
  or csa_tree_add_51_79_groupi_g39517(csa_tree_add_51_79_groupi_n_6565 ,csa_tree_add_51_79_groupi_n_5041 ,csa_tree_add_51_79_groupi_n_5824);
  or csa_tree_add_51_79_groupi_g39518(csa_tree_add_51_79_groupi_n_6564 ,csa_tree_add_51_79_groupi_n_5455 ,csa_tree_add_51_79_groupi_n_5876);
  or csa_tree_add_51_79_groupi_g39519(csa_tree_add_51_79_groupi_n_6563 ,csa_tree_add_51_79_groupi_n_5043 ,csa_tree_add_51_79_groupi_n_5821);
  or csa_tree_add_51_79_groupi_g39520(csa_tree_add_51_79_groupi_n_6562 ,csa_tree_add_51_79_groupi_n_5101 ,csa_tree_add_51_79_groupi_n_5715);
  or csa_tree_add_51_79_groupi_g39521(csa_tree_add_51_79_groupi_n_6561 ,csa_tree_add_51_79_groupi_n_5462 ,csa_tree_add_51_79_groupi_n_5818);
  nor csa_tree_add_51_79_groupi_g39522(csa_tree_add_51_79_groupi_n_6560 ,csa_tree_add_51_79_groupi_n_5451 ,csa_tree_add_51_79_groupi_n_5745);
  or csa_tree_add_51_79_groupi_g39523(csa_tree_add_51_79_groupi_n_6559 ,csa_tree_add_51_79_groupi_n_5500 ,csa_tree_add_51_79_groupi_n_5708);
  or csa_tree_add_51_79_groupi_g39524(csa_tree_add_51_79_groupi_n_6558 ,csa_tree_add_51_79_groupi_n_5459 ,csa_tree_add_51_79_groupi_n_5712);
  or csa_tree_add_51_79_groupi_g39525(csa_tree_add_51_79_groupi_n_6557 ,csa_tree_add_51_79_groupi_n_5077 ,csa_tree_add_51_79_groupi_n_5688);
  or csa_tree_add_51_79_groupi_g39526(csa_tree_add_51_79_groupi_n_6556 ,csa_tree_add_51_79_groupi_n_5018 ,csa_tree_add_51_79_groupi_n_5808);
  or csa_tree_add_51_79_groupi_g39527(csa_tree_add_51_79_groupi_n_6555 ,csa_tree_add_51_79_groupi_n_5011 ,csa_tree_add_51_79_groupi_n_6077);
  or csa_tree_add_51_79_groupi_g39528(csa_tree_add_51_79_groupi_n_6554 ,csa_tree_add_51_79_groupi_n_5460 ,csa_tree_add_51_79_groupi_n_5793);
  or csa_tree_add_51_79_groupi_g39529(csa_tree_add_51_79_groupi_n_6553 ,csa_tree_add_51_79_groupi_n_5069 ,csa_tree_add_51_79_groupi_n_5615);
  or csa_tree_add_51_79_groupi_g39530(csa_tree_add_51_79_groupi_n_6552 ,csa_tree_add_51_79_groupi_n_5469 ,csa_tree_add_51_79_groupi_n_6082);
  or csa_tree_add_51_79_groupi_g39531(csa_tree_add_51_79_groupi_n_6551 ,csa_tree_add_51_79_groupi_n_5449 ,csa_tree_add_51_79_groupi_n_5800);
  or csa_tree_add_51_79_groupi_g39532(csa_tree_add_51_79_groupi_n_6550 ,csa_tree_add_51_79_groupi_n_5075 ,csa_tree_add_51_79_groupi_n_5716);
  or csa_tree_add_51_79_groupi_g39533(csa_tree_add_51_79_groupi_n_6549 ,csa_tree_add_51_79_groupi_n_5047 ,csa_tree_add_51_79_groupi_n_5795);
  or csa_tree_add_51_79_groupi_g39534(csa_tree_add_51_79_groupi_n_6548 ,csa_tree_add_51_79_groupi_n_5108 ,csa_tree_add_51_79_groupi_n_5752);
  or csa_tree_add_51_79_groupi_g39535(csa_tree_add_51_79_groupi_n_6547 ,csa_tree_add_51_79_groupi_n_5466 ,csa_tree_add_51_79_groupi_n_5834);
  or csa_tree_add_51_79_groupi_g39536(csa_tree_add_51_79_groupi_n_6546 ,csa_tree_add_51_79_groupi_n_5438 ,csa_tree_add_51_79_groupi_n_5632);
  or csa_tree_add_51_79_groupi_g39537(csa_tree_add_51_79_groupi_n_6545 ,csa_tree_add_51_79_groupi_n_5092 ,csa_tree_add_51_79_groupi_n_5789);
  or csa_tree_add_51_79_groupi_g39538(csa_tree_add_51_79_groupi_n_6544 ,csa_tree_add_51_79_groupi_n_5050 ,csa_tree_add_51_79_groupi_n_5788);
  or csa_tree_add_51_79_groupi_g39539(csa_tree_add_51_79_groupi_n_6543 ,csa_tree_add_51_79_groupi_n_5436 ,csa_tree_add_51_79_groupi_n_5724);
  or csa_tree_add_51_79_groupi_g39540(csa_tree_add_51_79_groupi_n_6542 ,csa_tree_add_51_79_groupi_n_5048 ,csa_tree_add_51_79_groupi_n_5944);
  or csa_tree_add_51_79_groupi_g39541(csa_tree_add_51_79_groupi_n_6541 ,csa_tree_add_51_79_groupi_n_5452 ,csa_tree_add_51_79_groupi_n_5807);
  or csa_tree_add_51_79_groupi_g39542(csa_tree_add_51_79_groupi_n_6540 ,csa_tree_add_51_79_groupi_n_6141 ,csa_tree_add_51_79_groupi_n_6129);
  and csa_tree_add_51_79_groupi_g39543(csa_tree_add_51_79_groupi_n_6539 ,csa_tree_add_51_79_groupi_n_6141 ,csa_tree_add_51_79_groupi_n_6129);
  or csa_tree_add_51_79_groupi_g39544(csa_tree_add_51_79_groupi_n_6538 ,csa_tree_add_51_79_groupi_n_1528 ,csa_tree_add_51_79_groupi_n_5847);
  or csa_tree_add_51_79_groupi_g39545(csa_tree_add_51_79_groupi_n_6537 ,csa_tree_add_51_79_groupi_n_5468 ,csa_tree_add_51_79_groupi_n_5770);
  or csa_tree_add_51_79_groupi_g39546(csa_tree_add_51_79_groupi_n_6536 ,csa_tree_add_51_79_groupi_n_5054 ,csa_tree_add_51_79_groupi_n_5771);
  or csa_tree_add_51_79_groupi_g39547(csa_tree_add_51_79_groupi_n_6535 ,csa_tree_add_51_79_groupi_n_5055 ,csa_tree_add_51_79_groupi_n_5769);
  or csa_tree_add_51_79_groupi_g39548(csa_tree_add_51_79_groupi_n_6534 ,csa_tree_add_51_79_groupi_n_5064 ,csa_tree_add_51_79_groupi_n_5604);
  or csa_tree_add_51_79_groupi_g39549(csa_tree_add_51_79_groupi_n_6533 ,csa_tree_add_51_79_groupi_n_5106 ,csa_tree_add_51_79_groupi_n_5762);
  or csa_tree_add_51_79_groupi_g39550(csa_tree_add_51_79_groupi_n_6532 ,csa_tree_add_51_79_groupi_n_5122 ,csa_tree_add_51_79_groupi_n_5759);
  or csa_tree_add_51_79_groupi_g39551(csa_tree_add_51_79_groupi_n_6531 ,csa_tree_add_51_79_groupi_n_5502 ,csa_tree_add_51_79_groupi_n_5757);
  or csa_tree_add_51_79_groupi_g39552(csa_tree_add_51_79_groupi_n_6530 ,csa_tree_add_51_79_groupi_n_5098 ,csa_tree_add_51_79_groupi_n_5758);
  or csa_tree_add_51_79_groupi_g39553(csa_tree_add_51_79_groupi_n_6529 ,csa_tree_add_51_79_groupi_n_5563 ,csa_tree_add_51_79_groupi_n_5960);
  or csa_tree_add_51_79_groupi_g39554(csa_tree_add_51_79_groupi_n_6528 ,csa_tree_add_51_79_groupi_n_5487 ,csa_tree_add_51_79_groupi_n_5796);
  or csa_tree_add_51_79_groupi_g39555(csa_tree_add_51_79_groupi_n_6527 ,csa_tree_add_51_79_groupi_n_5060 ,csa_tree_add_51_79_groupi_n_5610);
  or csa_tree_add_51_79_groupi_g39556(csa_tree_add_51_79_groupi_n_6526 ,csa_tree_add_51_79_groupi_n_5079 ,csa_tree_add_51_79_groupi_n_5748);
  or csa_tree_add_51_79_groupi_g39557(csa_tree_add_51_79_groupi_n_6525 ,csa_tree_add_51_79_groupi_n_5056 ,csa_tree_add_51_79_groupi_n_5597);
  or csa_tree_add_51_79_groupi_g39558(csa_tree_add_51_79_groupi_n_6524 ,csa_tree_add_51_79_groupi_n_5545 ,csa_tree_add_51_79_groupi_n_5706);
  or csa_tree_add_51_79_groupi_g39559(csa_tree_add_51_79_groupi_n_6523 ,csa_tree_add_51_79_groupi_n_5115 ,csa_tree_add_51_79_groupi_n_5784);
  or csa_tree_add_51_79_groupi_g39560(csa_tree_add_51_79_groupi_n_6522 ,csa_tree_add_51_79_groupi_n_5073 ,csa_tree_add_51_79_groupi_n_5600);
  or csa_tree_add_51_79_groupi_g39561(csa_tree_add_51_79_groupi_n_6521 ,csa_tree_add_51_79_groupi_n_5855 ,csa_tree_add_51_79_groupi_n_5857);
  or csa_tree_add_51_79_groupi_g39562(csa_tree_add_51_79_groupi_n_6520 ,csa_tree_add_51_79_groupi_n_5096 ,csa_tree_add_51_79_groupi_n_5742);
  nor csa_tree_add_51_79_groupi_g39563(csa_tree_add_51_79_groupi_n_6519 ,csa_tree_add_51_79_groupi_n_5856 ,csa_tree_add_51_79_groupi_n_5858);
  or csa_tree_add_51_79_groupi_g39564(csa_tree_add_51_79_groupi_n_6518 ,csa_tree_add_51_79_groupi_n_5123 ,csa_tree_add_51_79_groupi_n_5739);
  or csa_tree_add_51_79_groupi_g39565(csa_tree_add_51_79_groupi_n_6517 ,csa_tree_add_51_79_groupi_n_5121 ,csa_tree_add_51_79_groupi_n_5925);
  or csa_tree_add_51_79_groupi_g39566(csa_tree_add_51_79_groupi_n_6516 ,csa_tree_add_51_79_groupi_n_5119 ,csa_tree_add_51_79_groupi_n_5737);
  or csa_tree_add_51_79_groupi_g39567(csa_tree_add_51_79_groupi_n_6515 ,csa_tree_add_51_79_groupi_n_5093 ,csa_tree_add_51_79_groupi_n_5735);
  or csa_tree_add_51_79_groupi_g39568(csa_tree_add_51_79_groupi_n_6514 ,csa_tree_add_51_79_groupi_n_5113 ,csa_tree_add_51_79_groupi_n_5734);
  or csa_tree_add_51_79_groupi_g39569(csa_tree_add_51_79_groupi_n_6513 ,csa_tree_add_51_79_groupi_n_5045 ,csa_tree_add_51_79_groupi_n_5690);
  or csa_tree_add_51_79_groupi_g39570(csa_tree_add_51_79_groupi_n_6512 ,csa_tree_add_51_79_groupi_n_5859 ,csa_tree_add_51_79_groupi_n_5842);
  or csa_tree_add_51_79_groupi_g39571(csa_tree_add_51_79_groupi_n_6511 ,csa_tree_add_51_79_groupi_n_5448 ,csa_tree_add_51_79_groupi_n_5683);
  or csa_tree_add_51_79_groupi_g39572(csa_tree_add_51_79_groupi_n_6510 ,csa_tree_add_51_79_groupi_n_5070 ,csa_tree_add_51_79_groupi_n_5815);
  and csa_tree_add_51_79_groupi_g39573(csa_tree_add_51_79_groupi_n_6509 ,csa_tree_add_51_79_groupi_n_6145 ,csa_tree_add_51_79_groupi_n_6146);
  or csa_tree_add_51_79_groupi_g39574(csa_tree_add_51_79_groupi_n_6508 ,csa_tree_add_51_79_groupi_n_5846 ,csa_tree_add_51_79_groupi_n_5845);
  or csa_tree_add_51_79_groupi_g39575(csa_tree_add_51_79_groupi_n_6507 ,csa_tree_add_51_79_groupi_n_5071 ,csa_tree_add_51_79_groupi_n_5725);
  and csa_tree_add_51_79_groupi_g39576(csa_tree_add_51_79_groupi_n_6506 ,csa_tree_add_51_79_groupi_n_5846 ,csa_tree_add_51_79_groupi_n_5845);
  or csa_tree_add_51_79_groupi_g39577(csa_tree_add_51_79_groupi_n_6505 ,csa_tree_add_51_79_groupi_n_6145 ,csa_tree_add_51_79_groupi_n_6146);
  nor csa_tree_add_51_79_groupi_g39578(csa_tree_add_51_79_groupi_n_6504 ,csa_tree_add_51_79_groupi_n_5446 ,csa_tree_add_51_79_groupi_n_5714);
  or csa_tree_add_51_79_groupi_g39579(csa_tree_add_51_79_groupi_n_6503 ,csa_tree_add_51_79_groupi_n_5105 ,csa_tree_add_51_79_groupi_n_5782);
  or csa_tree_add_51_79_groupi_g39580(csa_tree_add_51_79_groupi_n_6502 ,csa_tree_add_51_79_groupi_n_5513 ,csa_tree_add_51_79_groupi_n_5781);
  or csa_tree_add_51_79_groupi_g39581(csa_tree_add_51_79_groupi_n_6501 ,csa_tree_add_51_79_groupi_n_5125 ,csa_tree_add_51_79_groupi_n_5700);
  or csa_tree_add_51_79_groupi_g39582(csa_tree_add_51_79_groupi_n_6500 ,csa_tree_add_51_79_groupi_n_5124 ,csa_tree_add_51_79_groupi_n_5701);
  or csa_tree_add_51_79_groupi_g39583(csa_tree_add_51_79_groupi_n_6499 ,csa_tree_add_51_79_groupi_n_5081 ,csa_tree_add_51_79_groupi_n_5839);
  or csa_tree_add_51_79_groupi_g39584(csa_tree_add_51_79_groupi_n_6498 ,csa_tree_add_51_79_groupi_n_5497 ,csa_tree_add_51_79_groupi_n_5693);
  or csa_tree_add_51_79_groupi_g39585(csa_tree_add_51_79_groupi_n_6497 ,csa_tree_add_51_79_groupi_n_5118 ,csa_tree_add_51_79_groupi_n_5695);
  or csa_tree_add_51_79_groupi_g39586(csa_tree_add_51_79_groupi_n_6496 ,csa_tree_add_51_79_groupi_n_5114 ,csa_tree_add_51_79_groupi_n_5691);
  and csa_tree_add_51_79_groupi_g39587(csa_tree_add_51_79_groupi_n_6495 ,csa_tree_add_51_79_groupi_n_5859 ,csa_tree_add_51_79_groupi_n_5842);
  or csa_tree_add_51_79_groupi_g39588(csa_tree_add_51_79_groupi_n_6494 ,csa_tree_add_51_79_groupi_n_5110 ,csa_tree_add_51_79_groupi_n_5686);
  nor csa_tree_add_51_79_groupi_g39589(csa_tree_add_51_79_groupi_n_6493 ,csa_tree_add_51_79_groupi_n_5086 ,csa_tree_add_51_79_groupi_n_5635);
  or csa_tree_add_51_79_groupi_g39590(csa_tree_add_51_79_groupi_n_6492 ,csa_tree_add_51_79_groupi_n_5104 ,csa_tree_add_51_79_groupi_n_5681);
  or csa_tree_add_51_79_groupi_g39591(csa_tree_add_51_79_groupi_n_6491 ,csa_tree_add_51_79_groupi_n_5456 ,csa_tree_add_51_79_groupi_n_5810);
  or csa_tree_add_51_79_groupi_g39592(csa_tree_add_51_79_groupi_n_6490 ,csa_tree_add_51_79_groupi_n_5083 ,csa_tree_add_51_79_groupi_n_5679);
  or csa_tree_add_51_79_groupi_g39593(csa_tree_add_51_79_groupi_n_6489 ,csa_tree_add_51_79_groupi_n_5099 ,csa_tree_add_51_79_groupi_n_5675);
  or csa_tree_add_51_79_groupi_g39594(csa_tree_add_51_79_groupi_n_6488 ,csa_tree_add_51_79_groupi_n_5095 ,csa_tree_add_51_79_groupi_n_5672);
  or csa_tree_add_51_79_groupi_g39595(csa_tree_add_51_79_groupi_n_6487 ,csa_tree_add_51_79_groupi_n_5094 ,csa_tree_add_51_79_groupi_n_5671);
  or csa_tree_add_51_79_groupi_g39596(csa_tree_add_51_79_groupi_n_6486 ,csa_tree_add_51_79_groupi_n_5090 ,csa_tree_add_51_79_groupi_n_5667);
  or csa_tree_add_51_79_groupi_g39597(csa_tree_add_51_79_groupi_n_6485 ,csa_tree_add_51_79_groupi_n_5084 ,csa_tree_add_51_79_groupi_n_5665);
  or csa_tree_add_51_79_groupi_g39598(csa_tree_add_51_79_groupi_n_6484 ,csa_tree_add_51_79_groupi_n_5085 ,csa_tree_add_51_79_groupi_n_5663);
  or csa_tree_add_51_79_groupi_g39599(csa_tree_add_51_79_groupi_n_6483 ,csa_tree_add_51_79_groupi_n_5087 ,csa_tree_add_51_79_groupi_n_5662);
  or csa_tree_add_51_79_groupi_g39600(csa_tree_add_51_79_groupi_n_6482 ,csa_tree_add_51_79_groupi_n_5850 ,csa_tree_add_51_79_groupi_n_5849);
  and csa_tree_add_51_79_groupi_g39601(csa_tree_add_51_79_groupi_n_6481 ,csa_tree_add_51_79_groupi_n_5850 ,csa_tree_add_51_79_groupi_n_5849);
  or csa_tree_add_51_79_groupi_g39602(csa_tree_add_51_79_groupi_n_6480 ,csa_tree_add_51_79_groupi_n_5080 ,csa_tree_add_51_79_groupi_n_5658);
  nor csa_tree_add_51_79_groupi_g39603(csa_tree_add_51_79_groupi_n_6479 ,csa_tree_add_51_79_groupi_n_5074 ,csa_tree_add_51_79_groupi_n_5657);
  or csa_tree_add_51_79_groupi_g39604(csa_tree_add_51_79_groupi_n_6478 ,csa_tree_add_51_79_groupi_n_5458 ,csa_tree_add_51_79_groupi_n_5736);
  or csa_tree_add_51_79_groupi_g39605(csa_tree_add_51_79_groupi_n_6477 ,csa_tree_add_51_79_groupi_n_5066 ,csa_tree_add_51_79_groupi_n_5650);
  nor csa_tree_add_51_79_groupi_g39606(csa_tree_add_51_79_groupi_n_6476 ,csa_tree_add_51_79_groupi_n_5058 ,csa_tree_add_51_79_groupi_n_5640);
  or csa_tree_add_51_79_groupi_g39607(csa_tree_add_51_79_groupi_n_6475 ,csa_tree_add_51_79_groupi_n_5061 ,csa_tree_add_51_79_groupi_n_5648);
  or csa_tree_add_51_79_groupi_g39608(csa_tree_add_51_79_groupi_n_6474 ,csa_tree_add_51_79_groupi_n_5057 ,csa_tree_add_51_79_groupi_n_5645);
  or csa_tree_add_51_79_groupi_g39609(csa_tree_add_51_79_groupi_n_6473 ,csa_tree_add_51_79_groupi_n_5088 ,csa_tree_add_51_79_groupi_n_5643);
  or csa_tree_add_51_79_groupi_g39610(csa_tree_add_51_79_groupi_n_6472 ,csa_tree_add_51_79_groupi_n_5052 ,csa_tree_add_51_79_groupi_n_5638);
  or csa_tree_add_51_79_groupi_g39611(csa_tree_add_51_79_groupi_n_6471 ,csa_tree_add_51_79_groupi_n_5051 ,csa_tree_add_51_79_groupi_n_5639);
  or csa_tree_add_51_79_groupi_g39612(csa_tree_add_51_79_groupi_n_6470 ,csa_tree_add_51_79_groupi_n_5049 ,csa_tree_add_51_79_groupi_n_5633);
  or csa_tree_add_51_79_groupi_g39613(csa_tree_add_51_79_groupi_n_6469 ,csa_tree_add_51_79_groupi_n_5046 ,csa_tree_add_51_79_groupi_n_5631);
  nor csa_tree_add_51_79_groupi_g39614(csa_tree_add_51_79_groupi_n_6468 ,csa_tree_add_51_79_groupi_n_5042 ,csa_tree_add_51_79_groupi_n_5623);
  or csa_tree_add_51_79_groupi_g39615(csa_tree_add_51_79_groupi_n_6467 ,csa_tree_add_51_79_groupi_n_5040 ,csa_tree_add_51_79_groupi_n_5628);
  or csa_tree_add_51_79_groupi_g39616(csa_tree_add_51_79_groupi_n_6466 ,csa_tree_add_51_79_groupi_n_5038 ,csa_tree_add_51_79_groupi_n_5626);
  or csa_tree_add_51_79_groupi_g39617(csa_tree_add_51_79_groupi_n_6465 ,csa_tree_add_51_79_groupi_n_5026 ,csa_tree_add_51_79_groupi_n_5617);
  or csa_tree_add_51_79_groupi_g39618(csa_tree_add_51_79_groupi_n_6464 ,csa_tree_add_51_79_groupi_n_5437 ,csa_tree_add_51_79_groupi_n_5624);
  nor csa_tree_add_51_79_groupi_g39619(csa_tree_add_51_79_groupi_n_6463 ,csa_tree_add_51_79_groupi_n_5445 ,csa_tree_add_51_79_groupi_n_5619);
  and csa_tree_add_51_79_groupi_g39620(csa_tree_add_51_79_groupi_n_6462 ,csa_tree_add_51_79_groupi_n_5029 ,csa_tree_add_51_79_groupi_n_5616);
  and csa_tree_add_51_79_groupi_g39621(csa_tree_add_51_79_groupi_n_6461 ,csa_tree_add_51_79_groupi_n_5027 ,csa_tree_add_51_79_groupi_n_5614);
  and csa_tree_add_51_79_groupi_g39622(csa_tree_add_51_79_groupi_n_6762 ,csa_tree_add_51_79_groupi_n_4764 ,csa_tree_add_51_79_groupi_n_5661);
  and csa_tree_add_51_79_groupi_g39623(csa_tree_add_51_79_groupi_n_6761 ,csa_tree_add_51_79_groupi_n_4759 ,csa_tree_add_51_79_groupi_n_5595);
  and csa_tree_add_51_79_groupi_g39624(csa_tree_add_51_79_groupi_n_6760 ,csa_tree_add_51_79_groupi_n_4284 ,csa_tree_add_51_79_groupi_n_5862);
  and csa_tree_add_51_79_groupi_g39625(csa_tree_add_51_79_groupi_n_6759 ,csa_tree_add_51_79_groupi_n_4778 ,csa_tree_add_51_79_groupi_n_5774);
  and csa_tree_add_51_79_groupi_g39626(csa_tree_add_51_79_groupi_n_6758 ,csa_tree_add_51_79_groupi_n_4775 ,csa_tree_add_51_79_groupi_n_5673);
  and csa_tree_add_51_79_groupi_g39627(csa_tree_add_51_79_groupi_n_6756 ,csa_tree_add_51_79_groupi_n_4080 ,csa_tree_add_51_79_groupi_n_5811);
  and csa_tree_add_51_79_groupi_g39628(csa_tree_add_51_79_groupi_n_6755 ,csa_tree_add_51_79_groupi_n_5128 ,csa_tree_add_51_79_groupi_n_5728);
  and csa_tree_add_51_79_groupi_g39629(csa_tree_add_51_79_groupi_n_6753 ,csa_tree_add_51_79_groupi_n_5136 ,csa_tree_add_51_79_groupi_n_5896);
  or csa_tree_add_51_79_groupi_g39630(csa_tree_add_51_79_groupi_n_6752 ,csa_tree_add_51_79_groupi_n_4015 ,csa_tree_add_51_79_groupi_n_5707);
  and csa_tree_add_51_79_groupi_g39631(csa_tree_add_51_79_groupi_n_6749 ,csa_tree_add_51_79_groupi_n_4402 ,csa_tree_add_51_79_groupi_n_5750);
  and csa_tree_add_51_79_groupi_g39632(csa_tree_add_51_79_groupi_n_6747 ,csa_tree_add_51_79_groupi_n_4358 ,csa_tree_add_51_79_groupi_n_5755);
  and csa_tree_add_51_79_groupi_g39633(csa_tree_add_51_79_groupi_n_6746 ,csa_tree_add_51_79_groupi_n_4316 ,csa_tree_add_51_79_groupi_n_5721);
  or csa_tree_add_51_79_groupi_g39634(csa_tree_add_51_79_groupi_n_6745 ,csa_tree_add_51_79_groupi_n_4610 ,csa_tree_add_51_79_groupi_n_6059);
  and csa_tree_add_51_79_groupi_g39635(csa_tree_add_51_79_groupi_n_6743 ,csa_tree_add_51_79_groupi_n_4131 ,csa_tree_add_51_79_groupi_n_5947);
  or csa_tree_add_51_79_groupi_g39636(csa_tree_add_51_79_groupi_n_6741 ,csa_tree_add_51_79_groupi_n_4490 ,csa_tree_add_51_79_groupi_n_6126);
  or csa_tree_add_51_79_groupi_g39637(csa_tree_add_51_79_groupi_n_6740 ,csa_tree_add_51_79_groupi_n_4550 ,csa_tree_add_51_79_groupi_n_6020);
  and csa_tree_add_51_79_groupi_g39638(csa_tree_add_51_79_groupi_n_6738 ,csa_tree_add_51_79_groupi_n_4763 ,csa_tree_add_51_79_groupi_n_5618);
  and csa_tree_add_51_79_groupi_g39639(csa_tree_add_51_79_groupi_n_6737 ,csa_tree_add_51_79_groupi_n_4756 ,csa_tree_add_51_79_groupi_n_5596);
  and csa_tree_add_51_79_groupi_g39640(csa_tree_add_51_79_groupi_n_6735 ,csa_tree_add_51_79_groupi_n_3942 ,csa_tree_add_51_79_groupi_n_5655);
  and csa_tree_add_51_79_groupi_g39641(csa_tree_add_51_79_groupi_n_6734 ,csa_tree_add_51_79_groupi_n_4760 ,csa_tree_add_51_79_groupi_n_5651);
  and csa_tree_add_51_79_groupi_g39642(csa_tree_add_51_79_groupi_n_6733 ,csa_tree_add_51_79_groupi_n_4774 ,csa_tree_add_51_79_groupi_n_5727);
  and csa_tree_add_51_79_groupi_g39643(csa_tree_add_51_79_groupi_n_6731 ,csa_tree_add_51_79_groupi_n_4766 ,csa_tree_add_51_79_groupi_n_5659);
  and csa_tree_add_51_79_groupi_g39644(csa_tree_add_51_79_groupi_n_6729 ,csa_tree_add_51_79_groupi_n_4768 ,csa_tree_add_51_79_groupi_n_5660);
  and csa_tree_add_51_79_groupi_g39645(csa_tree_add_51_79_groupi_n_6728 ,csa_tree_add_51_79_groupi_n_4060 ,csa_tree_add_51_79_groupi_n_6041);
  and csa_tree_add_51_79_groupi_g39646(csa_tree_add_51_79_groupi_n_6727 ,csa_tree_add_51_79_groupi_n_4783 ,csa_tree_add_51_79_groupi_n_5677);
  and csa_tree_add_51_79_groupi_g39647(csa_tree_add_51_79_groupi_n_6725 ,csa_tree_add_51_79_groupi_n_4770 ,csa_tree_add_51_79_groupi_n_5756);
  and csa_tree_add_51_79_groupi_g39648(csa_tree_add_51_79_groupi_n_6723 ,csa_tree_add_51_79_groupi_n_4776 ,csa_tree_add_51_79_groupi_n_5765);
  or csa_tree_add_51_79_groupi_g39649(csa_tree_add_51_79_groupi_n_6722 ,csa_tree_add_51_79_groupi_n_4076 ,csa_tree_add_51_79_groupi_n_5773);
  and csa_tree_add_51_79_groupi_g39650(csa_tree_add_51_79_groupi_n_6720 ,csa_tree_add_51_79_groupi_n_3890 ,csa_tree_add_51_79_groupi_n_5719);
  not csa_tree_add_51_79_groupi_g39652(csa_tree_add_51_79_groupi_n_6436 ,csa_tree_add_51_79_groupi_n_6437);
  not csa_tree_add_51_79_groupi_g39653(csa_tree_add_51_79_groupi_n_6429 ,csa_tree_add_51_79_groupi_n_6430);
  not csa_tree_add_51_79_groupi_g39654(csa_tree_add_51_79_groupi_n_6427 ,csa_tree_add_51_79_groupi_n_6428);
  not csa_tree_add_51_79_groupi_g39655(csa_tree_add_51_79_groupi_n_6425 ,csa_tree_add_51_79_groupi_n_6426);
  not csa_tree_add_51_79_groupi_g39656(csa_tree_add_51_79_groupi_n_6423 ,csa_tree_add_51_79_groupi_n_6424);
  not csa_tree_add_51_79_groupi_g39657(csa_tree_add_51_79_groupi_n_6421 ,csa_tree_add_51_79_groupi_n_6422);
  not csa_tree_add_51_79_groupi_g39658(csa_tree_add_51_79_groupi_n_6419 ,csa_tree_add_51_79_groupi_n_6420);
  not csa_tree_add_51_79_groupi_g39659(csa_tree_add_51_79_groupi_n_6417 ,csa_tree_add_51_79_groupi_n_6418);
  not csa_tree_add_51_79_groupi_g39660(csa_tree_add_51_79_groupi_n_6414 ,csa_tree_add_51_79_groupi_n_6415);
  not csa_tree_add_51_79_groupi_g39661(csa_tree_add_51_79_groupi_n_6411 ,csa_tree_add_51_79_groupi_n_6412);
  not csa_tree_add_51_79_groupi_g39662(csa_tree_add_51_79_groupi_n_6408 ,csa_tree_add_51_79_groupi_n_6409);
  not csa_tree_add_51_79_groupi_g39663(csa_tree_add_51_79_groupi_n_6406 ,csa_tree_add_51_79_groupi_n_6407);
  not csa_tree_add_51_79_groupi_g39664(csa_tree_add_51_79_groupi_n_6403 ,csa_tree_add_51_79_groupi_n_6404);
  not csa_tree_add_51_79_groupi_g39665(csa_tree_add_51_79_groupi_n_6401 ,csa_tree_add_51_79_groupi_n_6402);
  not csa_tree_add_51_79_groupi_g39666(csa_tree_add_51_79_groupi_n_6398 ,csa_tree_add_51_79_groupi_n_6399);
  not csa_tree_add_51_79_groupi_g39667(csa_tree_add_51_79_groupi_n_6397 ,csa_tree_add_51_79_groupi_n_6396);
  not csa_tree_add_51_79_groupi_g39668(csa_tree_add_51_79_groupi_n_6395 ,csa_tree_add_51_79_groupi_n_6394);
  xnor csa_tree_add_51_79_groupi_g39669(csa_tree_add_51_79_groupi_n_6393 ,csa_tree_add_51_79_groupi_n_4828 ,csa_tree_add_51_79_groupi_n_5474);
  xnor csa_tree_add_51_79_groupi_g39670(csa_tree_add_51_79_groupi_n_6392 ,csa_tree_add_51_79_groupi_n_5506 ,csa_tree_add_51_79_groupi_n_5367);
  xnor csa_tree_add_51_79_groupi_g39671(csa_tree_add_51_79_groupi_n_6391 ,csa_tree_add_51_79_groupi_n_5294 ,csa_tree_add_51_79_groupi_n_5483);
  xnor csa_tree_add_51_79_groupi_g39672(csa_tree_add_51_79_groupi_n_6390 ,csa_tree_add_51_79_groupi_n_3767 ,csa_tree_add_51_79_groupi_n_5565);
  xnor csa_tree_add_51_79_groupi_g39673(csa_tree_add_51_79_groupi_n_6389 ,csa_tree_add_51_79_groupi_n_3734 ,csa_tree_add_51_79_groupi_n_5100);
  xnor csa_tree_add_51_79_groupi_g39674(csa_tree_add_51_79_groupi_n_6388 ,csa_tree_add_51_79_groupi_n_3309 ,csa_tree_add_51_79_groupi_n_5423);
  xnor csa_tree_add_51_79_groupi_g39675(csa_tree_add_51_79_groupi_n_6387 ,csa_tree_add_51_79_groupi_n_3213 ,csa_tree_add_51_79_groupi_n_5059);
  xnor csa_tree_add_51_79_groupi_g39676(csa_tree_add_51_79_groupi_n_6386 ,csa_tree_add_51_79_groupi_n_5075 ,csa_tree_add_51_79_groupi_n_5216);
  xnor csa_tree_add_51_79_groupi_g39677(csa_tree_add_51_79_groupi_n_6385 ,csa_tree_add_51_79_groupi_n_5467 ,csa_tree_add_51_79_groupi_n_5242);
  xnor csa_tree_add_51_79_groupi_g39678(csa_tree_add_51_79_groupi_n_6384 ,csa_tree_add_51_79_groupi_n_4957 ,csa_tree_add_51_79_groupi_n_5029);
  xor csa_tree_add_51_79_groupi_g39679(csa_tree_add_51_79_groupi_n_6383 ,csa_tree_add_51_79_groupi_n_4847 ,csa_tree_add_51_79_groupi_n_5497);
  xnor csa_tree_add_51_79_groupi_g39680(csa_tree_add_51_79_groupi_n_6382 ,csa_tree_add_51_79_groupi_n_3241 ,csa_tree_add_51_79_groupi_n_4796);
  xnor csa_tree_add_51_79_groupi_g39681(csa_tree_add_51_79_groupi_n_6381 ,csa_tree_add_51_79_groupi_n_3279 ,csa_tree_add_51_79_groupi_n_5117);
  xnor csa_tree_add_51_79_groupi_g39682(csa_tree_add_51_79_groupi_n_6380 ,csa_tree_add_51_79_groupi_n_4819 ,csa_tree_add_51_79_groupi_n_4818);
  xnor csa_tree_add_51_79_groupi_g39683(csa_tree_add_51_79_groupi_n_6379 ,csa_tree_add_51_79_groupi_n_4826 ,csa_tree_add_51_79_groupi_n_4834);
  xnor csa_tree_add_51_79_groupi_g39684(csa_tree_add_51_79_groupi_n_6378 ,csa_tree_add_51_79_groupi_n_3773 ,csa_tree_add_51_79_groupi_n_5275);
  xnor csa_tree_add_51_79_groupi_g39685(csa_tree_add_51_79_groupi_n_6377 ,csa_tree_add_51_79_groupi_n_3235 ,csa_tree_add_51_79_groupi_n_5323);
  xnor csa_tree_add_51_79_groupi_g39686(csa_tree_add_51_79_groupi_n_6376 ,csa_tree_add_51_79_groupi_n_3785 ,csa_tree_add_51_79_groupi_n_5556);
  xnor csa_tree_add_51_79_groupi_g39687(csa_tree_add_51_79_groupi_n_6375 ,csa_tree_add_51_79_groupi_n_4969 ,csa_tree_add_51_79_groupi_n_5513);
  xnor csa_tree_add_51_79_groupi_g39688(csa_tree_add_51_79_groupi_n_6374 ,csa_tree_add_51_79_groupi_n_3752 ,csa_tree_add_51_79_groupi_n_5266);
  xnor csa_tree_add_51_79_groupi_g39689(csa_tree_add_51_79_groupi_n_6373 ,csa_tree_add_51_79_groupi_n_4832 ,csa_tree_add_51_79_groupi_n_5113);
  xnor csa_tree_add_51_79_groupi_g39690(csa_tree_add_51_79_groupi_n_6372 ,csa_tree_add_51_79_groupi_n_4809 ,csa_tree_add_51_79_groupi_n_4822);
  xnor csa_tree_add_51_79_groupi_g39691(csa_tree_add_51_79_groupi_n_6371 ,csa_tree_add_51_79_groupi_n_5119 ,csa_tree_add_51_79_groupi_n_4829);
  xnor csa_tree_add_51_79_groupi_g39692(csa_tree_add_51_79_groupi_n_6370 ,csa_tree_add_51_79_groupi_n_3799 ,csa_tree_add_51_79_groupi_n_4866);
  xnor csa_tree_add_51_79_groupi_g39693(csa_tree_add_51_79_groupi_n_6369 ,csa_tree_add_51_79_groupi_n_3272 ,csa_tree_add_51_79_groupi_n_5292);
  xnor csa_tree_add_51_79_groupi_g39694(csa_tree_add_51_79_groupi_n_6368 ,csa_tree_add_51_79_groupi_n_5397 ,csa_tree_add_51_79_groupi_n_5562);
  xnor csa_tree_add_51_79_groupi_g39695(csa_tree_add_51_79_groupi_n_6367 ,csa_tree_add_51_79_groupi_n_3806 ,csa_tree_add_51_79_groupi_n_5560);
  xnor csa_tree_add_51_79_groupi_g39696(csa_tree_add_51_79_groupi_n_6366 ,csa_tree_add_51_79_groupi_n_3238 ,csa_tree_add_51_79_groupi_n_5244);
  xnor csa_tree_add_51_79_groupi_g39697(csa_tree_add_51_79_groupi_n_6365 ,csa_tree_add_51_79_groupi_n_5262 ,csa_tree_add_51_79_groupi_n_5472);
  xnor csa_tree_add_51_79_groupi_g39698(csa_tree_add_51_79_groupi_n_6364 ,csa_tree_add_51_79_groupi_n_5347 ,csa_tree_add_51_79_groupi_n_5314);
  xnor csa_tree_add_51_79_groupi_g39699(csa_tree_add_51_79_groupi_n_6363 ,csa_tree_add_51_79_groupi_n_3304 ,csa_tree_add_51_79_groupi_n_4959);
  xnor csa_tree_add_51_79_groupi_g39700(csa_tree_add_51_79_groupi_n_6362 ,csa_tree_add_51_79_groupi_n_3286 ,csa_tree_add_51_79_groupi_n_5426);
  xnor csa_tree_add_51_79_groupi_g39701(csa_tree_add_51_79_groupi_n_6361 ,csa_tree_add_51_79_groupi_n_4887 ,csa_tree_add_51_79_groupi_n_5074);
  xnor csa_tree_add_51_79_groupi_g39702(csa_tree_add_51_79_groupi_n_6360 ,csa_tree_add_51_79_groupi_n_4837 ,csa_tree_add_51_79_groupi_n_5538);
  xnor csa_tree_add_51_79_groupi_g39703(csa_tree_add_51_79_groupi_n_6359 ,csa_tree_add_51_79_groupi_n_5496 ,csa_tree_add_51_79_groupi_n_5360);
  xnor csa_tree_add_51_79_groupi_g39704(csa_tree_add_51_79_groupi_n_6358 ,csa_tree_add_51_79_groupi_n_3825 ,csa_tree_add_51_79_groupi_n_5511);
  xnor csa_tree_add_51_79_groupi_g39705(csa_tree_add_51_79_groupi_n_6357 ,csa_tree_add_51_79_groupi_n_3821 ,csa_tree_add_51_79_groupi_n_5337);
  xnor csa_tree_add_51_79_groupi_g39706(csa_tree_add_51_79_groupi_n_6356 ,csa_tree_add_51_79_groupi_n_5310 ,csa_tree_add_51_79_groupi_n_5264);
  xnor csa_tree_add_51_79_groupi_g39707(csa_tree_add_51_79_groupi_n_6355 ,csa_tree_add_51_79_groupi_n_3789 ,csa_tree_add_51_79_groupi_n_5300);
  xnor csa_tree_add_51_79_groupi_g39708(csa_tree_add_51_79_groupi_n_6354 ,csa_tree_add_51_79_groupi_n_5567 ,csa_tree_add_51_79_groupi_n_5321);
  xnor csa_tree_add_51_79_groupi_g39709(csa_tree_add_51_79_groupi_n_6353 ,csa_tree_add_51_79_groupi_n_4892 ,csa_tree_add_51_79_groupi_n_5303);
  xnor csa_tree_add_51_79_groupi_g39710(csa_tree_add_51_79_groupi_n_6352 ,csa_tree_add_51_79_groupi_n_3771 ,csa_tree_add_51_79_groupi_n_5241);
  xnor csa_tree_add_51_79_groupi_g39711(csa_tree_add_51_79_groupi_n_6351 ,csa_tree_add_51_79_groupi_n_3292 ,csa_tree_add_51_79_groupi_n_5080);
  xnor csa_tree_add_51_79_groupi_g39712(csa_tree_add_51_79_groupi_n_6350 ,csa_tree_add_51_79_groupi_n_3215 ,csa_tree_add_51_79_groupi_n_5403);
  xnor csa_tree_add_51_79_groupi_g39713(csa_tree_add_51_79_groupi_n_6349 ,csa_tree_add_51_79_groupi_n_5419 ,csa_tree_add_51_79_groupi_n_4859);
  xnor csa_tree_add_51_79_groupi_g39714(csa_tree_add_51_79_groupi_n_6348 ,csa_tree_add_51_79_groupi_n_5333 ,csa_tree_add_51_79_groupi_n_4900);
  xnor csa_tree_add_51_79_groupi_g39715(csa_tree_add_51_79_groupi_n_6347 ,csa_tree_add_51_79_groupi_n_5524 ,csa_tree_add_51_79_groupi_n_4799);
  xnor csa_tree_add_51_79_groupi_g39716(csa_tree_add_51_79_groupi_n_6346 ,csa_tree_add_51_79_groupi_n_5199 ,csa_tree_add_51_79_groupi_n_5184);
  xnor csa_tree_add_51_79_groupi_g39717(csa_tree_add_51_79_groupi_n_6345 ,csa_tree_add_51_79_groupi_n_4941 ,csa_tree_add_51_79_groupi_n_5445);
  xnor csa_tree_add_51_79_groupi_g39718(csa_tree_add_51_79_groupi_n_6344 ,csa_tree_add_51_79_groupi_n_3746 ,csa_tree_add_51_79_groupi_n_5062);
  xnor csa_tree_add_51_79_groupi_g39719(csa_tree_add_51_79_groupi_n_6343 ,csa_tree_add_51_79_groupi_n_5271 ,csa_tree_add_51_79_groupi_n_5532);
  xnor csa_tree_add_51_79_groupi_g39720(csa_tree_add_51_79_groupi_n_6342 ,csa_tree_add_51_79_groupi_n_5364 ,csa_tree_add_51_79_groupi_n_5573);
  xnor csa_tree_add_51_79_groupi_g39721(csa_tree_add_51_79_groupi_n_6341 ,csa_tree_add_51_79_groupi_n_3284 ,csa_tree_add_51_79_groupi_n_5441);
  xnor csa_tree_add_51_79_groupi_g39722(csa_tree_add_51_79_groupi_n_6340 ,csa_tree_add_51_79_groupi_n_3760 ,csa_tree_add_51_79_groupi_n_5484);
  xnor csa_tree_add_51_79_groupi_g39723(csa_tree_add_51_79_groupi_n_6339 ,csa_tree_add_51_79_groupi_n_5219 ,csa_tree_add_51_79_groupi_n_5220);
  xnor csa_tree_add_51_79_groupi_g39724(csa_tree_add_51_79_groupi_n_6338 ,csa_tree_add_51_79_groupi_n_3296 ,csa_tree_add_51_79_groupi_n_5237);
  xnor csa_tree_add_51_79_groupi_g39725(csa_tree_add_51_79_groupi_n_6337 ,csa_tree_add_51_79_groupi_n_3803 ,csa_tree_add_51_79_groupi_n_5160);
  xnor csa_tree_add_51_79_groupi_g39726(csa_tree_add_51_79_groupi_n_6336 ,csa_tree_add_51_79_groupi_n_3302 ,csa_tree_add_51_79_groupi_n_5455);
  xnor csa_tree_add_51_79_groupi_g39727(csa_tree_add_51_79_groupi_n_6335 ,csa_tree_add_51_79_groupi_n_5187 ,csa_tree_add_51_79_groupi_n_4813);
  xnor csa_tree_add_51_79_groupi_g39728(csa_tree_add_51_79_groupi_n_6334 ,csa_tree_add_51_79_groupi_n_5222 ,csa_tree_add_51_79_groupi_n_5223);
  xnor csa_tree_add_51_79_groupi_g39729(csa_tree_add_51_79_groupi_n_6333 ,csa_tree_add_51_79_groupi_n_5561 ,csa_tree_add_51_79_groupi_n_5376);
  xnor csa_tree_add_51_79_groupi_g39730(csa_tree_add_51_79_groupi_n_6332 ,csa_tree_add_51_79_groupi_n_4964 ,csa_tree_add_51_79_groupi_n_5478);
  xnor csa_tree_add_51_79_groupi_g39731(csa_tree_add_51_79_groupi_n_6331 ,csa_tree_add_51_79_groupi_n_3819 ,csa_tree_add_51_79_groupi_n_4932);
  xnor csa_tree_add_51_79_groupi_g39732(csa_tree_add_51_79_groupi_n_6330 ,csa_tree_add_51_79_groupi_n_5022 ,csa_tree_add_51_79_groupi_n_5370);
  xnor csa_tree_add_51_79_groupi_g39733(csa_tree_add_51_79_groupi_n_6329 ,csa_tree_add_51_79_groupi_n_4989 ,csa_tree_add_51_79_groupi_n_4840);
  xnor csa_tree_add_51_79_groupi_g39734(csa_tree_add_51_79_groupi_n_6328 ,csa_tree_add_51_79_groupi_n_5063 ,csa_tree_add_51_79_groupi_n_5326);
  xnor csa_tree_add_51_79_groupi_g39735(csa_tree_add_51_79_groupi_n_6327 ,csa_tree_add_51_79_groupi_n_5033 ,csa_tree_add_51_79_groupi_n_5255);
  xnor csa_tree_add_51_79_groupi_g39736(csa_tree_add_51_79_groupi_n_6326 ,csa_tree_add_51_79_groupi_n_4908 ,csa_tree_add_51_79_groupi_n_765);
  xnor csa_tree_add_51_79_groupi_g39737(csa_tree_add_51_79_groupi_n_6325 ,csa_tree_add_51_79_groupi_n_5393 ,csa_tree_add_51_79_groupi_n_5182);
  xnor csa_tree_add_51_79_groupi_g39738(csa_tree_add_51_79_groupi_n_6324 ,csa_tree_add_51_79_groupi_n_5193 ,csa_tree_add_51_79_groupi_n_5519);
  xnor csa_tree_add_51_79_groupi_g39739(csa_tree_add_51_79_groupi_n_6323 ,csa_tree_add_51_79_groupi_n_5044 ,csa_tree_add_51_79_groupi_n_5204);
  xnor csa_tree_add_51_79_groupi_g39740(csa_tree_add_51_79_groupi_n_6322 ,csa_tree_add_51_79_groupi_n_4808 ,csa_tree_add_51_79_groupi_n_4970);
  xnor csa_tree_add_51_79_groupi_g39741(csa_tree_add_51_79_groupi_n_6321 ,csa_tree_add_51_79_groupi_n_5156 ,csa_tree_add_51_79_groupi_n_4980);
  xnor csa_tree_add_51_79_groupi_g39742(csa_tree_add_51_79_groupi_n_6320 ,csa_tree_add_51_79_groupi_n_5124 ,csa_tree_add_51_79_groupi_n_4894);
  xnor csa_tree_add_51_79_groupi_g39743(csa_tree_add_51_79_groupi_n_6319 ,csa_tree_add_51_79_groupi_n_5383 ,csa_tree_add_51_79_groupi_n_4984);
  xnor csa_tree_add_51_79_groupi_g39744(csa_tree_add_51_79_groupi_n_6318 ,csa_tree_add_51_79_groupi_n_4850 ,csa_tree_add_51_79_groupi_n_4889);
  xnor csa_tree_add_51_79_groupi_g39745(csa_tree_add_51_79_groupi_n_6317 ,csa_tree_add_51_79_groupi_n_4877 ,csa_tree_add_51_79_groupi_n_4987);
  xnor csa_tree_add_51_79_groupi_g39746(csa_tree_add_51_79_groupi_n_6316 ,csa_tree_add_51_79_groupi_n_5026 ,csa_tree_add_51_79_groupi_n_4882);
  xnor csa_tree_add_51_79_groupi_g39747(csa_tree_add_51_79_groupi_n_6315 ,csa_tree_add_51_79_groupi_n_5114 ,csa_tree_add_51_79_groupi_n_4890);
  xnor csa_tree_add_51_79_groupi_g39748(csa_tree_add_51_79_groupi_n_6314 ,csa_tree_add_51_79_groupi_n_4927 ,csa_tree_add_51_79_groupi_n_4929);
  xnor csa_tree_add_51_79_groupi_g39749(csa_tree_add_51_79_groupi_n_6313 ,csa_tree_add_51_79_groupi_n_5427 ,csa_tree_add_51_79_groupi_n_5006);
  xnor csa_tree_add_51_79_groupi_g39750(csa_tree_add_51_79_groupi_n_6312 ,csa_tree_add_51_79_groupi_n_5424 ,csa_tree_add_51_79_groupi_n_4906);
  xnor csa_tree_add_51_79_groupi_g39751(csa_tree_add_51_79_groupi_n_6311 ,csa_tree_add_51_79_groupi_n_5421 ,csa_tree_add_51_79_groupi_n_5008);
  xnor csa_tree_add_51_79_groupi_g39752(csa_tree_add_51_79_groupi_n_6310 ,csa_tree_add_51_79_groupi_n_5269 ,csa_tree_add_51_79_groupi_n_4991);
  xnor csa_tree_add_51_79_groupi_g39753(csa_tree_add_51_79_groupi_n_6309 ,csa_tree_add_51_79_groupi_n_5247 ,csa_tree_add_51_79_groupi_n_4953);
  xnor csa_tree_add_51_79_groupi_g39754(csa_tree_add_51_79_groupi_n_6308 ,csa_tree_add_51_79_groupi_n_5263 ,csa_tree_add_51_79_groupi_n_4999);
  xnor csa_tree_add_51_79_groupi_g39755(csa_tree_add_51_79_groupi_n_6307 ,csa_tree_add_51_79_groupi_n_5186 ,csa_tree_add_51_79_groupi_n_4948);
  xnor csa_tree_add_51_79_groupi_g39756(csa_tree_add_51_79_groupi_n_6306 ,csa_tree_add_51_79_groupi_n_5318 ,csa_tree_add_51_79_groupi_n_4881);
  xnor csa_tree_add_51_79_groupi_g39757(csa_tree_add_51_79_groupi_n_6305 ,csa_tree_add_51_79_groupi_n_5428 ,csa_tree_add_51_79_groupi_n_4997);
  xnor csa_tree_add_51_79_groupi_g39758(csa_tree_add_51_79_groupi_n_6304 ,csa_tree_add_51_79_groupi_n_5196 ,csa_tree_add_51_79_groupi_n_4996);
  xnor csa_tree_add_51_79_groupi_g39759(csa_tree_add_51_79_groupi_n_6303 ,csa_tree_add_51_79_groupi_n_5167 ,csa_tree_add_51_79_groupi_n_5003);
  xnor csa_tree_add_51_79_groupi_g39760(csa_tree_add_51_79_groupi_n_6302 ,csa_tree_add_51_79_groupi_n_4812 ,csa_tree_add_51_79_groupi_n_4919);
  xnor csa_tree_add_51_79_groupi_g39761(csa_tree_add_51_79_groupi_n_6301 ,csa_tree_add_51_79_groupi_n_5248 ,csa_tree_add_51_79_groupi_n_5000);
  xnor csa_tree_add_51_79_groupi_g39762(csa_tree_add_51_79_groupi_n_6300 ,csa_tree_add_51_79_groupi_n_5157 ,csa_tree_add_51_79_groupi_n_4995);
  xnor csa_tree_add_51_79_groupi_g39763(csa_tree_add_51_79_groupi_n_6299 ,csa_tree_add_51_79_groupi_n_5414 ,csa_tree_add_51_79_groupi_n_5007);
  xnor csa_tree_add_51_79_groupi_g39764(csa_tree_add_51_79_groupi_n_6298 ,csa_tree_add_51_79_groupi_n_5161 ,csa_tree_add_51_79_groupi_n_4986);
  xnor csa_tree_add_51_79_groupi_g39765(csa_tree_add_51_79_groupi_n_6297 ,csa_tree_add_51_79_groupi_n_5176 ,csa_tree_add_51_79_groupi_n_4993);
  xnor csa_tree_add_51_79_groupi_g39766(csa_tree_add_51_79_groupi_n_6296 ,csa_tree_add_51_79_groupi_n_4933 ,csa_tree_add_51_79_groupi_n_4934);
  xnor csa_tree_add_51_79_groupi_g39767(csa_tree_add_51_79_groupi_n_6295 ,csa_tree_add_51_79_groupi_n_5202 ,csa_tree_add_51_79_groupi_n_4998);
  xnor csa_tree_add_51_79_groupi_g39768(csa_tree_add_51_79_groupi_n_6294 ,csa_tree_add_51_79_groupi_n_5249 ,csa_tree_add_51_79_groupi_n_4905);
  xnor csa_tree_add_51_79_groupi_g39769(csa_tree_add_51_79_groupi_n_6293 ,csa_tree_add_51_79_groupi_n_5190 ,csa_tree_add_51_79_groupi_n_5002);
  xnor csa_tree_add_51_79_groupi_g39770(csa_tree_add_51_79_groupi_n_6292 ,csa_tree_add_51_79_groupi_n_5171 ,csa_tree_add_51_79_groupi_n_4903);
  xnor csa_tree_add_51_79_groupi_g39771(csa_tree_add_51_79_groupi_n_6291 ,csa_tree_add_51_79_groupi_n_5379 ,csa_tree_add_51_79_groupi_n_4983);
  xnor csa_tree_add_51_79_groupi_g39772(csa_tree_add_51_79_groupi_n_6290 ,csa_tree_add_51_79_groupi_n_5353 ,csa_tree_add_51_79_groupi_n_4901);
  xnor csa_tree_add_51_79_groupi_g39773(csa_tree_add_51_79_groupi_n_6289 ,csa_tree_add_51_79_groupi_n_5330 ,csa_tree_add_51_79_groupi_n_4975);
  xnor csa_tree_add_51_79_groupi_g39774(csa_tree_add_51_79_groupi_n_6288 ,csa_tree_add_51_79_groupi_n_5165 ,csa_tree_add_51_79_groupi_n_4972);
  xnor csa_tree_add_51_79_groupi_g39775(csa_tree_add_51_79_groupi_n_6287 ,csa_tree_add_51_79_groupi_n_5311 ,csa_tree_add_51_79_groupi_n_4971);
  xnor csa_tree_add_51_79_groupi_g39776(csa_tree_add_51_79_groupi_n_6286 ,csa_tree_add_51_79_groupi_n_5420 ,csa_tree_add_51_79_groupi_n_4944);
  xnor csa_tree_add_51_79_groupi_g39777(csa_tree_add_51_79_groupi_n_6285 ,csa_tree_add_51_79_groupi_n_5057 ,csa_tree_add_51_79_groupi_n_4885);
  xnor csa_tree_add_51_79_groupi_g39778(csa_tree_add_51_79_groupi_n_6284 ,csa_tree_add_51_79_groupi_n_5365 ,csa_tree_add_51_79_groupi_n_4979);
  xnor csa_tree_add_51_79_groupi_g39779(csa_tree_add_51_79_groupi_n_6283 ,csa_tree_add_51_79_groupi_n_5203 ,csa_tree_add_51_79_groupi_n_4992);
  xnor csa_tree_add_51_79_groupi_g39780(csa_tree_add_51_79_groupi_n_6282 ,csa_tree_add_51_79_groupi_n_5239 ,csa_tree_add_51_79_groupi_n_4955);
  xnor csa_tree_add_51_79_groupi_g39781(csa_tree_add_51_79_groupi_n_6281 ,csa_tree_add_51_79_groupi_n_5261 ,csa_tree_add_51_79_groupi_n_4960);
  xnor csa_tree_add_51_79_groupi_g39782(csa_tree_add_51_79_groupi_n_6280 ,csa_tree_add_51_79_groupi_n_4926 ,csa_tree_add_51_79_groupi_n_4884);
  xnor csa_tree_add_51_79_groupi_g39783(csa_tree_add_51_79_groupi_n_6279 ,csa_tree_add_51_79_groupi_n_5246 ,csa_tree_add_51_79_groupi_n_4917);
  xnor csa_tree_add_51_79_groupi_g39784(csa_tree_add_51_79_groupi_n_6278 ,csa_tree_add_51_79_groupi_n_5290 ,csa_tree_add_51_79_groupi_n_4965);
  xnor csa_tree_add_51_79_groupi_g39785(csa_tree_add_51_79_groupi_n_6277 ,csa_tree_add_51_79_groupi_n_4848 ,csa_tree_add_51_79_groupi_n_4893);
  xnor csa_tree_add_51_79_groupi_g39786(csa_tree_add_51_79_groupi_n_6276 ,csa_tree_add_51_79_groupi_n_5312 ,csa_tree_add_51_79_groupi_n_5001);
  xnor csa_tree_add_51_79_groupi_g39787(csa_tree_add_51_79_groupi_n_6275 ,csa_tree_add_51_79_groupi_n_4897 ,csa_tree_add_51_79_groupi_n_3232);
  xnor csa_tree_add_51_79_groupi_g39788(csa_tree_add_51_79_groupi_n_6274 ,csa_tree_add_51_79_groupi_n_5412 ,csa_tree_add_51_79_groupi_n_4938);
  xnor csa_tree_add_51_79_groupi_g39789(csa_tree_add_51_79_groupi_n_6273 ,csa_tree_add_51_79_groupi_n_5180 ,csa_tree_add_51_79_groupi_n_4981);
  xnor csa_tree_add_51_79_groupi_g39790(csa_tree_add_51_79_groupi_n_6272 ,csa_tree_add_51_79_groupi_n_5212 ,csa_tree_add_51_79_groupi_n_4947);
  xnor csa_tree_add_51_79_groupi_g39791(csa_tree_add_51_79_groupi_n_6271 ,csa_tree_add_51_79_groupi_n_5209 ,csa_tree_add_51_79_groupi_n_4918);
  xnor csa_tree_add_51_79_groupi_g39792(csa_tree_add_51_79_groupi_n_6270 ,csa_tree_add_51_79_groupi_n_5177 ,csa_tree_add_51_79_groupi_n_4937);
  xnor csa_tree_add_51_79_groupi_g39793(csa_tree_add_51_79_groupi_n_6269 ,csa_tree_add_51_79_groupi_n_5173 ,csa_tree_add_51_79_groupi_n_4902);
  xnor csa_tree_add_51_79_groupi_g39794(csa_tree_add_51_79_groupi_n_6268 ,csa_tree_add_51_79_groupi_n_5158 ,csa_tree_add_51_79_groupi_n_4990);
  xnor csa_tree_add_51_79_groupi_g39795(csa_tree_add_51_79_groupi_n_6267 ,csa_tree_add_51_79_groupi_n_5169 ,csa_tree_add_51_79_groupi_n_4940);
  xnor csa_tree_add_51_79_groupi_g39796(csa_tree_add_51_79_groupi_n_6266 ,csa_tree_add_51_79_groupi_n_5192 ,csa_tree_add_51_79_groupi_n_4916);
  xnor csa_tree_add_51_79_groupi_g39797(csa_tree_add_51_79_groupi_n_6265 ,csa_tree_add_51_79_groupi_n_4802 ,csa_tree_add_51_79_groupi_n_4994);
  xnor csa_tree_add_51_79_groupi_g39798(csa_tree_add_51_79_groupi_n_6264 ,csa_tree_add_51_79_groupi_n_4924 ,csa_tree_add_51_79_groupi_n_4925);
  xnor csa_tree_add_51_79_groupi_g39799(csa_tree_add_51_79_groupi_n_6263 ,csa_tree_add_51_79_groupi_n_5005 ,csa_tree_add_51_79_groupi_n_4915);
  xnor csa_tree_add_51_79_groupi_g39800(csa_tree_add_51_79_groupi_n_6262 ,csa_tree_add_51_79_groupi_n_4907 ,csa_tree_add_51_79_groupi_n_4982);
  xnor csa_tree_add_51_79_groupi_g39801(csa_tree_add_51_79_groupi_n_6261 ,csa_tree_add_51_79_groupi_n_4913 ,csa_tree_add_51_79_groupi_n_4899);
  xnor csa_tree_add_51_79_groupi_g39802(csa_tree_add_51_79_groupi_n_6260 ,csa_tree_add_51_79_groupi_n_5226 ,csa_tree_add_51_79_groupi_n_4952);
  xnor csa_tree_add_51_79_groupi_g39803(csa_tree_add_51_79_groupi_n_6259 ,csa_tree_add_51_79_groupi_n_5009 ,csa_tree_add_51_79_groupi_n_4911);
  xnor csa_tree_add_51_79_groupi_g39804(csa_tree_add_51_79_groupi_n_6258 ,csa_tree_add_51_79_groupi_n_5164 ,csa_tree_add_51_79_groupi_n_5045);
  xnor csa_tree_add_51_79_groupi_g39805(csa_tree_add_51_79_groupi_n_6257 ,csa_tree_add_51_79_groupi_n_5105 ,csa_tree_add_51_79_groupi_n_4935);
  xnor csa_tree_add_51_79_groupi_g39806(csa_tree_add_51_79_groupi_n_6256 ,csa_tree_add_51_79_groupi_n_5101 ,csa_tree_add_51_79_groupi_n_4974);
  xnor csa_tree_add_51_79_groupi_g39807(csa_tree_add_51_79_groupi_n_6255 ,csa_tree_add_51_79_groupi_n_4798 ,csa_tree_add_51_79_groupi_n_5055);
  xnor csa_tree_add_51_79_groupi_g39808(csa_tree_add_51_79_groupi_n_6254 ,csa_tree_add_51_79_groupi_n_5170 ,csa_tree_add_51_79_groupi_n_5071);
  xnor csa_tree_add_51_79_groupi_g39809(csa_tree_add_51_79_groupi_n_6253 ,csa_tree_add_51_79_groupi_n_5108 ,csa_tree_add_51_79_groupi_n_4985);
  xnor csa_tree_add_51_79_groupi_g39810(csa_tree_add_51_79_groupi_n_6252 ,csa_tree_add_51_79_groupi_n_5523 ,csa_tree_add_51_79_groupi_n_4898);
  xor csa_tree_add_51_79_groupi_g39811(csa_tree_add_51_79_groupi_n_6251 ,csa_tree_add_51_79_groupi_n_3204 ,csa_tree_add_51_79_groupi_n_5058);
  xnor csa_tree_add_51_79_groupi_g39812(csa_tree_add_51_79_groupi_n_6250 ,csa_tree_add_51_79_groupi_n_5357 ,csa_tree_add_51_79_groupi_n_4853);
  xnor csa_tree_add_51_79_groupi_g39813(csa_tree_add_51_79_groupi_n_6249 ,csa_tree_add_51_79_groupi_n_5429 ,csa_tree_add_51_79_groupi_n_5433);
  xnor csa_tree_add_51_79_groupi_g39814(csa_tree_add_51_79_groupi_n_6248 ,csa_tree_add_51_79_groupi_n_5566 ,csa_tree_add_51_79_groupi_n_5341);
  xnor csa_tree_add_51_79_groupi_g39815(csa_tree_add_51_79_groupi_n_6247 ,csa_tree_add_51_79_groupi_n_5276 ,csa_tree_add_51_79_groupi_n_5277);
  xnor csa_tree_add_51_79_groupi_g39816(csa_tree_add_51_79_groupi_n_6246 ,csa_tree_add_51_79_groupi_n_5218 ,csa_tree_add_51_79_groupi_n_5197);
  xnor csa_tree_add_51_79_groupi_g39817(csa_tree_add_51_79_groupi_n_6245 ,csa_tree_add_51_79_groupi_n_5557 ,csa_tree_add_51_79_groupi_n_5345);
  xor csa_tree_add_51_79_groupi_g39818(csa_tree_add_51_79_groupi_n_6244 ,csa_tree_add_51_79_groupi_n_3290 ,csa_tree_add_51_79_groupi_n_5451);
  xnor csa_tree_add_51_79_groupi_g39819(csa_tree_add_51_79_groupi_n_6243 ,csa_tree_add_51_79_groupi_n_5498 ,csa_tree_add_51_79_groupi_n_5343);
  xnor csa_tree_add_51_79_groupi_g39820(csa_tree_add_51_79_groupi_n_6242 ,csa_tree_add_51_79_groupi_n_5225 ,csa_tree_add_51_79_groupi_n_5227);
  xnor csa_tree_add_51_79_groupi_g39821(csa_tree_add_51_79_groupi_n_6241 ,csa_tree_add_51_79_groupi_n_4852 ,csa_tree_add_51_79_groupi_n_5356);
  xnor csa_tree_add_51_79_groupi_g39822(csa_tree_add_51_79_groupi_n_6240 ,csa_tree_add_51_79_groupi_n_5245 ,csa_tree_add_51_79_groupi_n_5575);
  xnor csa_tree_add_51_79_groupi_g39823(csa_tree_add_51_79_groupi_n_6239 ,csa_tree_add_51_79_groupi_n_5260 ,csa_tree_add_51_79_groupi_n_5515);
  xnor csa_tree_add_51_79_groupi_g39824(csa_tree_add_51_79_groupi_n_6238 ,csa_tree_add_51_79_groupi_n_5378 ,csa_tree_add_51_79_groupi_n_5382);
  xor csa_tree_add_51_79_groupi_g39825(csa_tree_add_51_79_groupi_n_6237 ,csa_tree_add_51_79_groupi_n_5362 ,csa_tree_add_51_79_groupi_n_5577);
  xnor csa_tree_add_51_79_groupi_g39826(csa_tree_add_51_79_groupi_n_6236 ,csa_tree_add_51_79_groupi_n_5230 ,csa_tree_add_51_79_groupi_n_5233);
  xnor csa_tree_add_51_79_groupi_g39827(csa_tree_add_51_79_groupi_n_6235 ,csa_tree_add_51_79_groupi_n_5447 ,csa_tree_add_51_79_groupi_n_5287);
  xor csa_tree_add_51_79_groupi_g39828(csa_tree_add_51_79_groupi_n_6234 ,csa_tree_add_51_79_groupi_n_5163 ,csa_tree_add_51_79_groupi_n_5461);
  xnor csa_tree_add_51_79_groupi_g39829(csa_tree_add_51_79_groupi_n_6233 ,csa_tree_add_51_79_groupi_n_5253 ,csa_tree_add_51_79_groupi_n_5256);
  xnor csa_tree_add_51_79_groupi_g39830(csa_tree_add_51_79_groupi_n_6232 ,csa_tree_add_51_79_groupi_n_5284 ,csa_tree_add_51_79_groupi_n_5285);
  xnor csa_tree_add_51_79_groupi_g39831(csa_tree_add_51_79_groupi_n_6231 ,csa_tree_add_51_79_groupi_n_5510 ,csa_tree_add_51_79_groupi_n_4895);
  xnor csa_tree_add_51_79_groupi_g39832(csa_tree_add_51_79_groupi_n_6230 ,csa_tree_add_51_79_groupi_n_5501 ,csa_tree_add_51_79_groupi_n_4797);
  xor csa_tree_add_51_79_groupi_g39833(csa_tree_add_51_79_groupi_n_6229 ,csa_tree_add_51_79_groupi_n_3280 ,csa_tree_add_51_79_groupi_n_5042);
  xnor csa_tree_add_51_79_groupi_g39834(csa_tree_add_51_79_groupi_n_6228 ,csa_tree_add_51_79_groupi_n_4810 ,csa_tree_add_51_79_groupi_n_5122);
  xnor csa_tree_add_51_79_groupi_g39835(csa_tree_add_51_79_groupi_n_6227 ,csa_tree_add_51_79_groupi_n_4836 ,csa_tree_add_51_79_groupi_n_5448);
  xnor csa_tree_add_51_79_groupi_g39836(csa_tree_add_51_79_groupi_n_6226 ,csa_tree_add_51_79_groupi_n_4816 ,csa_tree_add_51_79_groupi_n_5487);
  xnor csa_tree_add_51_79_groupi_g39837(csa_tree_add_51_79_groupi_n_6225 ,csa_tree_add_51_79_groupi_n_5297 ,csa_tree_add_51_79_groupi_n_5516);
  xnor csa_tree_add_51_79_groupi_g39838(csa_tree_add_51_79_groupi_n_6224 ,csa_tree_add_51_79_groupi_n_5494 ,csa_tree_add_51_79_groupi_n_5211);
  xnor csa_tree_add_51_79_groupi_g39839(csa_tree_add_51_79_groupi_n_6223 ,csa_tree_add_51_79_groupi_n_4914 ,csa_tree_add_51_79_groupi_n_5061);
  xnor csa_tree_add_51_79_groupi_g39840(csa_tree_add_51_79_groupi_n_6222 ,csa_tree_add_51_79_groupi_n_4910 ,csa_tree_add_51_79_groupi_n_4909);
  xnor csa_tree_add_51_79_groupi_g39841(csa_tree_add_51_79_groupi_n_6221 ,csa_tree_add_51_79_groupi_n_4977 ,csa_tree_add_51_79_groupi_n_5508);
  xnor csa_tree_add_51_79_groupi_g39842(csa_tree_add_51_79_groupi_n_6220 ,csa_tree_add_51_79_groupi_n_5338 ,csa_tree_add_51_79_groupi_n_5096);
  xor csa_tree_add_51_79_groupi_g39843(csa_tree_add_51_79_groupi_n_6219 ,csa_tree_add_51_79_groupi_n_3264 ,csa_tree_add_51_79_groupi_n_5446);
  xnor csa_tree_add_51_79_groupi_g39844(csa_tree_add_51_79_groupi_n_6218 ,csa_tree_add_51_79_groupi_n_4923 ,csa_tree_add_51_79_groupi_n_3260);
  xnor csa_tree_add_51_79_groupi_g39845(csa_tree_add_51_79_groupi_n_6217 ,csa_tree_add_51_79_groupi_n_5201 ,csa_tree_add_51_79_groupi_n_5531);
  xnor csa_tree_add_51_79_groupi_g39846(csa_tree_add_51_79_groupi_n_6216 ,csa_tree_add_51_79_groupi_n_4879 ,csa_tree_add_51_79_groupi_n_5085);
  xnor csa_tree_add_51_79_groupi_g39847(csa_tree_add_51_79_groupi_n_6215 ,csa_tree_add_51_79_groupi_n_4851 ,csa_tree_add_51_79_groupi_n_5293);
  xnor csa_tree_add_51_79_groupi_g39848(csa_tree_add_51_79_groupi_n_6214 ,csa_tree_add_51_79_groupi_n_5094 ,csa_tree_add_51_79_groupi_n_4870);
  xnor csa_tree_add_51_79_groupi_g39849(csa_tree_add_51_79_groupi_n_6213 ,csa_tree_add_51_79_groupi_n_4868 ,csa_tree_add_51_79_groupi_n_4867);
  xnor csa_tree_add_51_79_groupi_g39850(csa_tree_add_51_79_groupi_n_6212 ,csa_tree_add_51_79_groupi_n_4876 ,csa_tree_add_51_79_groupi_n_5095);
  xnor csa_tree_add_51_79_groupi_g39851(csa_tree_add_51_79_groupi_n_6211 ,csa_tree_add_51_79_groupi_n_5038 ,csa_tree_add_51_79_groupi_n_5010);
  xnor csa_tree_add_51_79_groupi_g39852(csa_tree_add_51_79_groupi_n_6210 ,csa_tree_add_51_79_groupi_n_4943 ,csa_tree_add_51_79_groupi_n_5040);
  xnor csa_tree_add_51_79_groupi_g39853(csa_tree_add_51_79_groupi_n_6209 ,csa_tree_add_51_79_groupi_n_4872 ,csa_tree_add_51_79_groupi_n_5099);
  xnor csa_tree_add_51_79_groupi_g39854(csa_tree_add_51_79_groupi_n_6208 ,csa_tree_add_51_79_groupi_n_5051 ,csa_tree_add_51_79_groupi_n_4928);
  xnor csa_tree_add_51_79_groupi_g39855(csa_tree_add_51_79_groupi_n_6207 ,csa_tree_add_51_79_groupi_n_4883 ,csa_tree_add_51_79_groupi_n_4880);
  xnor csa_tree_add_51_79_groupi_g39856(csa_tree_add_51_79_groupi_n_6206 ,csa_tree_add_51_79_groupi_n_4888 ,csa_tree_add_51_79_groupi_n_4886);
  xnor csa_tree_add_51_79_groupi_g39857(csa_tree_add_51_79_groupi_n_6205 ,csa_tree_add_51_79_groupi_n_5437 ,csa_tree_add_51_79_groupi_n_4951);
  xnor csa_tree_add_51_79_groupi_g39858(csa_tree_add_51_79_groupi_n_6204 ,csa_tree_add_51_79_groupi_n_5399 ,csa_tree_add_51_79_groupi_n_5525);
  xnor csa_tree_add_51_79_groupi_g39859(csa_tree_add_51_79_groupi_n_6203 ,csa_tree_add_51_79_groupi_n_5304 ,csa_tree_add_51_79_groupi_n_5485);
  xnor csa_tree_add_51_79_groupi_g39860(csa_tree_add_51_79_groupi_n_6202 ,csa_tree_add_51_79_groupi_n_5495 ,csa_tree_add_51_79_groupi_n_5332);
  xnor csa_tree_add_51_79_groupi_g39861(csa_tree_add_51_79_groupi_n_6201 ,csa_tree_add_51_79_groupi_n_5121 ,csa_tree_add_51_79_groupi_n_4824);
  xnor csa_tree_add_51_79_groupi_g39862(csa_tree_add_51_79_groupi_n_6200 ,csa_tree_add_51_79_groupi_n_4838 ,csa_tree_add_51_79_groupi_n_5404);
  xnor csa_tree_add_51_79_groupi_g39863(csa_tree_add_51_79_groupi_n_6199 ,csa_tree_add_51_79_groupi_n_5320 ,csa_tree_add_51_79_groupi_n_5392);
  xnor csa_tree_add_51_79_groupi_g39864(csa_tree_add_51_79_groupi_n_6198 ,csa_tree_add_51_79_groupi_n_5391 ,csa_tree_add_51_79_groupi_n_5405);
  xnor csa_tree_add_51_79_groupi_g39865(csa_tree_add_51_79_groupi_n_6197 ,csa_tree_add_51_79_groupi_n_5390 ,csa_tree_add_51_79_groupi_n_3748);
  xnor csa_tree_add_51_79_groupi_g39866(csa_tree_add_51_79_groupi_n_6196 ,csa_tree_add_51_79_groupi_n_5340 ,csa_tree_add_51_79_groupi_n_5339);
  xnor csa_tree_add_51_79_groupi_g39867(csa_tree_add_51_79_groupi_n_6195 ,csa_tree_add_51_79_groupi_n_5115 ,csa_tree_add_51_79_groupi_n_5208);
  xnor csa_tree_add_51_79_groupi_g39868(csa_tree_add_51_79_groupi_n_6194 ,csa_tree_add_51_79_groupi_n_4856 ,csa_tree_add_51_79_groupi_n_5110);
  xnor csa_tree_add_51_79_groupi_g39869(csa_tree_add_51_79_groupi_n_6193 ,csa_tree_add_51_79_groupi_n_5232 ,csa_tree_add_51_79_groupi_n_5238);
  xnor csa_tree_add_51_79_groupi_g39870(csa_tree_add_51_79_groupi_n_6192 ,csa_tree_add_51_79_groupi_n_5477 ,csa_tree_add_51_79_groupi_n_5355);
  xnor csa_tree_add_51_79_groupi_g39871(csa_tree_add_51_79_groupi_n_6191 ,csa_tree_add_51_79_groupi_n_5125 ,csa_tree_add_51_79_groupi_n_4845);
  xnor csa_tree_add_51_79_groupi_g39872(csa_tree_add_51_79_groupi_n_6190 ,csa_tree_add_51_79_groupi_n_5089 ,csa_tree_add_51_79_groupi_n_5334);
  xor csa_tree_add_51_79_groupi_g39873(csa_tree_add_51_79_groupi_n_6189 ,csa_tree_add_51_79_groupi_n_3757 ,csa_tree_add_51_79_groupi_n_5522);
  xnor csa_tree_add_51_79_groupi_g39874(csa_tree_add_51_79_groupi_n_6188 ,csa_tree_add_51_79_groupi_n_5416 ,csa_tree_add_51_79_groupi_n_5521);
  xnor csa_tree_add_51_79_groupi_g39875(csa_tree_add_51_79_groupi_n_6187 ,csa_tree_add_51_79_groupi_n_5384 ,csa_tree_add_51_79_groupi_n_5479);
  xnor csa_tree_add_51_79_groupi_g39876(csa_tree_add_51_79_groupi_n_6186 ,csa_tree_add_51_79_groupi_n_5278 ,csa_tree_add_51_79_groupi_n_5546);
  xnor csa_tree_add_51_79_groupi_g39877(csa_tree_add_51_79_groupi_n_6185 ,csa_tree_add_51_79_groupi_n_5407 ,csa_tree_add_51_79_groupi_n_5408);
  xnor csa_tree_add_51_79_groupi_g39878(csa_tree_add_51_79_groupi_n_6184 ,csa_tree_add_51_79_groupi_n_5569 ,csa_tree_add_51_79_groupi_n_5410);
  xnor csa_tree_add_51_79_groupi_g39879(csa_tree_add_51_79_groupi_n_6183 ,csa_tree_add_51_79_groupi_n_5224 ,csa_tree_add_51_79_groupi_n_5235);
  xnor csa_tree_add_51_79_groupi_g39880(csa_tree_add_51_79_groupi_n_6182 ,csa_tree_add_51_79_groupi_n_5166 ,csa_tree_add_51_79_groupi_n_5168);
  xnor csa_tree_add_51_79_groupi_g39881(csa_tree_add_51_79_groupi_n_6181 ,csa_tree_add_51_79_groupi_n_5153 ,csa_tree_add_51_79_groupi_n_5120);
  xnor csa_tree_add_51_79_groupi_g39882(csa_tree_add_51_79_groupi_n_6180 ,csa_tree_add_51_79_groupi_n_5155 ,csa_tree_add_51_79_groupi_n_5528);
  xnor csa_tree_add_51_79_groupi_g39883(csa_tree_add_51_79_groupi_n_6179 ,csa_tree_add_51_79_groupi_n_5352 ,csa_tree_add_51_79_groupi_n_5544);
  xnor csa_tree_add_51_79_groupi_g39884(csa_tree_add_51_79_groupi_n_6178 ,csa_tree_add_51_79_groupi_n_5102 ,csa_tree_add_51_79_groupi_n_5234);
  xnor csa_tree_add_51_79_groupi_g39885(csa_tree_add_51_79_groupi_n_6177 ,csa_tree_add_51_79_groupi_n_5183 ,csa_tree_add_51_79_groupi_n_5188);
  xnor csa_tree_add_51_79_groupi_g39886(csa_tree_add_51_79_groupi_n_6176 ,csa_tree_add_51_79_groupi_n_5213 ,csa_tree_add_51_79_groupi_n_5214);
  xnor csa_tree_add_51_79_groupi_g39887(csa_tree_add_51_79_groupi_n_6175 ,csa_tree_add_51_79_groupi_n_5283 ,csa_tree_add_51_79_groupi_n_4841);
  xnor csa_tree_add_51_79_groupi_g39888(csa_tree_add_51_79_groupi_n_6174 ,csa_tree_add_51_79_groupi_n_5172 ,csa_tree_add_51_79_groupi_n_5174);
  xnor csa_tree_add_51_79_groupi_g39889(csa_tree_add_51_79_groupi_n_6173 ,csa_tree_add_51_79_groupi_n_5206 ,csa_tree_add_51_79_groupi_n_5539);
  xnor csa_tree_add_51_79_groupi_g39890(csa_tree_add_51_79_groupi_n_6172 ,csa_tree_add_51_79_groupi_n_5191 ,csa_tree_add_51_79_groupi_n_5195);
  xnor csa_tree_add_51_79_groupi_g39891(csa_tree_add_51_79_groupi_n_6171 ,csa_tree_add_51_79_groupi_n_5348 ,csa_tree_add_51_79_groupi_n_5439);
  xnor csa_tree_add_51_79_groupi_g39892(csa_tree_add_51_79_groupi_n_6170 ,csa_tree_add_51_79_groupi_n_5315 ,csa_tree_add_51_79_groupi_n_5551);
  xnor csa_tree_add_51_79_groupi_g39893(csa_tree_add_51_79_groupi_n_6169 ,csa_tree_add_51_79_groupi_n_5553 ,csa_tree_add_51_79_groupi_n_5181);
  xnor csa_tree_add_51_79_groupi_g39894(csa_tree_add_51_79_groupi_n_6168 ,csa_tree_add_51_79_groupi_n_5046 ,csa_tree_add_51_79_groupi_n_4936);
  xnor csa_tree_add_51_79_groupi_g39895(csa_tree_add_51_79_groupi_n_6167 ,csa_tree_add_51_79_groupi_n_5221 ,csa_tree_add_51_79_groupi_n_5194);
  xnor csa_tree_add_51_79_groupi_g39896(csa_tree_add_51_79_groupi_n_6166 ,csa_tree_add_51_79_groupi_n_5373 ,csa_tree_add_51_79_groupi_n_5319);
  xnor csa_tree_add_51_79_groupi_g39897(csa_tree_add_51_79_groupi_n_6165 ,csa_tree_add_51_79_groupi_n_5328 ,csa_tree_add_51_79_groupi_n_5189);
  xnor csa_tree_add_51_79_groupi_g39898(csa_tree_add_51_79_groupi_n_6164 ,csa_tree_add_51_79_groupi_n_5368 ,csa_tree_add_51_79_groupi_n_5349);
  xnor csa_tree_add_51_79_groupi_g39899(csa_tree_add_51_79_groupi_n_6163 ,csa_tree_add_51_79_groupi_n_5358 ,csa_tree_add_51_79_groupi_n_5361);
  xnor csa_tree_add_51_79_groupi_g39900(csa_tree_add_51_79_groupi_n_6162 ,csa_tree_add_51_79_groupi_n_5430 ,csa_tree_add_51_79_groupi_n_5530);
  xor csa_tree_add_51_79_groupi_g39901(csa_tree_add_51_79_groupi_n_6161 ,csa_tree_add_51_79_groupi_n_3758 ,csa_tree_add_51_79_groupi_n_5555);
  xnor csa_tree_add_51_79_groupi_g39902(csa_tree_add_51_79_groupi_n_6160 ,csa_tree_add_51_79_groupi_n_5077 ,csa_tree_add_51_79_groupi_n_4814);
  xor csa_tree_add_51_79_groupi_g39903(csa_tree_add_51_79_groupi_n_6159 ,csa_tree_add_51_79_groupi_n_4860 ,csa_tree_add_51_79_groupi_n_5086);
  xnor csa_tree_add_51_79_groupi_g39904(csa_tree_add_51_79_groupi_n_6158 ,csa_tree_add_51_79_groupi_n_5377 ,csa_tree_add_51_79_groupi_n_5406);
  xnor csa_tree_add_51_79_groupi_g39905(csa_tree_add_51_79_groupi_n_6157 ,csa_tree_add_51_79_groupi_n_5175 ,csa_tree_add_51_79_groupi_n_5205);
  xnor csa_tree_add_51_79_groupi_g39906(csa_tree_add_51_79_groupi_n_6460 ,csa_tree_add_51_79_groupi_n_3205 ,csa_tree_add_51_79_groupi_n_4732);
  xnor csa_tree_add_51_79_groupi_g39907(csa_tree_add_51_79_groupi_n_6459 ,csa_tree_add_51_79_groupi_n_3318 ,csa_tree_add_51_79_groupi_n_4737);
  xnor csa_tree_add_51_79_groupi_g39908(csa_tree_add_51_79_groupi_n_6458 ,csa_tree_add_51_79_groupi_n_3312 ,csa_tree_add_51_79_groupi_n_4730);
  xnor csa_tree_add_51_79_groupi_g39909(csa_tree_add_51_79_groupi_n_6457 ,csa_tree_add_51_79_groupi_n_3220 ,csa_tree_add_51_79_groupi_n_4720);
  xnor csa_tree_add_51_79_groupi_g39910(csa_tree_add_51_79_groupi_n_6456 ,csa_tree_add_51_79_groupi_n_3313 ,csa_tree_add_51_79_groupi_n_4723);
  xnor csa_tree_add_51_79_groupi_g39911(csa_tree_add_51_79_groupi_n_6455 ,csa_tree_add_51_79_groupi_n_8 ,csa_tree_add_51_79_groupi_n_7);
  xnor csa_tree_add_51_79_groupi_g39912(csa_tree_add_51_79_groupi_n_6454 ,csa_tree_add_51_79_groupi_n_3270 ,csa_tree_add_51_79_groupi_n_4733);
  xnor csa_tree_add_51_79_groupi_g39913(csa_tree_add_51_79_groupi_n_6453 ,csa_tree_add_51_79_groupi_n_4800 ,csa_tree_add_51_79_groupi_n_3191);
  xnor csa_tree_add_51_79_groupi_g39915(csa_tree_add_51_79_groupi_n_6452 ,csa_tree_add_51_79_groupi_n_5463 ,csa_tree_add_51_79_groupi_n_5453);
  xnor csa_tree_add_51_79_groupi_g39916(csa_tree_add_51_79_groupi_n_6451 ,csa_tree_add_51_79_groupi_n_5076 ,csa_tree_add_51_79_groupi_n_5558);
  xnor csa_tree_add_51_79_groupi_g39917(csa_tree_add_51_79_groupi_n_6450 ,csa_tree_add_51_79_groupi_n_3261 ,csa_tree_add_51_79_groupi_n_4729);
  xnor csa_tree_add_51_79_groupi_g39919(csa_tree_add_51_79_groupi_n_6449 ,csa_tree_add_51_79_groupi_n_3314 ,csa_tree_add_51_79_groupi_n_4728);
  xnor csa_tree_add_51_79_groupi_g39920(csa_tree_add_51_79_groupi_n_6448 ,csa_tree_add_51_79_groupi_n_3323 ,csa_tree_add_51_79_groupi_n_4716);
  xnor csa_tree_add_51_79_groupi_g39921(csa_tree_add_51_79_groupi_n_6447 ,csa_tree_add_51_79_groupi_n_3332 ,csa_tree_add_51_79_groupi_n_4726);
  xnor csa_tree_add_51_79_groupi_g39922(csa_tree_add_51_79_groupi_n_6446 ,csa_tree_add_51_79_groupi_n_3329 ,csa_tree_add_51_79_groupi_n_4725);
  xnor csa_tree_add_51_79_groupi_g39923(csa_tree_add_51_79_groupi_n_6445 ,csa_tree_add_51_79_groupi_n_5443 ,csa_tree_add_51_79_groupi_n_5034);
  xnor csa_tree_add_51_79_groupi_g39924(csa_tree_add_51_79_groupi_n_6444 ,csa_tree_add_51_79_groupi_n_3217 ,csa_tree_add_51_79_groupi_n_4727);
  xnor csa_tree_add_51_79_groupi_g39925(csa_tree_add_51_79_groupi_n_6443 ,csa_tree_add_51_79_groupi_n_3316 ,csa_tree_add_51_79_groupi_n_4722);
  xnor csa_tree_add_51_79_groupi_g39926(csa_tree_add_51_79_groupi_n_6442 ,csa_tree_add_51_79_groupi_n_5534 ,csa_tree_add_51_79_groupi_n_4744);
  xnor csa_tree_add_51_79_groupi_g39927(csa_tree_add_51_79_groupi_n_6441 ,csa_tree_add_51_79_groupi_n_3321 ,csa_tree_add_51_79_groupi_n_4721);
  xnor csa_tree_add_51_79_groupi_g39928(csa_tree_add_51_79_groupi_n_6440 ,csa_tree_add_51_79_groupi_n_3324 ,csa_tree_add_51_79_groupi_n_4724);
  xnor csa_tree_add_51_79_groupi_g39929(csa_tree_add_51_79_groupi_n_6439 ,csa_tree_add_51_79_groupi_n_3225 ,csa_tree_add_51_79_groupi_n_4719);
  xnor csa_tree_add_51_79_groupi_g39930(csa_tree_add_51_79_groupi_n_6438 ,csa_tree_add_51_79_groupi_n_3328 ,csa_tree_add_51_79_groupi_n_4717);
  xnor csa_tree_add_51_79_groupi_g39931(csa_tree_add_51_79_groupi_n_6437 ,csa_tree_add_51_79_groupi_n_5103 ,csa_tree_add_51_79_groupi_n_4738);
  xnor csa_tree_add_51_79_groupi_g39932(csa_tree_add_51_79_groupi_n_6435 ,csa_tree_add_51_79_groupi_n_3331 ,csa_tree_add_51_79_groupi_n_4734);
  xnor csa_tree_add_51_79_groupi_g39933(csa_tree_add_51_79_groupi_n_6434 ,csa_tree_add_51_79_groupi_n_4806 ,csa_tree_add_51_79_groupi_n_3193);
  xnor csa_tree_add_51_79_groupi_g39934(csa_tree_add_51_79_groupi_n_6433 ,csa_tree_add_51_79_groupi_n_4807 ,csa_tree_add_51_79_groupi_n_3192);
  xnor csa_tree_add_51_79_groupi_g39935(csa_tree_add_51_79_groupi_n_6432 ,csa_tree_add_51_79_groupi_n_4800 ,csa_tree_add_51_79_groupi_n_1178);
  xnor csa_tree_add_51_79_groupi_g39936(csa_tree_add_51_79_groupi_n_6431 ,csa_tree_add_51_79_groupi_n_4806 ,csa_tree_add_51_79_groupi_n_1176);
  xnor csa_tree_add_51_79_groupi_g39937(csa_tree_add_51_79_groupi_n_6430 ,csa_tree_add_51_79_groupi_n_4807 ,csa_tree_add_51_79_groupi_n_1174);
  xnor csa_tree_add_51_79_groupi_g39938(csa_tree_add_51_79_groupi_n_6428 ,csa_tree_add_51_79_groupi_n_3833 ,csa_tree_add_51_79_groupi_n_4715);
  xnor csa_tree_add_51_79_groupi_g39939(csa_tree_add_51_79_groupi_n_6426 ,csa_tree_add_51_79_groupi_n_5499 ,csa_tree_add_51_79_groupi_n_4739);
  xnor csa_tree_add_51_79_groupi_g39940(csa_tree_add_51_79_groupi_n_6424 ,csa_tree_add_51_79_groupi_n_5571 ,csa_tree_add_51_79_groupi_n_4748);
  xnor csa_tree_add_51_79_groupi_g39941(csa_tree_add_51_79_groupi_n_6422 ,csa_tree_add_51_79_groupi_n_3828 ,csa_tree_add_51_79_groupi_n_5434);
  xnor csa_tree_add_51_79_groupi_g39942(csa_tree_add_51_79_groupi_n_6420 ,csa_tree_add_51_79_groupi_n_5549 ,csa_tree_add_51_79_groupi_n_4747);
  xnor csa_tree_add_51_79_groupi_g39943(csa_tree_add_51_79_groupi_n_6418 ,csa_tree_add_51_79_groupi_n_3334 ,csa_tree_add_51_79_groupi_n_4746);
  xnor csa_tree_add_51_79_groupi_g39944(csa_tree_add_51_79_groupi_n_6416 ,csa_tree_add_51_79_groupi_n_3298 ,csa_tree_add_51_79_groupi_n_4736);
  xnor csa_tree_add_51_79_groupi_g39945(csa_tree_add_51_79_groupi_n_6415 ,csa_tree_add_51_79_groupi_n_3327 ,csa_tree_add_51_79_groupi_n_4745);
  xnor csa_tree_add_51_79_groupi_g39946(csa_tree_add_51_79_groupi_n_6413 ,csa_tree_add_51_79_groupi_n_3832 ,csa_tree_add_51_79_groupi_n_4743);
  xnor csa_tree_add_51_79_groupi_g39947(csa_tree_add_51_79_groupi_n_6412 ,csa_tree_add_51_79_groupi_n_3830 ,csa_tree_add_51_79_groupi_n_4714);
  xnor csa_tree_add_51_79_groupi_g39948(csa_tree_add_51_79_groupi_n_6410 ,csa_tree_add_51_79_groupi_n_3310 ,csa_tree_add_51_79_groupi_n_4735);
  xnor csa_tree_add_51_79_groupi_g39949(csa_tree_add_51_79_groupi_n_6409 ,csa_tree_add_51_79_groupi_n_5109 ,csa_tree_add_51_79_groupi_n_4741);
  xnor csa_tree_add_51_79_groupi_g39950(csa_tree_add_51_79_groupi_n_6407 ,csa_tree_add_51_79_groupi_n_3317 ,csa_tree_add_51_79_groupi_n_4742);
  xnor csa_tree_add_51_79_groupi_g39951(csa_tree_add_51_79_groupi_n_6405 ,csa_tree_add_51_79_groupi_n_3831 ,csa_tree_add_51_79_groupi_n_4731);
  xnor csa_tree_add_51_79_groupi_g39952(csa_tree_add_51_79_groupi_n_6404 ,csa_tree_add_51_79_groupi_n_5091 ,csa_tree_add_51_79_groupi_n_4749);
  xnor csa_tree_add_51_79_groupi_g39953(csa_tree_add_51_79_groupi_n_6402 ,csa_tree_add_51_79_groupi_n_3330 ,csa_tree_add_51_79_groupi_n_4740);
  and csa_tree_add_51_79_groupi_g39954(csa_tree_add_51_79_groupi_n_6400 ,csa_tree_add_51_79_groupi_n_4785 ,csa_tree_add_51_79_groupi_n_5787);
  xnor csa_tree_add_51_79_groupi_g39955(csa_tree_add_51_79_groupi_n_6399 ,csa_tree_add_51_79_groupi_n_5509 ,csa_tree_add_51_79_groupi_n_4718);
  and csa_tree_add_51_79_groupi_g39956(csa_tree_add_51_79_groupi_n_6396 ,csa_tree_add_51_79_groupi_n_4773 ,csa_tree_add_51_79_groupi_n_5817);
  and csa_tree_add_51_79_groupi_g39957(csa_tree_add_51_79_groupi_n_6394 ,csa_tree_add_51_79_groupi_n_4784 ,csa_tree_add_51_79_groupi_n_5799);
  not csa_tree_add_51_79_groupi_g39958(csa_tree_add_51_79_groupi_n_6142 ,csa_tree_add_51_79_groupi_n_6143);
  not csa_tree_add_51_79_groupi_g39959(csa_tree_add_51_79_groupi_n_6135 ,csa_tree_add_51_79_groupi_n_6136);
  not csa_tree_add_51_79_groupi_g39960(csa_tree_add_51_79_groupi_n_6133 ,csa_tree_add_51_79_groupi_n_6134);
  not csa_tree_add_51_79_groupi_g39961(csa_tree_add_51_79_groupi_n_6130 ,csa_tree_add_51_79_groupi_n_6131);
  nor csa_tree_add_51_79_groupi_g39962(csa_tree_add_51_79_groupi_n_6126 ,csa_tree_add_51_79_groupi_n_4573 ,csa_tree_add_51_79_groupi_n_5534);
  or csa_tree_add_51_79_groupi_g39963(csa_tree_add_51_79_groupi_n_6125 ,csa_tree_add_51_79_groupi_n_3256 ,csa_tree_add_51_79_groupi_n_5153);
  and csa_tree_add_51_79_groupi_g39964(csa_tree_add_51_79_groupi_n_6124 ,csa_tree_add_51_79_groupi_n_4976 ,csa_tree_add_51_79_groupi_n_4977);
  or csa_tree_add_51_79_groupi_g39965(csa_tree_add_51_79_groupi_n_6123 ,csa_tree_add_51_79_groupi_n_3766 ,csa_tree_add_51_79_groupi_n_5316);
  or csa_tree_add_51_79_groupi_g39966(csa_tree_add_51_79_groupi_n_6122 ,csa_tree_add_51_79_groupi_n_4980 ,csa_tree_add_51_79_groupi_n_5156);
  or csa_tree_add_51_79_groupi_g39967(csa_tree_add_51_79_groupi_n_6121 ,csa_tree_add_51_79_groupi_n_4815 ,csa_tree_add_51_79_groupi_n_4816);
  or csa_tree_add_51_79_groupi_g39968(csa_tree_add_51_79_groupi_n_6120 ,csa_tree_add_51_79_groupi_n_5386 ,csa_tree_add_51_79_groupi_n_5348);
  or csa_tree_add_51_79_groupi_g39969(csa_tree_add_51_79_groupi_n_6119 ,csa_tree_add_51_79_groupi_n_3741 ,csa_tree_add_51_79_groupi_n_5242);
  and csa_tree_add_51_79_groupi_g39970(csa_tree_add_51_79_groupi_n_6118 ,csa_tree_add_51_79_groupi_n_3758 ,csa_tree_add_51_79_groupi_n_765);
  and csa_tree_add_51_79_groupi_g39971(csa_tree_add_51_79_groupi_n_6117 ,csa_tree_add_51_79_groupi_n_4905 ,csa_tree_add_51_79_groupi_n_5249);
  or csa_tree_add_51_79_groupi_g39972(csa_tree_add_51_79_groupi_n_6116 ,csa_tree_add_51_79_groupi_n_4986 ,csa_tree_add_51_79_groupi_n_5161);
  nor csa_tree_add_51_79_groupi_g39973(csa_tree_add_51_79_groupi_n_6115 ,csa_tree_add_51_79_groupi_n_3767 ,csa_tree_add_51_79_groupi_n_5317);
  and csa_tree_add_51_79_groupi_g39974(csa_tree_add_51_79_groupi_n_6114 ,csa_tree_add_51_79_groupi_n_5204 ,csa_tree_add_51_79_groupi_n_5273);
  nor csa_tree_add_51_79_groupi_g39975(csa_tree_add_51_79_groupi_n_6113 ,csa_tree_add_51_79_groupi_n_3758 ,csa_tree_add_51_79_groupi_n_4793);
  or csa_tree_add_51_79_groupi_g39976(csa_tree_add_51_79_groupi_n_6112 ,csa_tree_add_51_79_groupi_n_5260 ,csa_tree_add_51_79_groupi_n_5431);
  or csa_tree_add_51_79_groupi_g39977(csa_tree_add_51_79_groupi_n_6111 ,csa_tree_add_51_79_groupi_n_3764 ,csa_tree_add_51_79_groupi_n_5201);
  nor csa_tree_add_51_79_groupi_g39978(csa_tree_add_51_79_groupi_n_6110 ,csa_tree_add_51_79_groupi_n_5271 ,csa_tree_add_51_79_groupi_n_5396);
  or csa_tree_add_51_79_groupi_g39979(csa_tree_add_51_79_groupi_n_6109 ,csa_tree_add_51_79_groupi_n_4981 ,csa_tree_add_51_79_groupi_n_5180);
  nor csa_tree_add_51_79_groupi_g39980(csa_tree_add_51_79_groupi_n_6108 ,csa_tree_add_51_79_groupi_n_3765 ,csa_tree_add_51_79_groupi_n_5200);
  or csa_tree_add_51_79_groupi_g39981(csa_tree_add_51_79_groupi_n_6107 ,csa_tree_add_51_79_groupi_n_5406 ,csa_tree_add_51_79_groupi_n_5377);
  or csa_tree_add_51_79_groupi_g39982(csa_tree_add_51_79_groupi_n_6106 ,csa_tree_add_51_79_groupi_n_3788 ,csa_tree_add_51_79_groupi_n_5300);
  or csa_tree_add_51_79_groupi_g39983(csa_tree_add_51_79_groupi_n_6105 ,csa_tree_add_51_79_groupi_n_3814 ,csa_tree_add_51_79_groupi_n_4845);
  and csa_tree_add_51_79_groupi_g39984(csa_tree_add_51_79_groupi_n_6104 ,csa_tree_add_51_79_groupi_n_6 ,csa_tree_add_51_79_groupi_n_2);
  and csa_tree_add_51_79_groupi_g39985(csa_tree_add_51_79_groupi_n_6103 ,csa_tree_add_51_79_groupi_n_5406 ,csa_tree_add_51_79_groupi_n_5377);
  or csa_tree_add_51_79_groupi_g39986(csa_tree_add_51_79_groupi_n_6102 ,csa_tree_add_51_79_groupi_n_3768 ,csa_tree_add_51_79_groupi_n_5332);
  or csa_tree_add_51_79_groupi_g39987(csa_tree_add_51_79_groupi_n_6101 ,csa_tree_add_51_79_groupi_n_4813 ,csa_tree_add_51_79_groupi_n_5187);
  nor csa_tree_add_51_79_groupi_g39988(csa_tree_add_51_79_groupi_n_6100 ,csa_tree_add_51_79_groupi_n_5432 ,csa_tree_add_51_79_groupi_n_5259);
  or csa_tree_add_51_79_groupi_g39989(csa_tree_add_51_79_groupi_n_6099 ,csa_tree_add_51_79_groupi_n_5205 ,csa_tree_add_51_79_groupi_n_5175);
  nor csa_tree_add_51_79_groupi_g39990(csa_tree_add_51_79_groupi_n_6098 ,csa_tree_add_51_79_groupi_n_3769 ,csa_tree_add_51_79_groupi_n_5331);
  or csa_tree_add_51_79_groupi_g39991(csa_tree_add_51_79_groupi_n_6097 ,csa_tree_add_51_79_groupi_n_4992 ,csa_tree_add_51_79_groupi_n_5203);
  and csa_tree_add_51_79_groupi_g39992(csa_tree_add_51_79_groupi_n_6096 ,csa_tree_add_51_79_groupi_n_4992 ,csa_tree_add_51_79_groupi_n_5203);
  or csa_tree_add_51_79_groupi_g39993(csa_tree_add_51_79_groupi_n_6095 ,csa_tree_add_51_79_groupi_n_3285 ,csa_tree_add_51_79_groupi_n_5426);
  or csa_tree_add_51_79_groupi_g39994(csa_tree_add_51_79_groupi_n_6094 ,csa_tree_add_51_79_groupi_n_4997 ,csa_tree_add_51_79_groupi_n_5428);
  and csa_tree_add_51_79_groupi_g39995(csa_tree_add_51_79_groupi_n_6093 ,csa_tree_add_51_79_groupi_n_4997 ,csa_tree_add_51_79_groupi_n_5428);
  or csa_tree_add_51_79_groupi_g39996(csa_tree_add_51_79_groupi_n_6092 ,csa_tree_add_51_79_groupi_n_5405 ,csa_tree_add_51_79_groupi_n_5391);
  nor csa_tree_add_51_79_groupi_g39997(csa_tree_add_51_79_groupi_n_6091 ,csa_tree_add_51_79_groupi_n_3286 ,csa_tree_add_51_79_groupi_n_5425);
  or csa_tree_add_51_79_groupi_g39998(csa_tree_add_51_79_groupi_n_6090 ,csa_tree_add_51_79_groupi_n_5385 ,csa_tree_add_51_79_groupi_n_5384);
  and csa_tree_add_51_79_groupi_g39999(csa_tree_add_51_79_groupi_n_6089 ,csa_tree_add_51_79_groupi_n_5405 ,csa_tree_add_51_79_groupi_n_5391);
  and csa_tree_add_51_79_groupi_g40000(csa_tree_add_51_79_groupi_n_6088 ,csa_tree_add_51_79_groupi_n_5205 ,csa_tree_add_51_79_groupi_n_5175);
  or csa_tree_add_51_79_groupi_g40001(csa_tree_add_51_79_groupi_n_6087 ,csa_tree_add_51_79_groupi_n_5382 ,csa_tree_add_51_79_groupi_n_5378);
  nor csa_tree_add_51_79_groupi_g40002(csa_tree_add_51_79_groupi_n_6086 ,csa_tree_add_51_79_groupi_n_3789 ,csa_tree_add_51_79_groupi_n_5299);
  or csa_tree_add_51_79_groupi_g40003(csa_tree_add_51_79_groupi_n_6085 ,csa_tree_add_51_79_groupi_n_5257 ,csa_tree_add_51_79_groupi_n_5254);
  or csa_tree_add_51_79_groupi_g40004(csa_tree_add_51_79_groupi_n_6084 ,csa_tree_add_51_79_groupi_n_5363 ,csa_tree_add_51_79_groupi_n_5288);
  and csa_tree_add_51_79_groupi_g40005(csa_tree_add_51_79_groupi_n_6083 ,csa_tree_add_51_79_groupi_n_5382 ,csa_tree_add_51_79_groupi_n_5378);
  and csa_tree_add_51_79_groupi_g40006(csa_tree_add_51_79_groupi_n_6082 ,csa_tree_add_51_79_groupi_n_4917 ,csa_tree_add_51_79_groupi_n_5246);
  and csa_tree_add_51_79_groupi_g40007(csa_tree_add_51_79_groupi_n_6081 ,csa_tree_add_51_79_groupi_n_5385 ,csa_tree_add_51_79_groupi_n_5384);
  or csa_tree_add_51_79_groupi_g40008(csa_tree_add_51_79_groupi_n_6080 ,csa_tree_add_51_79_groupi_n_3793 ,csa_tree_add_51_79_groupi_n_5355);
  nor csa_tree_add_51_79_groupi_g40009(csa_tree_add_51_79_groupi_n_6079 ,csa_tree_add_51_79_groupi_n_3794 ,csa_tree_add_51_79_groupi_n_5354);
  or csa_tree_add_51_79_groupi_g40010(csa_tree_add_51_79_groupi_n_6078 ,csa_tree_add_51_79_groupi_n_4905 ,csa_tree_add_51_79_groupi_n_5249);
  and csa_tree_add_51_79_groupi_g40011(csa_tree_add_51_79_groupi_n_6077 ,csa_tree_add_51_79_groupi_n_4996 ,csa_tree_add_51_79_groupi_n_5196);
  and csa_tree_add_51_79_groupi_g40012(csa_tree_add_51_79_groupi_n_6076 ,csa_tree_add_51_79_groupi_n_5256 ,csa_tree_add_51_79_groupi_n_5253);
  or csa_tree_add_51_79_groupi_g40013(csa_tree_add_51_79_groupi_n_6075 ,csa_tree_add_51_79_groupi_n_3791 ,csa_tree_add_51_79_groupi_n_5287);
  or csa_tree_add_51_79_groupi_g40014(csa_tree_add_51_79_groupi_n_6074 ,csa_tree_add_51_79_groupi_n_4999 ,csa_tree_add_51_79_groupi_n_5263);
  nor csa_tree_add_51_79_groupi_g40015(csa_tree_add_51_79_groupi_n_6073 ,csa_tree_add_51_79_groupi_n_3792 ,csa_tree_add_51_79_groupi_n_5286);
  or csa_tree_add_51_79_groupi_g40016(csa_tree_add_51_79_groupi_n_6072 ,csa_tree_add_51_79_groupi_n_5251 ,csa_tree_add_51_79_groupi_n_5245);
  and csa_tree_add_51_79_groupi_g40017(csa_tree_add_51_79_groupi_n_6071 ,csa_tree_add_51_79_groupi_n_4999 ,csa_tree_add_51_79_groupi_n_5263);
  or csa_tree_add_51_79_groupi_g40018(csa_tree_add_51_79_groupi_n_6070 ,csa_tree_add_51_79_groupi_n_5235 ,csa_tree_add_51_79_groupi_n_5224);
  and csa_tree_add_51_79_groupi_g40019(csa_tree_add_51_79_groupi_n_6069 ,csa_tree_add_51_79_groupi_n_5235 ,csa_tree_add_51_79_groupi_n_5224);
  or csa_tree_add_51_79_groupi_g40020(csa_tree_add_51_79_groupi_n_6068 ,csa_tree_add_51_79_groupi_n_5002 ,csa_tree_add_51_79_groupi_n_5190);
  and csa_tree_add_51_79_groupi_g40021(csa_tree_add_51_79_groupi_n_6067 ,csa_tree_add_51_79_groupi_n_5251 ,csa_tree_add_51_79_groupi_n_5245);
  and csa_tree_add_51_79_groupi_g40022(csa_tree_add_51_79_groupi_n_6066 ,csa_tree_add_51_79_groupi_n_5002 ,csa_tree_add_51_79_groupi_n_5190);
  or csa_tree_add_51_79_groupi_g40023(csa_tree_add_51_79_groupi_n_6065 ,csa_tree_add_51_79_groupi_n_5168 ,csa_tree_add_51_79_groupi_n_5166);
  and csa_tree_add_51_79_groupi_g40024(csa_tree_add_51_79_groupi_n_6064 ,csa_tree_add_51_79_groupi_n_5168 ,csa_tree_add_51_79_groupi_n_5166);
  or csa_tree_add_51_79_groupi_g40025(csa_tree_add_51_79_groupi_n_6063 ,csa_tree_add_51_79_groupi_n_5433 ,csa_tree_add_51_79_groupi_n_5429);
  and csa_tree_add_51_79_groupi_g40026(csa_tree_add_51_79_groupi_n_6062 ,csa_tree_add_51_79_groupi_n_5433 ,csa_tree_add_51_79_groupi_n_5429);
  or csa_tree_add_51_79_groupi_g40027(csa_tree_add_51_79_groupi_n_6061 ,csa_tree_add_51_79_groupi_n_5006 ,csa_tree_add_51_79_groupi_n_5427);
  and csa_tree_add_51_79_groupi_g40028(csa_tree_add_51_79_groupi_n_6060 ,csa_tree_add_51_79_groupi_n_5006 ,csa_tree_add_51_79_groupi_n_5427);
  and csa_tree_add_51_79_groupi_g40029(csa_tree_add_51_79_groupi_n_6059 ,csa_tree_add_51_79_groupi_n_4603 ,csa_tree_add_51_79_groupi_n_5571);
  or csa_tree_add_51_79_groupi_g40030(csa_tree_add_51_79_groupi_n_6058 ,csa_tree_add_51_79_groupi_n_4906 ,csa_tree_add_51_79_groupi_n_5424);
  and csa_tree_add_51_79_groupi_g40031(csa_tree_add_51_79_groupi_n_6057 ,csa_tree_add_51_79_groupi_n_4906 ,csa_tree_add_51_79_groupi_n_5424);
  or csa_tree_add_51_79_groupi_g40032(csa_tree_add_51_79_groupi_n_6056 ,csa_tree_add_51_79_groupi_n_5008 ,csa_tree_add_51_79_groupi_n_5421);
  and csa_tree_add_51_79_groupi_g40033(csa_tree_add_51_79_groupi_n_6055 ,csa_tree_add_51_79_groupi_n_5008 ,csa_tree_add_51_79_groupi_n_5421);
  nor csa_tree_add_51_79_groupi_g40034(csa_tree_add_51_79_groupi_n_6054 ,csa_tree_add_51_79_groupi_n_5364 ,csa_tree_add_51_79_groupi_n_5289);
  or csa_tree_add_51_79_groupi_g40035(csa_tree_add_51_79_groupi_n_6053 ,csa_tree_add_51_79_groupi_n_4953 ,csa_tree_add_51_79_groupi_n_5247);
  and csa_tree_add_51_79_groupi_g40036(csa_tree_add_51_79_groupi_n_6052 ,csa_tree_add_51_79_groupi_n_4953 ,csa_tree_add_51_79_groupi_n_5247);
  and csa_tree_add_51_79_groupi_g40037(csa_tree_add_51_79_groupi_n_6051 ,csa_tree_add_51_79_groupi_n_3742 ,csa_tree_add_51_79_groupi_n_5321);
  or csa_tree_add_51_79_groupi_g40038(csa_tree_add_51_79_groupi_n_6050 ,csa_tree_add_51_79_groupi_n_3809 ,csa_tree_add_51_79_groupi_n_5410);
  or csa_tree_add_51_79_groupi_g40039(csa_tree_add_51_79_groupi_n_6049 ,csa_tree_add_51_79_groupi_n_5007 ,csa_tree_add_51_79_groupi_n_5414);
  or csa_tree_add_51_79_groupi_g40040(csa_tree_add_51_79_groupi_n_6048 ,csa_tree_add_51_79_groupi_n_5339 ,csa_tree_add_51_79_groupi_n_5340);
  and csa_tree_add_51_79_groupi_g40041(csa_tree_add_51_79_groupi_n_6047 ,csa_tree_add_51_79_groupi_n_5339 ,csa_tree_add_51_79_groupi_n_5340);
  and csa_tree_add_51_79_groupi_g40042(csa_tree_add_51_79_groupi_n_6046 ,csa_tree_add_51_79_groupi_n_5408 ,csa_tree_add_51_79_groupi_n_5407);
  or csa_tree_add_51_79_groupi_g40043(csa_tree_add_51_79_groupi_n_6045 ,csa_tree_add_51_79_groupi_n_4975 ,csa_tree_add_51_79_groupi_n_5330);
  nor csa_tree_add_51_79_groupi_g40044(csa_tree_add_51_79_groupi_n_6044 ,csa_tree_add_51_79_groupi_n_3810 ,csa_tree_add_51_79_groupi_n_5409);
  or csa_tree_add_51_79_groupi_g40045(csa_tree_add_51_79_groupi_n_6043 ,csa_tree_add_51_79_groupi_n_5256 ,csa_tree_add_51_79_groupi_n_5253);
  or csa_tree_add_51_79_groupi_g40046(csa_tree_add_51_79_groupi_n_6042 ,csa_tree_add_51_79_groupi_n_5341 ,csa_tree_add_51_79_groupi_n_5394);
  or csa_tree_add_51_79_groupi_g40047(csa_tree_add_51_79_groupi_n_6041 ,csa_tree_add_51_79_groupi_n_4393 ,csa_tree_add_51_79_groupi_n_5117);
  and csa_tree_add_51_79_groupi_g40048(csa_tree_add_51_79_groupi_n_6040 ,csa_tree_add_51_79_groupi_n_4990 ,csa_tree_add_51_79_groupi_n_5158);
  and csa_tree_add_51_79_groupi_g40049(csa_tree_add_51_79_groupi_n_6039 ,csa_tree_add_51_79_groupi_n_5341 ,csa_tree_add_51_79_groupi_n_5394);
  or csa_tree_add_51_79_groupi_g40050(csa_tree_add_51_79_groupi_n_6038 ,csa_tree_add_51_79_groupi_n_3239 ,csa_tree_add_51_79_groupi_n_5376);
  nor csa_tree_add_51_79_groupi_g40051(csa_tree_add_51_79_groupi_n_6037 ,csa_tree_add_51_79_groupi_n_3742 ,csa_tree_add_51_79_groupi_n_5321);
  or csa_tree_add_51_79_groupi_g40052(csa_tree_add_51_79_groupi_n_6036 ,csa_tree_add_51_79_groupi_n_3805 ,csa_tree_add_51_79_groupi_n_5375);
  nor csa_tree_add_51_79_groupi_g40053(csa_tree_add_51_79_groupi_n_6035 ,csa_tree_add_51_79_groupi_n_3806 ,csa_tree_add_51_79_groupi_n_5374);
  or csa_tree_add_51_79_groupi_g40054(csa_tree_add_51_79_groupi_n_6034 ,csa_tree_add_51_79_groupi_n_5314 ,csa_tree_add_51_79_groupi_n_5346);
  and csa_tree_add_51_79_groupi_g40055(csa_tree_add_51_79_groupi_n_6033 ,csa_tree_add_51_79_groupi_n_4960 ,csa_tree_add_51_79_groupi_n_5261);
  and csa_tree_add_51_79_groupi_g40056(csa_tree_add_51_79_groupi_n_6032 ,csa_tree_add_51_79_groupi_n_5386 ,csa_tree_add_51_79_groupi_n_5348);
  or csa_tree_add_51_79_groupi_g40057(csa_tree_add_51_79_groupi_n_6031 ,csa_tree_add_51_79_groupi_n_5345 ,csa_tree_add_51_79_groupi_n_5344);
  and csa_tree_add_51_79_groupi_g40058(csa_tree_add_51_79_groupi_n_6030 ,csa_tree_add_51_79_groupi_n_5345 ,csa_tree_add_51_79_groupi_n_5344);
  or csa_tree_add_51_79_groupi_g40059(csa_tree_add_51_79_groupi_n_6029 ,csa_tree_add_51_79_groupi_n_5181 ,csa_tree_add_51_79_groupi_n_5324);
  nor csa_tree_add_51_79_groupi_g40060(csa_tree_add_51_79_groupi_n_6028 ,csa_tree_add_51_79_groupi_n_3233 ,csa_tree_add_51_79_groupi_n_5362);
  nor csa_tree_add_51_79_groupi_g40061(csa_tree_add_51_79_groupi_n_6027 ,csa_tree_add_51_79_groupi_n_5347 ,csa_tree_add_51_79_groupi_n_5313);
  or csa_tree_add_51_79_groupi_g40062(csa_tree_add_51_79_groupi_n_6026 ,csa_tree_add_51_79_groupi_n_4881 ,csa_tree_add_51_79_groupi_n_5318);
  and csa_tree_add_51_79_groupi_g40063(csa_tree_add_51_79_groupi_n_6025 ,csa_tree_add_51_79_groupi_n_5181 ,csa_tree_add_51_79_groupi_n_5324);
  or csa_tree_add_51_79_groupi_g40064(csa_tree_add_51_79_groupi_n_6024 ,csa_tree_add_51_79_groupi_n_4892 ,csa_tree_add_51_79_groupi_n_5302);
  or csa_tree_add_51_79_groupi_g40065(csa_tree_add_51_79_groupi_n_6023 ,csa_tree_add_51_79_groupi_n_4861 ,csa_tree_add_51_79_groupi_n_5315);
  and csa_tree_add_51_79_groupi_g40066(csa_tree_add_51_79_groupi_n_6022 ,csa_tree_add_51_79_groupi_n_4881 ,csa_tree_add_51_79_groupi_n_5318);
  or csa_tree_add_51_79_groupi_g40067(csa_tree_add_51_79_groupi_n_6021 ,csa_tree_add_51_79_groupi_n_5001 ,csa_tree_add_51_79_groupi_n_5312);
  and csa_tree_add_51_79_groupi_g40068(csa_tree_add_51_79_groupi_n_6020 ,csa_tree_add_51_79_groupi_n_4534 ,csa_tree_add_51_79_groupi_n_5549);
  and csa_tree_add_51_79_groupi_g40069(csa_tree_add_51_79_groupi_n_6019 ,csa_tree_add_51_79_groupi_n_5001 ,csa_tree_add_51_79_groupi_n_5312);
  or csa_tree_add_51_79_groupi_g40070(csa_tree_add_51_79_groupi_n_6018 ,csa_tree_add_51_79_groupi_n_4841 ,csa_tree_add_51_79_groupi_n_5283);
  or csa_tree_add_51_79_groupi_g40071(csa_tree_add_51_79_groupi_n_6017 ,csa_tree_add_51_79_groupi_n_3756 ,csa_tree_add_51_79_groupi_n_5178);
  and csa_tree_add_51_79_groupi_g40072(csa_tree_add_51_79_groupi_n_6016 ,csa_tree_add_51_79_groupi_n_4861 ,csa_tree_add_51_79_groupi_n_5315);
  or csa_tree_add_51_79_groupi_g40073(csa_tree_add_51_79_groupi_n_6015 ,csa_tree_add_51_79_groupi_n_5282 ,csa_tree_add_51_79_groupi_n_5278);
  and csa_tree_add_51_79_groupi_g40074(csa_tree_add_51_79_groupi_n_6014 ,csa_tree_add_51_79_groupi_n_4841 ,csa_tree_add_51_79_groupi_n_5283);
  or csa_tree_add_51_79_groupi_g40075(csa_tree_add_51_79_groupi_n_6013 ,csa_tree_add_51_79_groupi_n_5277 ,csa_tree_add_51_79_groupi_n_5276);
  and csa_tree_add_51_79_groupi_g40076(csa_tree_add_51_79_groupi_n_6012 ,csa_tree_add_51_79_groupi_n_5282 ,csa_tree_add_51_79_groupi_n_5278);
  and csa_tree_add_51_79_groupi_g40077(csa_tree_add_51_79_groupi_n_6011 ,csa_tree_add_51_79_groupi_n_5277 ,csa_tree_add_51_79_groupi_n_5276);
  nor csa_tree_add_51_79_groupi_g40078(csa_tree_add_51_79_groupi_n_6010 ,csa_tree_add_51_79_groupi_n_5303 ,csa_tree_add_51_79_groupi_n_4891);
  or csa_tree_add_51_79_groupi_g40079(csa_tree_add_51_79_groupi_n_6009 ,csa_tree_add_51_79_groupi_n_3237 ,csa_tree_add_51_79_groupi_n_5244);
  or csa_tree_add_51_79_groupi_g40080(csa_tree_add_51_79_groupi_n_6008 ,csa_tree_add_51_79_groupi_n_5000 ,csa_tree_add_51_79_groupi_n_5248);
  and csa_tree_add_51_79_groupi_g40081(csa_tree_add_51_79_groupi_n_6007 ,csa_tree_add_51_79_groupi_n_5000 ,csa_tree_add_51_79_groupi_n_5248);
  or csa_tree_add_51_79_groupi_g40082(csa_tree_add_51_79_groupi_n_6006 ,csa_tree_add_51_79_groupi_n_5194 ,csa_tree_add_51_79_groupi_n_5221);
  nor csa_tree_add_51_79_groupi_g40083(csa_tree_add_51_79_groupi_n_6005 ,csa_tree_add_51_79_groupi_n_3238 ,csa_tree_add_51_79_groupi_n_5243);
  and csa_tree_add_51_79_groupi_g40084(csa_tree_add_51_79_groupi_n_6004 ,csa_tree_add_51_79_groupi_n_5194 ,csa_tree_add_51_79_groupi_n_5221);
  or csa_tree_add_51_79_groupi_g40085(csa_tree_add_51_79_groupi_n_6003 ,csa_tree_add_51_79_groupi_n_5215 ,csa_tree_add_51_79_groupi_n_5206);
  or csa_tree_add_51_79_groupi_g40086(csa_tree_add_51_79_groupi_n_6002 ,csa_tree_add_51_79_groupi_n_5214 ,csa_tree_add_51_79_groupi_n_5213);
  or csa_tree_add_51_79_groupi_g40087(csa_tree_add_51_79_groupi_n_6001 ,csa_tree_add_51_79_groupi_n_4818 ,csa_tree_add_51_79_groupi_n_4819);
  and csa_tree_add_51_79_groupi_g40088(csa_tree_add_51_79_groupi_n_6000 ,csa_tree_add_51_79_groupi_n_5214 ,csa_tree_add_51_79_groupi_n_5213);
  or csa_tree_add_51_79_groupi_g40089(csa_tree_add_51_79_groupi_n_5999 ,csa_tree_add_51_79_groupi_n_4998 ,csa_tree_add_51_79_groupi_n_5202);
  or csa_tree_add_51_79_groupi_g40090(csa_tree_add_51_79_groupi_n_5998 ,csa_tree_add_51_79_groupi_n_5199 ,csa_tree_add_51_79_groupi_n_5185);
  and csa_tree_add_51_79_groupi_g40091(csa_tree_add_51_79_groupi_n_5997 ,csa_tree_add_51_79_groupi_n_5215 ,csa_tree_add_51_79_groupi_n_5206);
  or csa_tree_add_51_79_groupi_g40092(csa_tree_add_51_79_groupi_n_5996 ,csa_tree_add_51_79_groupi_n_5198 ,csa_tree_add_51_79_groupi_n_5193);
  and csa_tree_add_51_79_groupi_g40093(csa_tree_add_51_79_groupi_n_5995 ,csa_tree_add_51_79_groupi_n_4998 ,csa_tree_add_51_79_groupi_n_5202);
  or csa_tree_add_51_79_groupi_g40094(csa_tree_add_51_79_groupi_n_5994 ,csa_tree_add_51_79_groupi_n_5195 ,csa_tree_add_51_79_groupi_n_5191);
  and csa_tree_add_51_79_groupi_g40095(csa_tree_add_51_79_groupi_n_5993 ,csa_tree_add_51_79_groupi_n_5195 ,csa_tree_add_51_79_groupi_n_5191);
  and csa_tree_add_51_79_groupi_g40096(csa_tree_add_51_79_groupi_n_5992 ,csa_tree_add_51_79_groupi_n_5198 ,csa_tree_add_51_79_groupi_n_5193);
  or csa_tree_add_51_79_groupi_g40097(csa_tree_add_51_79_groupi_n_5991 ,csa_tree_add_51_79_groupi_n_3761 ,csa_tree_add_51_79_groupi_n_5155);
  or csa_tree_add_51_79_groupi_g40098(csa_tree_add_51_79_groupi_n_5990 ,csa_tree_add_51_79_groupi_n_4996 ,csa_tree_add_51_79_groupi_n_5196);
  and csa_tree_add_51_79_groupi_g40099(csa_tree_add_51_79_groupi_n_5989 ,csa_tree_add_51_79_groupi_n_5188 ,csa_tree_add_51_79_groupi_n_5183);
  or csa_tree_add_51_79_groupi_g40100(csa_tree_add_51_79_groupi_n_5988 ,csa_tree_add_51_79_groupi_n_4993 ,csa_tree_add_51_79_groupi_n_5176);
  nor csa_tree_add_51_79_groupi_g40101(csa_tree_add_51_79_groupi_n_5987 ,csa_tree_add_51_79_groupi_n_3783 ,csa_tree_add_51_79_groupi_n_5398);
  and csa_tree_add_51_79_groupi_g40102(csa_tree_add_51_79_groupi_n_5986 ,csa_tree_add_51_79_groupi_n_4993 ,csa_tree_add_51_79_groupi_n_5176);
  or csa_tree_add_51_79_groupi_g40103(csa_tree_add_51_79_groupi_n_5985 ,csa_tree_add_51_79_groupi_n_5174 ,csa_tree_add_51_79_groupi_n_5172);
  nor csa_tree_add_51_79_groupi_g40104(csa_tree_add_51_79_groupi_n_5984 ,csa_tree_add_51_79_groupi_n_5258 ,csa_tree_add_51_79_groupi_n_5255);
  and csa_tree_add_51_79_groupi_g40105(csa_tree_add_51_79_groupi_n_5983 ,csa_tree_add_51_79_groupi_n_5174 ,csa_tree_add_51_79_groupi_n_5172);
  or csa_tree_add_51_79_groupi_g40106(csa_tree_add_51_79_groupi_n_5982 ,csa_tree_add_51_79_groupi_n_4995 ,csa_tree_add_51_79_groupi_n_5157);
  and csa_tree_add_51_79_groupi_g40107(csa_tree_add_51_79_groupi_n_5981 ,csa_tree_add_51_79_groupi_n_4995 ,csa_tree_add_51_79_groupi_n_5157);
  or csa_tree_add_51_79_groupi_g40108(csa_tree_add_51_79_groupi_n_5980 ,csa_tree_add_51_79_groupi_n_5325 ,csa_tree_add_51_79_groupi_n_5430);
  or csa_tree_add_51_79_groupi_g40109(csa_tree_add_51_79_groupi_n_5979 ,csa_tree_add_51_79_groupi_n_4960 ,csa_tree_add_51_79_groupi_n_5261);
  nor csa_tree_add_51_79_groupi_g40110(csa_tree_add_51_79_groupi_n_5978 ,csa_tree_add_51_79_groupi_n_3775 ,csa_tree_add_51_79_groupi_n_4827);
  and csa_tree_add_51_79_groupi_g40111(csa_tree_add_51_79_groupi_n_5977 ,csa_tree_add_51_79_groupi_n_5325 ,csa_tree_add_51_79_groupi_n_5430);
  or csa_tree_add_51_79_groupi_g40112(csa_tree_add_51_79_groupi_n_5976 ,csa_tree_add_51_79_groupi_n_5252 ,csa_tree_add_51_79_groupi_n_5262);
  and csa_tree_add_51_79_groupi_g40113(csa_tree_add_51_79_groupi_n_5975 ,csa_tree_add_51_79_groupi_n_4986 ,csa_tree_add_51_79_groupi_n_5161);
  or csa_tree_add_51_79_groupi_g40114(csa_tree_add_51_79_groupi_n_5974 ,csa_tree_add_51_79_groupi_n_4937 ,csa_tree_add_51_79_groupi_n_5177);
  and csa_tree_add_51_79_groupi_g40115(csa_tree_add_51_79_groupi_n_5973 ,csa_tree_add_51_79_groupi_n_5272 ,csa_tree_add_51_79_groupi_n_5397);
  or csa_tree_add_51_79_groupi_g40116(csa_tree_add_51_79_groupi_n_5972 ,csa_tree_add_51_79_groupi_n_3782 ,csa_tree_add_51_79_groupi_n_5399);
  and csa_tree_add_51_79_groupi_g40117(csa_tree_add_51_79_groupi_n_5971 ,csa_tree_add_51_79_groupi_n_4991 ,csa_tree_add_51_79_groupi_n_5269);
  nor csa_tree_add_51_79_groupi_g40118(csa_tree_add_51_79_groupi_n_5970 ,csa_tree_add_51_79_groupi_n_3762 ,csa_tree_add_51_79_groupi_n_5154);
  or csa_tree_add_51_79_groupi_g40119(csa_tree_add_51_79_groupi_n_5969 ,csa_tree_add_51_79_groupi_n_4921 ,csa_tree_add_51_79_groupi_n_5327);
  or csa_tree_add_51_79_groupi_g40120(csa_tree_add_51_79_groupi_n_5968 ,csa_tree_add_51_79_groupi_n_3228 ,csa_tree_add_51_79_groupi_n_5416);
  nor csa_tree_add_51_79_groupi_g40121(csa_tree_add_51_79_groupi_n_5967 ,csa_tree_add_51_79_groupi_n_4895 ,csa_tree_add_51_79_groupi_n_5418);
  and csa_tree_add_51_79_groupi_g40122(csa_tree_add_51_79_groupi_n_5966 ,csa_tree_add_51_79_groupi_n_4895 ,csa_tree_add_51_79_groupi_n_5418);
  or csa_tree_add_51_79_groupi_g40123(csa_tree_add_51_79_groupi_n_5965 ,csa_tree_add_51_79_groupi_n_5408 ,csa_tree_add_51_79_groupi_n_5407);
  or csa_tree_add_51_79_groupi_g40124(csa_tree_add_51_79_groupi_n_5964 ,csa_tree_add_51_79_groupi_n_4974 ,csa_tree_add_51_79_groupi_n_4842);
  or csa_tree_add_51_79_groupi_g40125(csa_tree_add_51_79_groupi_n_5963 ,csa_tree_add_51_79_groupi_n_3807 ,csa_tree_add_51_79_groupi_n_5360);
  or csa_tree_add_51_79_groupi_g40126(csa_tree_add_51_79_groupi_n_5962 ,csa_tree_add_51_79_groupi_n_5188 ,csa_tree_add_51_79_groupi_n_5183);
  nor csa_tree_add_51_79_groupi_g40127(csa_tree_add_51_79_groupi_n_5961 ,csa_tree_add_51_79_groupi_n_3229 ,csa_tree_add_51_79_groupi_n_5415);
  and csa_tree_add_51_79_groupi_g40128(csa_tree_add_51_79_groupi_n_5960 ,csa_tree_add_51_79_groupi_n_4813 ,csa_tree_add_51_79_groupi_n_5187);
  or csa_tree_add_51_79_groupi_g40129(csa_tree_add_51_79_groupi_n_5959 ,csa_tree_add_51_79_groupi_n_3308 ,csa_tree_add_51_79_groupi_n_5423);
  or csa_tree_add_51_79_groupi_g40130(csa_tree_add_51_79_groupi_n_5958 ,csa_tree_add_51_79_groupi_n_3774 ,csa_tree_add_51_79_groupi_n_4828);
  nor csa_tree_add_51_79_groupi_g40131(csa_tree_add_51_79_groupi_n_5957 ,csa_tree_add_51_79_groupi_n_3309 ,csa_tree_add_51_79_groupi_n_5422);
  or csa_tree_add_51_79_groupi_g40132(csa_tree_add_51_79_groupi_n_5956 ,csa_tree_add_51_79_groupi_n_3745 ,csa_tree_add_51_79_groupi_n_5388);
  nor csa_tree_add_51_79_groupi_g40133(csa_tree_add_51_79_groupi_n_5955 ,csa_tree_add_51_79_groupi_n_3746 ,csa_tree_add_51_79_groupi_n_5387);
  or csa_tree_add_51_79_groupi_g40134(csa_tree_add_51_79_groupi_n_5954 ,csa_tree_add_51_79_groupi_n_4988 ,csa_tree_add_51_79_groupi_n_4840);
  or csa_tree_add_51_79_groupi_g40135(csa_tree_add_51_79_groupi_n_5953 ,csa_tree_add_51_79_groupi_n_3752 ,csa_tree_add_51_79_groupi_n_5265);
  nor csa_tree_add_51_79_groupi_g40136(csa_tree_add_51_79_groupi_n_5952 ,csa_tree_add_51_79_groupi_n_4989 ,csa_tree_add_51_79_groupi_n_4839);
  or csa_tree_add_51_79_groupi_g40137(csa_tree_add_51_79_groupi_n_5951 ,csa_tree_add_51_79_groupi_n_3824 ,csa_tree_add_51_79_groupi_n_5381);
  and csa_tree_add_51_79_groupi_g40138(csa_tree_add_51_79_groupi_n_5950 ,csa_tree_add_51_79_groupi_n_4984 ,csa_tree_add_51_79_groupi_n_5383);
  or csa_tree_add_51_79_groupi_g40139(csa_tree_add_51_79_groupi_n_5949 ,csa_tree_add_51_79_groupi_n_4983 ,csa_tree_add_51_79_groupi_n_5379);
  nor csa_tree_add_51_79_groupi_g40140(csa_tree_add_51_79_groupi_n_5948 ,csa_tree_add_51_79_groupi_n_3751 ,csa_tree_add_51_79_groupi_n_5266);
  or csa_tree_add_51_79_groupi_g40141(csa_tree_add_51_79_groupi_n_5947 ,csa_tree_add_51_79_groupi_n_4361 ,csa_tree_add_51_79_groupi_n_5509);
  and csa_tree_add_51_79_groupi_g40142(csa_tree_add_51_79_groupi_n_5946 ,csa_tree_add_51_79_groupi_n_4983 ,csa_tree_add_51_79_groupi_n_5379);
  or csa_tree_add_51_79_groupi_g40143(csa_tree_add_51_79_groupi_n_5945 ,csa_tree_add_51_79_groupi_n_5319 ,csa_tree_add_51_79_groupi_n_5373);
  and csa_tree_add_51_79_groupi_g40144(csa_tree_add_51_79_groupi_n_5944 ,csa_tree_add_51_79_groupi_n_4916 ,csa_tree_add_51_79_groupi_n_5192);
  nor csa_tree_add_51_79_groupi_g40145(csa_tree_add_51_79_groupi_n_5943 ,csa_tree_add_51_79_groupi_n_3825 ,csa_tree_add_51_79_groupi_n_5380);
  nor csa_tree_add_51_79_groupi_g40146(csa_tree_add_51_79_groupi_n_5942 ,csa_tree_add_51_79_groupi_n_5372 ,csa_tree_add_51_79_groupi_n_5370);
  and csa_tree_add_51_79_groupi_g40147(csa_tree_add_51_79_groupi_n_5941 ,csa_tree_add_51_79_groupi_n_5319 ,csa_tree_add_51_79_groupi_n_5373);
  or csa_tree_add_51_79_groupi_g40148(csa_tree_add_51_79_groupi_n_5940 ,csa_tree_add_51_79_groupi_n_5349 ,csa_tree_add_51_79_groupi_n_5368);
  or csa_tree_add_51_79_groupi_g40149(csa_tree_add_51_79_groupi_n_5939 ,csa_tree_add_51_79_groupi_n_3779 ,csa_tree_add_51_79_groupi_n_5367);
  and csa_tree_add_51_79_groupi_g40150(csa_tree_add_51_79_groupi_n_5938 ,csa_tree_add_51_79_groupi_n_5349 ,csa_tree_add_51_79_groupi_n_5368);
  or csa_tree_add_51_79_groupi_g40151(csa_tree_add_51_79_groupi_n_5937 ,csa_tree_add_51_79_groupi_n_4979 ,csa_tree_add_51_79_groupi_n_5365);
  or csa_tree_add_51_79_groupi_g40152(csa_tree_add_51_79_groupi_n_5936 ,csa_tree_add_51_79_groupi_n_3811 ,csa_tree_add_51_79_groupi_n_5352);
  or csa_tree_add_51_79_groupi_g40153(csa_tree_add_51_79_groupi_n_5935 ,csa_tree_add_51_79_groupi_n_5371 ,csa_tree_add_51_79_groupi_n_5369);
  or csa_tree_add_51_79_groupi_g40154(csa_tree_add_51_79_groupi_n_5934 ,csa_tree_add_51_79_groupi_n_4853 ,csa_tree_add_51_79_groupi_n_5357);
  and csa_tree_add_51_79_groupi_g40155(csa_tree_add_51_79_groupi_n_5933 ,csa_tree_add_51_79_groupi_n_4979 ,csa_tree_add_51_79_groupi_n_5365);
  or csa_tree_add_51_79_groupi_g40156(csa_tree_add_51_79_groupi_n_5932 ,csa_tree_add_51_79_groupi_n_5361 ,csa_tree_add_51_79_groupi_n_5358);
  and csa_tree_add_51_79_groupi_g40157(csa_tree_add_51_79_groupi_n_5931 ,csa_tree_add_51_79_groupi_n_5361 ,csa_tree_add_51_79_groupi_n_5358);
  or csa_tree_add_51_79_groupi_g40158(csa_tree_add_51_79_groupi_n_5930 ,csa_tree_add_51_79_groupi_n_4901 ,csa_tree_add_51_79_groupi_n_5353);
  nor csa_tree_add_51_79_groupi_g40159(csa_tree_add_51_79_groupi_n_5929 ,csa_tree_add_51_79_groupi_n_3780 ,csa_tree_add_51_79_groupi_n_5366);
  and csa_tree_add_51_79_groupi_g40160(csa_tree_add_51_79_groupi_n_5928 ,csa_tree_add_51_79_groupi_n_4853 ,csa_tree_add_51_79_groupi_n_5357);
  or csa_tree_add_51_79_groupi_g40161(csa_tree_add_51_79_groupi_n_5927 ,csa_tree_add_51_79_groupi_n_3802 ,csa_tree_add_51_79_groupi_n_5160);
  nor csa_tree_add_51_79_groupi_g40162(csa_tree_add_51_79_groupi_n_5926 ,csa_tree_add_51_79_groupi_n_3757 ,csa_tree_add_51_79_groupi_n_5179);
  nor csa_tree_add_51_79_groupi_g40163(csa_tree_add_51_79_groupi_n_5925 ,csa_tree_add_51_79_groupi_n_3227 ,csa_tree_add_51_79_groupi_n_4823);
  nor csa_tree_add_51_79_groupi_g40164(csa_tree_add_51_79_groupi_n_5924 ,csa_tree_add_51_79_groupi_n_3803 ,csa_tree_add_51_79_groupi_n_5159);
  or csa_tree_add_51_79_groupi_g40165(csa_tree_add_51_79_groupi_n_5923 ,csa_tree_add_51_79_groupi_n_4945 ,csa_tree_add_51_79_groupi_n_5343);
  or csa_tree_add_51_79_groupi_g40166(csa_tree_add_51_79_groupi_n_5922 ,csa_tree_add_51_79_groupi_n_4843 ,csa_tree_add_51_79_groupi_n_5217);
  and csa_tree_add_51_79_groupi_g40167(csa_tree_add_51_79_groupi_n_5921 ,csa_tree_add_51_79_groupi_n_4797 ,csa_tree_add_51_79_groupi_n_5350);
  and csa_tree_add_51_79_groupi_g40168(csa_tree_add_51_79_groupi_n_5920 ,csa_tree_add_51_79_groupi_n_4799 ,csa_tree_add_51_79_groupi_n_4801);
  nor csa_tree_add_51_79_groupi_g40169(csa_tree_add_51_79_groupi_n_5919 ,csa_tree_add_51_79_groupi_n_4946 ,csa_tree_add_51_79_groupi_n_5342);
  or csa_tree_add_51_79_groupi_g40170(csa_tree_add_51_79_groupi_n_5918 ,csa_tree_add_51_79_groupi_n_4990 ,csa_tree_add_51_79_groupi_n_5158);
  and csa_tree_add_51_79_groupi_g40171(csa_tree_add_51_79_groupi_n_5917 ,csa_tree_add_51_79_groupi_n_5238 ,csa_tree_add_51_79_groupi_n_5232);
  and csa_tree_add_51_79_groupi_g40172(csa_tree_add_51_79_groupi_n_5916 ,csa_tree_add_51_79_groupi_n_5007 ,csa_tree_add_51_79_groupi_n_5414);
  or csa_tree_add_51_79_groupi_g40173(csa_tree_add_51_79_groupi_n_5915 ,csa_tree_add_51_79_groupi_n_5270 ,csa_tree_add_51_79_groupi_n_5395);
  nor csa_tree_add_51_79_groupi_g40174(csa_tree_add_51_79_groupi_n_5914 ,csa_tree_add_51_79_groupi_n_3820 ,csa_tree_add_51_79_groupi_n_5337);
  or csa_tree_add_51_79_groupi_g40175(csa_tree_add_51_79_groupi_n_5913 ,csa_tree_add_51_79_groupi_n_5272 ,csa_tree_add_51_79_groupi_n_5397);
  nor csa_tree_add_51_79_groupi_g40176(csa_tree_add_51_79_groupi_n_5912 ,csa_tree_add_51_79_groupi_n_3808 ,csa_tree_add_51_79_groupi_n_5359);
  or csa_tree_add_51_79_groupi_g40177(csa_tree_add_51_79_groupi_n_5911 ,csa_tree_add_51_79_groupi_n_4900 ,csa_tree_add_51_79_groupi_n_5333);
  or csa_tree_add_51_79_groupi_g40178(csa_tree_add_51_79_groupi_n_5910 ,csa_tree_add_51_79_groupi_n_3821 ,csa_tree_add_51_79_groupi_n_5336);
  nor csa_tree_add_51_79_groupi_g40179(csa_tree_add_51_79_groupi_n_5909 ,csa_tree_add_51_79_groupi_n_3812 ,csa_tree_add_51_79_groupi_n_5351);
  nor csa_tree_add_51_79_groupi_g40180(csa_tree_add_51_79_groupi_n_5908 ,csa_tree_add_51_79_groupi_n_3817 ,csa_tree_add_51_79_groupi_n_5210);
  and csa_tree_add_51_79_groupi_g40181(csa_tree_add_51_79_groupi_n_5907 ,csa_tree_add_51_79_groupi_n_4975 ,csa_tree_add_51_79_groupi_n_5330);
  or csa_tree_add_51_79_groupi_g40182(csa_tree_add_51_79_groupi_n_5906 ,csa_tree_add_51_79_groupi_n_5189 ,csa_tree_add_51_79_groupi_n_5328);
  and csa_tree_add_51_79_groupi_g40183(csa_tree_add_51_79_groupi_n_5905 ,csa_tree_add_51_79_groupi_n_3290 ,csa_tree_add_51_79_groupi_n_5250);
  and csa_tree_add_51_79_groupi_g40184(csa_tree_add_51_79_groupi_n_5904 ,csa_tree_add_51_79_groupi_n_5189 ,csa_tree_add_51_79_groupi_n_5328);
  and csa_tree_add_51_79_groupi_g40185(csa_tree_add_51_79_groupi_n_5903 ,csa_tree_add_51_79_groupi_n_4900 ,csa_tree_add_51_79_groupi_n_5333);
  nor csa_tree_add_51_79_groupi_g40186(csa_tree_add_51_79_groupi_n_5902 ,csa_tree_add_51_79_groupi_n_4964 ,csa_tree_add_51_79_groupi_n_5280);
  or csa_tree_add_51_79_groupi_g40187(csa_tree_add_51_79_groupi_n_5901 ,csa_tree_add_51_79_groupi_n_3733 ,csa_tree_add_51_79_groupi_n_5268);
  or csa_tree_add_51_79_groupi_g40188(csa_tree_add_51_79_groupi_n_5900 ,csa_tree_add_51_79_groupi_n_4938 ,csa_tree_add_51_79_groupi_n_5412);
  nor csa_tree_add_51_79_groupi_g40189(csa_tree_add_51_79_groupi_n_5899 ,csa_tree_add_51_79_groupi_n_3734 ,csa_tree_add_51_79_groupi_n_5267);
  nor csa_tree_add_51_79_groupi_g40190(csa_tree_add_51_79_groupi_n_5898 ,csa_tree_add_51_79_groupi_n_3215 ,csa_tree_add_51_79_groupi_n_5402);
  and csa_tree_add_51_79_groupi_g40191(csa_tree_add_51_79_groupi_n_5897 ,csa_tree_add_51_79_groupi_n_5285 ,csa_tree_add_51_79_groupi_n_5284);
  or csa_tree_add_51_79_groupi_g40192(csa_tree_add_51_79_groupi_n_5896 ,csa_tree_add_51_79_groupi_n_2570 ,csa_tree_add_51_79_groupi_n_4790);
  or csa_tree_add_51_79_groupi_g40193(csa_tree_add_51_79_groupi_n_5895 ,csa_tree_add_51_79_groupi_n_3295 ,csa_tree_add_51_79_groupi_n_5237);
  or csa_tree_add_51_79_groupi_g40194(csa_tree_add_51_79_groupi_n_5894 ,csa_tree_add_51_79_groupi_n_4971 ,csa_tree_add_51_79_groupi_n_5311);
  or csa_tree_add_51_79_groupi_g40195(csa_tree_add_51_79_groupi_n_5893 ,csa_tree_add_51_79_groupi_n_4963 ,csa_tree_add_51_79_groupi_n_5281);
  and csa_tree_add_51_79_groupi_g40196(csa_tree_add_51_79_groupi_n_5892 ,csa_tree_add_51_79_groupi_n_4971 ,csa_tree_add_51_79_groupi_n_5311);
  or csa_tree_add_51_79_groupi_g40197(csa_tree_add_51_79_groupi_n_5891 ,csa_tree_add_51_79_groupi_n_5264 ,csa_tree_add_51_79_groupi_n_5310);
  and csa_tree_add_51_79_groupi_g40198(csa_tree_add_51_79_groupi_n_5890 ,csa_tree_add_51_79_groupi_n_5264 ,csa_tree_add_51_79_groupi_n_5310);
  nor csa_tree_add_51_79_groupi_g40199(csa_tree_add_51_79_groupi_n_5889 ,csa_tree_add_51_79_groupi_n_3235 ,csa_tree_add_51_79_groupi_n_5322);
  or csa_tree_add_51_79_groupi_g40200(csa_tree_add_51_79_groupi_n_5888 ,csa_tree_add_51_79_groupi_n_3214 ,csa_tree_add_51_79_groupi_n_5403);
  and csa_tree_add_51_79_groupi_g40201(csa_tree_add_51_79_groupi_n_5887 ,csa_tree_add_51_79_groupi_n_4965 ,csa_tree_add_51_79_groupi_n_5290);
  or csa_tree_add_51_79_groupi_g40202(csa_tree_add_51_79_groupi_n_5886 ,csa_tree_add_51_79_groupi_n_4965 ,csa_tree_add_51_79_groupi_n_5290);
  or csa_tree_add_51_79_groupi_g40203(csa_tree_add_51_79_groupi_n_5885 ,csa_tree_add_51_79_groupi_n_3759 ,csa_tree_add_51_79_groupi_n_5306);
  or csa_tree_add_51_79_groupi_g40204(csa_tree_add_51_79_groupi_n_5884 ,csa_tree_add_51_79_groupi_n_5307 ,csa_tree_add_51_79_groupi_n_5304);
  and csa_tree_add_51_79_groupi_g40205(csa_tree_add_51_79_groupi_n_5883 ,csa_tree_add_51_79_groupi_n_5307 ,csa_tree_add_51_79_groupi_n_5304);
  or csa_tree_add_51_79_groupi_g40206(csa_tree_add_51_79_groupi_n_5882 ,csa_tree_add_51_79_groupi_n_4967 ,csa_tree_add_51_79_groupi_n_5297);
  or csa_tree_add_51_79_groupi_g40207(csa_tree_add_51_79_groupi_n_5881 ,csa_tree_add_51_79_groupi_n_4969 ,csa_tree_add_51_79_groupi_n_5298);
  nor csa_tree_add_51_79_groupi_g40208(csa_tree_add_51_79_groupi_n_5880 ,csa_tree_add_51_79_groupi_n_3760 ,csa_tree_add_51_79_groupi_n_5305);
  or csa_tree_add_51_79_groupi_g40209(csa_tree_add_51_79_groupi_n_5879 ,csa_tree_add_51_79_groupi_n_4973 ,csa_tree_add_51_79_groupi_n_5164);
  or csa_tree_add_51_79_groupi_g40210(csa_tree_add_51_79_groupi_n_5878 ,csa_tree_add_51_79_groupi_n_5295 ,csa_tree_add_51_79_groupi_n_5294);
  or csa_tree_add_51_79_groupi_g40211(csa_tree_add_51_79_groupi_n_5877 ,csa_tree_add_51_79_groupi_n_4918 ,csa_tree_add_51_79_groupi_n_5209);
  nor csa_tree_add_51_79_groupi_g40212(csa_tree_add_51_79_groupi_n_5876 ,csa_tree_add_51_79_groupi_n_3302 ,csa_tree_add_51_79_groupi_n_5228);
  or csa_tree_add_51_79_groupi_g40213(csa_tree_add_51_79_groupi_n_5875 ,csa_tree_add_51_79_groupi_n_4994 ,csa_tree_add_51_79_groupi_n_4802);
  nor csa_tree_add_51_79_groupi_g40214(csa_tree_add_51_79_groupi_n_5874 ,csa_tree_add_51_79_groupi_n_4968 ,csa_tree_add_51_79_groupi_n_5296);
  nor csa_tree_add_51_79_groupi_g40215(csa_tree_add_51_79_groupi_n_5873 ,csa_tree_add_51_79_groupi_n_3296 ,csa_tree_add_51_79_groupi_n_5236);
  nor csa_tree_add_51_79_groupi_g40216(csa_tree_add_51_79_groupi_n_5872 ,csa_tree_add_51_79_groupi_n_3271 ,csa_tree_add_51_79_groupi_n_5292);
  and csa_tree_add_51_79_groupi_g40217(csa_tree_add_51_79_groupi_n_5871 ,csa_tree_add_51_79_groupi_n_5295 ,csa_tree_add_51_79_groupi_n_5294);
  and csa_tree_add_51_79_groupi_g40218(csa_tree_add_51_79_groupi_n_5870 ,csa_tree_add_51_79_groupi_n_1210 ,csa_tree_add_51_79_groupi_n_763);
  or csa_tree_add_51_79_groupi_g40219(csa_tree_add_51_79_groupi_n_5869 ,csa_tree_add_51_79_groupi_n_1210 ,csa_tree_add_51_79_groupi_n_11);
  or csa_tree_add_51_79_groupi_g40220(csa_tree_add_51_79_groupi_n_6156 ,csa_tree_add_51_79_groupi_n_4304 ,csa_tree_add_51_79_groupi_n_5135);
  and csa_tree_add_51_79_groupi_g40221(csa_tree_add_51_79_groupi_n_6155 ,csa_tree_add_51_79_groupi_n_4478 ,csa_tree_add_51_79_groupi_n_5143);
  and csa_tree_add_51_79_groupi_g40222(csa_tree_add_51_79_groupi_n_6154 ,csa_tree_add_51_79_groupi_n_4136 ,csa_tree_add_51_79_groupi_n_5142);
  or csa_tree_add_51_79_groupi_g40223(csa_tree_add_51_79_groupi_n_6153 ,csa_tree_add_51_79_groupi_n_5463 ,csa_tree_add_51_79_groupi_n_5454);
  and csa_tree_add_51_79_groupi_g40224(csa_tree_add_51_79_groupi_n_6152 ,csa_tree_add_51_79_groupi_n_4396 ,csa_tree_add_51_79_groupi_n_4788);
  or csa_tree_add_51_79_groupi_g40225(csa_tree_add_51_79_groupi_n_6151 ,csa_tree_add_51_79_groupi_n_3320 ,csa_tree_add_51_79_groupi_n_5107);
  or csa_tree_add_51_79_groupi_g40226(csa_tree_add_51_79_groupi_n_6150 ,csa_tree_add_51_79_groupi_n_3829 ,csa_tree_add_51_79_groupi_n_5434);
  and csa_tree_add_51_79_groupi_g40227(csa_tree_add_51_79_groupi_n_6149 ,csa_tree_add_51_79_groupi_n_4117 ,csa_tree_add_51_79_groupi_n_5132);
  and csa_tree_add_51_79_groupi_g40228(csa_tree_add_51_79_groupi_n_6148 ,csa_tree_add_51_79_groupi_n_4698 ,csa_tree_add_51_79_groupi_n_5152);
  and csa_tree_add_51_79_groupi_g40229(csa_tree_add_51_79_groupi_n_6147 ,csa_tree_add_51_79_groupi_n_4365 ,csa_tree_add_51_79_groupi_n_5138);
  or csa_tree_add_51_79_groupi_g40230(csa_tree_add_51_79_groupi_n_6146 ,csa_tree_add_51_79_groupi_n_4712 ,csa_tree_add_51_79_groupi_n_5139);
  or csa_tree_add_51_79_groupi_g40231(csa_tree_add_51_79_groupi_n_6145 ,csa_tree_add_51_79_groupi_n_4305 ,csa_tree_add_51_79_groupi_n_5140);
  and csa_tree_add_51_79_groupi_g40232(csa_tree_add_51_79_groupi_n_6144 ,csa_tree_add_51_79_groupi_n_4483 ,csa_tree_add_51_79_groupi_n_5145);
  and csa_tree_add_51_79_groupi_g40233(csa_tree_add_51_79_groupi_n_6143 ,csa_tree_add_51_79_groupi_n_5518 ,csa_tree_add_51_79_groupi_n_5097);
  and csa_tree_add_51_79_groupi_g40234(csa_tree_add_51_79_groupi_n_6141 ,csa_tree_add_51_79_groupi_n_4456 ,csa_tree_add_51_79_groupi_n_5130);
  and csa_tree_add_51_79_groupi_g40235(csa_tree_add_51_79_groupi_n_6140 ,csa_tree_add_51_79_groupi_n_4045 ,csa_tree_add_51_79_groupi_n_5133);
  and csa_tree_add_51_79_groupi_g40236(csa_tree_add_51_79_groupi_n_6139 ,csa_tree_add_51_79_groupi_n_5035 ,csa_tree_add_51_79_groupi_n_5444);
  and csa_tree_add_51_79_groupi_g40237(csa_tree_add_51_79_groupi_n_6138 ,csa_tree_add_51_79_groupi_n_4687 ,csa_tree_add_51_79_groupi_n_5144);
  and csa_tree_add_51_79_groupi_g40238(csa_tree_add_51_79_groupi_n_6137 ,csa_tree_add_51_79_groupi_n_4367 ,csa_tree_add_51_79_groupi_n_5137);
  or csa_tree_add_51_79_groupi_g40239(csa_tree_add_51_79_groupi_n_6136 ,csa_tree_add_51_79_groupi_n_4554 ,csa_tree_add_51_79_groupi_n_5146);
  or csa_tree_add_51_79_groupi_g40240(csa_tree_add_51_79_groupi_n_6134 ,csa_tree_add_51_79_groupi_n_4352 ,csa_tree_add_51_79_groupi_n_5150);
  and csa_tree_add_51_79_groupi_g40241(csa_tree_add_51_79_groupi_n_6132 ,csa_tree_add_51_79_groupi_n_4668 ,csa_tree_add_51_79_groupi_n_5127);
  or csa_tree_add_51_79_groupi_g40242(csa_tree_add_51_79_groupi_n_6131 ,csa_tree_add_51_79_groupi_n_4640 ,csa_tree_add_51_79_groupi_n_5149);
  and csa_tree_add_51_79_groupi_g40243(csa_tree_add_51_79_groupi_n_6129 ,csa_tree_add_51_79_groupi_n_4390 ,csa_tree_add_51_79_groupi_n_4771);
  or csa_tree_add_51_79_groupi_g40244(csa_tree_add_51_79_groupi_n_6128 ,csa_tree_add_51_79_groupi_n_4058 ,csa_tree_add_51_79_groupi_n_5151);
  or csa_tree_add_51_79_groupi_g40245(csa_tree_add_51_79_groupi_n_6127 ,csa_tree_add_51_79_groupi_n_4447 ,csa_tree_add_51_79_groupi_n_5131);
  not csa_tree_add_51_79_groupi_g40246(csa_tree_add_51_79_groupi_n_5862 ,csa_tree_add_51_79_groupi_n_5861);
  not csa_tree_add_51_79_groupi_g40247(csa_tree_add_51_79_groupi_n_5857 ,csa_tree_add_51_79_groupi_n_5858);
  not csa_tree_add_51_79_groupi_g40248(csa_tree_add_51_79_groupi_n_5855 ,csa_tree_add_51_79_groupi_n_5856);
  not csa_tree_add_51_79_groupi_g40250(csa_tree_add_51_79_groupi_n_5852 ,csa_tree_add_51_79_groupi_n_5853);
  not csa_tree_add_51_79_groupi_g40251(csa_tree_add_51_79_groupi_n_5847 ,csa_tree_add_51_79_groupi_n_5848);
  not csa_tree_add_51_79_groupi_g40252(csa_tree_add_51_79_groupi_n_5843 ,csa_tree_add_51_79_groupi_n_5844);
  not csa_tree_add_51_79_groupi_g40253(csa_tree_add_51_79_groupi_n_5840 ,csa_tree_add_51_79_groupi_n_5841);
  and csa_tree_add_51_79_groupi_g40254(csa_tree_add_51_79_groupi_n_5839 ,csa_tree_add_51_79_groupi_n_4893 ,csa_tree_add_51_79_groupi_n_4848);
  or csa_tree_add_51_79_groupi_g40255(csa_tree_add_51_79_groupi_n_5838 ,csa_tree_add_51_79_groupi_n_5182 ,csa_tree_add_51_79_groupi_n_5393);
  or csa_tree_add_51_79_groupi_g40256(csa_tree_add_51_79_groupi_n_5837 ,csa_tree_add_51_79_groupi_n_3770 ,csa_tree_add_51_79_groupi_n_5241);
  and csa_tree_add_51_79_groupi_g40257(csa_tree_add_51_79_groupi_n_5836 ,csa_tree_add_51_79_groupi_n_5182 ,csa_tree_add_51_79_groupi_n_5393);
  and csa_tree_add_51_79_groupi_g40258(csa_tree_add_51_79_groupi_n_5835 ,csa_tree_add_51_79_groupi_n_4955 ,csa_tree_add_51_79_groupi_n_5239);
  nor csa_tree_add_51_79_groupi_g40259(csa_tree_add_51_79_groupi_n_5834 ,csa_tree_add_51_79_groupi_n_3771 ,csa_tree_add_51_79_groupi_n_5240);
  or csa_tree_add_51_79_groupi_g40260(csa_tree_add_51_79_groupi_n_5833 ,csa_tree_add_51_79_groupi_n_5234 ,csa_tree_add_51_79_groupi_n_5231);
  and csa_tree_add_51_79_groupi_g40261(csa_tree_add_51_79_groupi_n_5832 ,csa_tree_add_51_79_groupi_n_3741 ,csa_tree_add_51_79_groupi_n_5242);
  or csa_tree_add_51_79_groupi_g40262(csa_tree_add_51_79_groupi_n_5831 ,csa_tree_add_51_79_groupi_n_3301 ,csa_tree_add_51_79_groupi_n_5229);
  or csa_tree_add_51_79_groupi_g40263(csa_tree_add_51_79_groupi_n_5830 ,csa_tree_add_51_79_groupi_n_5233 ,csa_tree_add_51_79_groupi_n_5230);
  and csa_tree_add_51_79_groupi_g40264(csa_tree_add_51_79_groupi_n_5829 ,csa_tree_add_51_79_groupi_n_5233 ,csa_tree_add_51_79_groupi_n_5230);
  and csa_tree_add_51_79_groupi_g40265(csa_tree_add_51_79_groupi_n_5828 ,csa_tree_add_51_79_groupi_n_5234 ,csa_tree_add_51_79_groupi_n_5231);
  or csa_tree_add_51_79_groupi_g40266(csa_tree_add_51_79_groupi_n_5827 ,csa_tree_add_51_79_groupi_n_5227 ,csa_tree_add_51_79_groupi_n_5225);
  and csa_tree_add_51_79_groupi_g40267(csa_tree_add_51_79_groupi_n_5826 ,csa_tree_add_51_79_groupi_n_4952 ,csa_tree_add_51_79_groupi_n_5226);
  or csa_tree_add_51_79_groupi_g40268(csa_tree_add_51_79_groupi_n_5825 ,csa_tree_add_51_79_groupi_n_5223 ,csa_tree_add_51_79_groupi_n_5222);
  and csa_tree_add_51_79_groupi_g40269(csa_tree_add_51_79_groupi_n_5824 ,csa_tree_add_51_79_groupi_n_5223 ,csa_tree_add_51_79_groupi_n_5222);
  and csa_tree_add_51_79_groupi_g40270(csa_tree_add_51_79_groupi_n_5823 ,csa_tree_add_51_79_groupi_n_5227 ,csa_tree_add_51_79_groupi_n_5225);
  or csa_tree_add_51_79_groupi_g40271(csa_tree_add_51_79_groupi_n_5822 ,csa_tree_add_51_79_groupi_n_5220 ,csa_tree_add_51_79_groupi_n_5219);
  and csa_tree_add_51_79_groupi_g40272(csa_tree_add_51_79_groupi_n_5821 ,csa_tree_add_51_79_groupi_n_4994 ,csa_tree_add_51_79_groupi_n_4802);
  or csa_tree_add_51_79_groupi_g40273(csa_tree_add_51_79_groupi_n_5820 ,csa_tree_add_51_79_groupi_n_4944 ,csa_tree_add_51_79_groupi_n_5420);
  or csa_tree_add_51_79_groupi_g40274(csa_tree_add_51_79_groupi_n_5819 ,csa_tree_add_51_79_groupi_n_3772 ,csa_tree_add_51_79_groupi_n_5275);
  and csa_tree_add_51_79_groupi_g40275(csa_tree_add_51_79_groupi_n_5818 ,csa_tree_add_51_79_groupi_n_5220 ,csa_tree_add_51_79_groupi_n_5219);
  or csa_tree_add_51_79_groupi_g40276(csa_tree_add_51_79_groupi_n_5817 ,csa_tree_add_51_79_groupi_n_4290 ,csa_tree_add_51_79_groupi_n_4780);
  or csa_tree_add_51_79_groupi_g40277(csa_tree_add_51_79_groupi_n_5816 ,csa_tree_add_51_79_groupi_n_4991 ,csa_tree_add_51_79_groupi_n_5269);
  and csa_tree_add_51_79_groupi_g40278(csa_tree_add_51_79_groupi_n_5815 ,csa_tree_add_51_79_groupi_n_4947 ,csa_tree_add_51_79_groupi_n_5212);
  or csa_tree_add_51_79_groupi_g40279(csa_tree_add_51_79_groupi_n_5814 ,csa_tree_add_51_79_groupi_n_4947 ,csa_tree_add_51_79_groupi_n_5212);
  and csa_tree_add_51_79_groupi_g40280(csa_tree_add_51_79_groupi_n_5813 ,csa_tree_add_51_79_groupi_n_5185 ,csa_tree_add_51_79_groupi_n_5199);
  and csa_tree_add_51_79_groupi_g40281(csa_tree_add_51_79_groupi_n_5812 ,csa_tree_add_51_79_groupi_n_3239 ,csa_tree_add_51_79_groupi_n_5376);
  or csa_tree_add_51_79_groupi_g40282(csa_tree_add_51_79_groupi_n_5811 ,csa_tree_add_51_79_groupi_n_4042 ,csa_tree_add_51_79_groupi_n_5441);
  nor csa_tree_add_51_79_groupi_g40283(csa_tree_add_51_79_groupi_n_5810 ,csa_tree_add_51_79_groupi_n_3232 ,csa_tree_add_51_79_groupi_n_4897);
  or csa_tree_add_51_79_groupi_g40284(csa_tree_add_51_79_groupi_n_5809 ,csa_tree_add_51_79_groupi_n_5204 ,csa_tree_add_51_79_groupi_n_5273);
  and csa_tree_add_51_79_groupi_g40285(csa_tree_add_51_79_groupi_n_5808 ,csa_tree_add_51_79_groupi_n_4938 ,csa_tree_add_51_79_groupi_n_5412);
  nor csa_tree_add_51_79_groupi_g40286(csa_tree_add_51_79_groupi_n_5807 ,csa_tree_add_51_79_groupi_n_3241 ,csa_tree_add_51_79_groupi_n_4795);
  or csa_tree_add_51_79_groupi_g40287(csa_tree_add_51_79_groupi_n_5806 ,csa_tree_add_51_79_groupi_n_5404 ,csa_tree_add_51_79_groupi_n_4838);
  and csa_tree_add_51_79_groupi_g40288(csa_tree_add_51_79_groupi_n_5805 ,csa_tree_add_51_79_groupi_n_4972 ,csa_tree_add_51_79_groupi_n_5165);
  or csa_tree_add_51_79_groupi_g40289(csa_tree_add_51_79_groupi_n_5804 ,csa_tree_add_51_79_groupi_n_3231 ,csa_tree_add_51_79_groupi_n_4896);
  and csa_tree_add_51_79_groupi_g40290(csa_tree_add_51_79_groupi_n_5803 ,csa_tree_add_51_79_groupi_n_3256 ,csa_tree_add_51_79_groupi_n_5153);
  or csa_tree_add_51_79_groupi_g40291(csa_tree_add_51_79_groupi_n_5802 ,csa_tree_add_51_79_groupi_n_4955 ,csa_tree_add_51_79_groupi_n_5239);
  or csa_tree_add_51_79_groupi_g40292(csa_tree_add_51_79_groupi_n_5801 ,csa_tree_add_51_79_groupi_n_4859 ,csa_tree_add_51_79_groupi_n_5419);
  and csa_tree_add_51_79_groupi_g40293(csa_tree_add_51_79_groupi_n_5800 ,csa_tree_add_51_79_groupi_n_5404 ,csa_tree_add_51_79_groupi_n_4838);
  or csa_tree_add_51_79_groupi_g40294(csa_tree_add_51_79_groupi_n_5799 ,csa_tree_add_51_79_groupi_n_4301 ,csa_tree_add_51_79_groupi_n_4772);
  nor csa_tree_add_51_79_groupi_g40295(csa_tree_add_51_79_groupi_n_5798 ,csa_tree_add_51_79_groupi_n_3303 ,csa_tree_add_51_79_groupi_n_4959);
  or csa_tree_add_51_79_groupi_g40296(csa_tree_add_51_79_groupi_n_5797 ,csa_tree_add_51_79_groupi_n_4948 ,csa_tree_add_51_79_groupi_n_5186);
  and csa_tree_add_51_79_groupi_g40297(csa_tree_add_51_79_groupi_n_5796 ,csa_tree_add_51_79_groupi_n_4815 ,csa_tree_add_51_79_groupi_n_4816);
  and csa_tree_add_51_79_groupi_g40298(csa_tree_add_51_79_groupi_n_5795 ,csa_tree_add_51_79_groupi_n_4948 ,csa_tree_add_51_79_groupi_n_5186);
  or csa_tree_add_51_79_groupi_g40299(csa_tree_add_51_79_groupi_n_5794 ,csa_tree_add_51_79_groupi_n_5411 ,csa_tree_add_51_79_groupi_n_4836);
  and csa_tree_add_51_79_groupi_g40300(csa_tree_add_51_79_groupi_n_5793 ,csa_tree_add_51_79_groupi_n_4981 ,csa_tree_add_51_79_groupi_n_5180);
  and csa_tree_add_51_79_groupi_g40301(csa_tree_add_51_79_groupi_n_5792 ,csa_tree_add_51_79_groupi_n_4937 ,csa_tree_add_51_79_groupi_n_5177);
  nor csa_tree_add_51_79_groupi_g40302(csa_tree_add_51_79_groupi_n_5791 ,csa_tree_add_51_79_groupi_n_3306 ,csa_tree_add_51_79_groupi_n_5163);
  or csa_tree_add_51_79_groupi_g40303(csa_tree_add_51_79_groupi_n_5790 ,csa_tree_add_51_79_groupi_n_4903 ,csa_tree_add_51_79_groupi_n_5171);
  and csa_tree_add_51_79_groupi_g40304(csa_tree_add_51_79_groupi_n_5789 ,csa_tree_add_51_79_groupi_n_4903 ,csa_tree_add_51_79_groupi_n_5171);
  and csa_tree_add_51_79_groupi_g40305(csa_tree_add_51_79_groupi_n_5788 ,csa_tree_add_51_79_groupi_n_4940 ,csa_tree_add_51_79_groupi_n_5169);
  or csa_tree_add_51_79_groupi_g40306(csa_tree_add_51_79_groupi_n_5787 ,csa_tree_add_51_79_groupi_n_4291 ,csa_tree_add_51_79_groupi_n_4779);
  or csa_tree_add_51_79_groupi_g40307(csa_tree_add_51_79_groupi_n_5786 ,csa_tree_add_51_79_groupi_n_5003 ,csa_tree_add_51_79_groupi_n_5167);
  or csa_tree_add_51_79_groupi_g40308(csa_tree_add_51_79_groupi_n_5785 ,csa_tree_add_51_79_groupi_n_3305 ,csa_tree_add_51_79_groupi_n_5162);
  nor csa_tree_add_51_79_groupi_g40309(csa_tree_add_51_79_groupi_n_5784 ,csa_tree_add_51_79_groupi_n_3197 ,csa_tree_add_51_79_groupi_n_5207);
  or csa_tree_add_51_79_groupi_g40310(csa_tree_add_51_79_groupi_n_5783 ,csa_tree_add_51_79_groupi_n_4984 ,csa_tree_add_51_79_groupi_n_5383);
  and csa_tree_add_51_79_groupi_g40311(csa_tree_add_51_79_groupi_n_5782 ,csa_tree_add_51_79_groupi_n_4935 ,csa_tree_add_51_79_groupi_n_4794);
  and csa_tree_add_51_79_groupi_g40312(csa_tree_add_51_79_groupi_n_5781 ,csa_tree_add_51_79_groupi_n_4969 ,csa_tree_add_51_79_groupi_n_5298);
  or csa_tree_add_51_79_groupi_g40313(csa_tree_add_51_79_groupi_n_5780 ,csa_tree_add_51_79_groupi_n_4940 ,csa_tree_add_51_79_groupi_n_5169);
  or csa_tree_add_51_79_groupi_g40314(csa_tree_add_51_79_groupi_n_5779 ,csa_tree_add_51_79_groupi_n_4935 ,csa_tree_add_51_79_groupi_n_4794);
  and csa_tree_add_51_79_groupi_g40315(csa_tree_add_51_79_groupi_n_5778 ,csa_tree_add_51_79_groupi_n_5197 ,csa_tree_add_51_79_groupi_n_5218);
  or csa_tree_add_51_79_groupi_g40316(csa_tree_add_51_79_groupi_n_5777 ,csa_tree_add_51_79_groupi_n_4972 ,csa_tree_add_51_79_groupi_n_5165);
  or csa_tree_add_51_79_groupi_g40317(csa_tree_add_51_79_groupi_n_5776 ,csa_tree_add_51_79_groupi_n_4952 ,csa_tree_add_51_79_groupi_n_5226);
  or csa_tree_add_51_79_groupi_g40318(csa_tree_add_51_79_groupi_n_5775 ,csa_tree_add_51_79_groupi_n_5356 ,csa_tree_add_51_79_groupi_n_4852);
  or csa_tree_add_51_79_groupi_g40319(csa_tree_add_51_79_groupi_n_5774 ,csa_tree_add_51_79_groupi_n_4293 ,csa_tree_add_51_79_groupi_n_4787);
  and csa_tree_add_51_79_groupi_g40320(csa_tree_add_51_79_groupi_n_5773 ,csa_tree_add_51_79_groupi_n_4399 ,csa_tree_add_51_79_groupi_n_5091);
  or csa_tree_add_51_79_groupi_g40321(csa_tree_add_51_79_groupi_n_5772 ,csa_tree_add_51_79_groupi_n_3818 ,csa_tree_add_51_79_groupi_n_4932);
  nor csa_tree_add_51_79_groupi_g40322(csa_tree_add_51_79_groupi_n_5771 ,csa_tree_add_51_79_groupi_n_3819 ,csa_tree_add_51_79_groupi_n_4931);
  and csa_tree_add_51_79_groupi_g40323(csa_tree_add_51_79_groupi_n_5770 ,csa_tree_add_51_79_groupi_n_5392 ,csa_tree_add_51_79_groupi_n_5320);
  and csa_tree_add_51_79_groupi_g40324(csa_tree_add_51_79_groupi_n_5769 ,csa_tree_add_51_79_groupi_n_4835 ,csa_tree_add_51_79_groupi_n_4798);
  or csa_tree_add_51_79_groupi_g40325(csa_tree_add_51_79_groupi_n_5768 ,csa_tree_add_51_79_groupi_n_4799 ,csa_tree_add_51_79_groupi_n_4801);
  or csa_tree_add_51_79_groupi_g40326(csa_tree_add_51_79_groupi_n_5767 ,csa_tree_add_51_79_groupi_n_3747 ,csa_tree_add_51_79_groupi_n_5389);
  or csa_tree_add_51_79_groupi_g40327(csa_tree_add_51_79_groupi_n_5766 ,csa_tree_add_51_79_groupi_n_4797 ,csa_tree_add_51_79_groupi_n_5350);
  or csa_tree_add_51_79_groupi_g40328(csa_tree_add_51_79_groupi_n_5765 ,csa_tree_add_51_79_groupi_n_4294 ,csa_tree_add_51_79_groupi_n_4777);
  or csa_tree_add_51_79_groupi_g40329(csa_tree_add_51_79_groupi_n_5764 ,csa_tree_add_51_79_groupi_n_5392 ,csa_tree_add_51_79_groupi_n_5320);
  and csa_tree_add_51_79_groupi_g40330(csa_tree_add_51_79_groupi_n_5763 ,csa_tree_add_51_79_groupi_n_4901 ,csa_tree_add_51_79_groupi_n_5353);
  and csa_tree_add_51_79_groupi_g40331(csa_tree_add_51_79_groupi_n_5762 ,csa_tree_add_51_79_groupi_n_4970 ,csa_tree_add_51_79_groupi_n_4808);
  or csa_tree_add_51_79_groupi_g40332(csa_tree_add_51_79_groupi_n_5761 ,csa_tree_add_51_79_groupi_n_5004 ,csa_tree_add_51_79_groupi_n_4810);
  or csa_tree_add_51_79_groupi_g40333(csa_tree_add_51_79_groupi_n_5760 ,csa_tree_add_51_79_groupi_n_4919 ,csa_tree_add_51_79_groupi_n_4812);
  and csa_tree_add_51_79_groupi_g40334(csa_tree_add_51_79_groupi_n_5759 ,csa_tree_add_51_79_groupi_n_5004 ,csa_tree_add_51_79_groupi_n_4810);
  nor csa_tree_add_51_79_groupi_g40335(csa_tree_add_51_79_groupi_n_5758 ,csa_tree_add_51_79_groupi_n_3748 ,csa_tree_add_51_79_groupi_n_5390);
  and csa_tree_add_51_79_groupi_g40336(csa_tree_add_51_79_groupi_n_5757 ,csa_tree_add_51_79_groupi_n_4919 ,csa_tree_add_51_79_groupi_n_4812);
  or csa_tree_add_51_79_groupi_g40337(csa_tree_add_51_79_groupi_n_5756 ,csa_tree_add_51_79_groupi_n_4295 ,csa_tree_add_51_79_groupi_n_4765);
  or csa_tree_add_51_79_groupi_g40338(csa_tree_add_51_79_groupi_n_5755 ,csa_tree_add_51_79_groupi_n_4090 ,csa_tree_add_51_79_groupi_n_5556);
  or csa_tree_add_51_79_groupi_g40339(csa_tree_add_51_79_groupi_n_5754 ,csa_tree_add_51_79_groupi_n_4985 ,csa_tree_add_51_79_groupi_n_4817);
  or csa_tree_add_51_79_groupi_g40340(csa_tree_add_51_79_groupi_n_5753 ,csa_tree_add_51_79_groupi_n_3268 ,csa_tree_add_51_79_groupi_n_763);
  and csa_tree_add_51_79_groupi_g40341(csa_tree_add_51_79_groupi_n_5752 ,csa_tree_add_51_79_groupi_n_4985 ,csa_tree_add_51_79_groupi_n_4817);
  or csa_tree_add_51_79_groupi_g40342(csa_tree_add_51_79_groupi_n_5751 ,csa_tree_add_51_79_groupi_n_4898 ,csa_tree_add_51_79_groupi_n_4805);
  or csa_tree_add_51_79_groupi_g40343(csa_tree_add_51_79_groupi_n_5750 ,csa_tree_add_51_79_groupi_n_4401 ,csa_tree_add_51_79_groupi_n_5109);
  or csa_tree_add_51_79_groupi_g40344(csa_tree_add_51_79_groupi_n_5749 ,csa_tree_add_51_79_groupi_n_6 ,csa_tree_add_51_79_groupi_n_2);
  and csa_tree_add_51_79_groupi_g40345(csa_tree_add_51_79_groupi_n_5748 ,csa_tree_add_51_79_groupi_n_4818 ,csa_tree_add_51_79_groupi_n_4819);
  or csa_tree_add_51_79_groupi_g40346(csa_tree_add_51_79_groupi_n_5747 ,csa_tree_add_51_79_groupi_n_4835 ,csa_tree_add_51_79_groupi_n_4798);
  or csa_tree_add_51_79_groupi_g40347(csa_tree_add_51_79_groupi_n_5746 ,csa_tree_add_51_79_groupi_n_4820 ,csa_tree_add_51_79_groupi_n_5338);
  nor csa_tree_add_51_79_groupi_g40348(csa_tree_add_51_79_groupi_n_5745 ,csa_tree_add_51_79_groupi_n_3290 ,csa_tree_add_51_79_groupi_n_5250);
  or csa_tree_add_51_79_groupi_g40349(csa_tree_add_51_79_groupi_n_5744 ,csa_tree_add_51_79_groupi_n_4978 ,csa_tree_add_51_79_groupi_n_5170);
  or csa_tree_add_51_79_groupi_g40350(csa_tree_add_51_79_groupi_n_5743 ,csa_tree_add_51_79_groupi_n_3226 ,csa_tree_add_51_79_groupi_n_4824);
  and csa_tree_add_51_79_groupi_g40351(csa_tree_add_51_79_groupi_n_5742 ,csa_tree_add_51_79_groupi_n_4820 ,csa_tree_add_51_79_groupi_n_5338);
  or csa_tree_add_51_79_groupi_g40352(csa_tree_add_51_79_groupi_n_5741 ,csa_tree_add_51_79_groupi_n_4822 ,csa_tree_add_51_79_groupi_n_4809);
  or csa_tree_add_51_79_groupi_g40353(csa_tree_add_51_79_groupi_n_5740 ,csa_tree_add_51_79_groupi_n_4826 ,csa_tree_add_51_79_groupi_n_4833);
  and csa_tree_add_51_79_groupi_g40354(csa_tree_add_51_79_groupi_n_5739 ,csa_tree_add_51_79_groupi_n_4822 ,csa_tree_add_51_79_groupi_n_4809);
  or csa_tree_add_51_79_groupi_g40355(csa_tree_add_51_79_groupi_n_5738 ,csa_tree_add_51_79_groupi_n_4829 ,csa_tree_add_51_79_groupi_n_4830);
  and csa_tree_add_51_79_groupi_g40356(csa_tree_add_51_79_groupi_n_5737 ,csa_tree_add_51_79_groupi_n_4829 ,csa_tree_add_51_79_groupi_n_4830);
  and csa_tree_add_51_79_groupi_g40357(csa_tree_add_51_79_groupi_n_5736 ,csa_tree_add_51_79_groupi_n_4918 ,csa_tree_add_51_79_groupi_n_5209);
  nor csa_tree_add_51_79_groupi_g40358(csa_tree_add_51_79_groupi_n_5735 ,csa_tree_add_51_79_groupi_n_4834 ,csa_tree_add_51_79_groupi_n_4825);
  and csa_tree_add_51_79_groupi_g40359(csa_tree_add_51_79_groupi_n_5734 ,csa_tree_add_51_79_groupi_n_4831 ,csa_tree_add_51_79_groupi_n_4832);
  or csa_tree_add_51_79_groupi_g40360(csa_tree_add_51_79_groupi_n_5733 ,csa_tree_add_51_79_groupi_n_5197 ,csa_tree_add_51_79_groupi_n_5218);
  or csa_tree_add_51_79_groupi_g40361(csa_tree_add_51_79_groupi_n_5732 ,csa_tree_add_51_79_groupi_n_4917 ,csa_tree_add_51_79_groupi_n_5246);
  or csa_tree_add_51_79_groupi_g40362(csa_tree_add_51_79_groupi_n_5731 ,csa_tree_add_51_79_groupi_n_3234 ,csa_tree_add_51_79_groupi_n_5323);
  and csa_tree_add_51_79_groupi_g40363(csa_tree_add_51_79_groupi_n_5730 ,csa_tree_add_51_79_groupi_n_4921 ,csa_tree_add_51_79_groupi_n_5327);
  or csa_tree_add_51_79_groupi_g40364(csa_tree_add_51_79_groupi_n_5729 ,csa_tree_add_51_79_groupi_n_3196 ,csa_tree_add_51_79_groupi_n_5208);
  or csa_tree_add_51_79_groupi_g40365(csa_tree_add_51_79_groupi_n_5728 ,csa_tree_add_51_79_groupi_n_4285 ,csa_tree_add_51_79_groupi_n_4789);
  or csa_tree_add_51_79_groupi_g40366(csa_tree_add_51_79_groupi_n_5727 ,csa_tree_add_51_79_groupi_n_4296 ,csa_tree_add_51_79_groupi_n_4782);
  or csa_tree_add_51_79_groupi_g40367(csa_tree_add_51_79_groupi_n_5726 ,csa_tree_add_51_79_groupi_n_4837 ,csa_tree_add_51_79_groupi_n_5329);
  and csa_tree_add_51_79_groupi_g40368(csa_tree_add_51_79_groupi_n_5725 ,csa_tree_add_51_79_groupi_n_4978 ,csa_tree_add_51_79_groupi_n_5170);
  and csa_tree_add_51_79_groupi_g40369(csa_tree_add_51_79_groupi_n_5724 ,csa_tree_add_51_79_groupi_n_5003 ,csa_tree_add_51_79_groupi_n_5167);
  or csa_tree_add_51_79_groupi_g40370(csa_tree_add_51_79_groupi_n_5723 ,csa_tree_add_51_79_groupi_n_4916 ,csa_tree_add_51_79_groupi_n_5192);
  or csa_tree_add_51_79_groupi_g40371(csa_tree_add_51_79_groupi_n_5722 ,csa_tree_add_51_79_groupi_n_4902 ,csa_tree_add_51_79_groupi_n_5173);
  or csa_tree_add_51_79_groupi_g40372(csa_tree_add_51_79_groupi_n_5721 ,csa_tree_add_51_79_groupi_n_4029 ,csa_tree_add_51_79_groupi_n_5103);
  and csa_tree_add_51_79_groupi_g40373(csa_tree_add_51_79_groupi_n_5720 ,csa_tree_add_51_79_groupi_n_5252 ,csa_tree_add_51_79_groupi_n_5262);
  or csa_tree_add_51_79_groupi_g40374(csa_tree_add_51_79_groupi_n_5719 ,csa_tree_add_51_79_groupi_n_4576 ,csa_tree_add_51_79_groupi_n_8);
  and csa_tree_add_51_79_groupi_g40375(csa_tree_add_51_79_groupi_n_5718 ,csa_tree_add_51_79_groupi_n_4898 ,csa_tree_add_51_79_groupi_n_4805);
  and csa_tree_add_51_79_groupi_g40376(csa_tree_add_51_79_groupi_n_5717 ,csa_tree_add_51_79_groupi_n_3264 ,csa_tree_add_51_79_groupi_n_4864);
  and csa_tree_add_51_79_groupi_g40377(csa_tree_add_51_79_groupi_n_5716 ,csa_tree_add_51_79_groupi_n_5217 ,csa_tree_add_51_79_groupi_n_4843);
  and csa_tree_add_51_79_groupi_g40378(csa_tree_add_51_79_groupi_n_5715 ,csa_tree_add_51_79_groupi_n_4974 ,csa_tree_add_51_79_groupi_n_4842);
  nor csa_tree_add_51_79_groupi_g40379(csa_tree_add_51_79_groupi_n_5714 ,csa_tree_add_51_79_groupi_n_3264 ,csa_tree_add_51_79_groupi_n_4864);
  or csa_tree_add_51_79_groupi_g40380(csa_tree_add_51_79_groupi_n_5713 ,csa_tree_add_51_79_groupi_n_5334 ,csa_tree_add_51_79_groupi_n_4844);
  nor csa_tree_add_51_79_groupi_g40381(csa_tree_add_51_79_groupi_n_5712 ,csa_tree_add_51_79_groupi_n_3773 ,csa_tree_add_51_79_groupi_n_5274);
  and csa_tree_add_51_79_groupi_g40382(csa_tree_add_51_79_groupi_n_5711 ,csa_tree_add_51_79_groupi_n_4837 ,csa_tree_add_51_79_groupi_n_5329);
  and csa_tree_add_51_79_groupi_g40383(csa_tree_add_51_79_groupi_n_5710 ,csa_tree_add_51_79_groupi_n_3269 ,csa_tree_add_51_79_groupi_n_4860);
  and csa_tree_add_51_79_groupi_g40384(csa_tree_add_51_79_groupi_n_5709 ,csa_tree_add_51_79_groupi_n_5334 ,csa_tree_add_51_79_groupi_n_4844);
  and csa_tree_add_51_79_groupi_g40385(csa_tree_add_51_79_groupi_n_5708 ,csa_tree_add_51_79_groupi_n_4944 ,csa_tree_add_51_79_groupi_n_5420);
  and csa_tree_add_51_79_groupi_g40386(csa_tree_add_51_79_groupi_n_5707 ,csa_tree_add_51_79_groupi_n_4186 ,csa_tree_add_51_79_groupi_n_5499);
  and csa_tree_add_51_79_groupi_g40387(csa_tree_add_51_79_groupi_n_5706 ,csa_tree_add_51_79_groupi_n_4859 ,csa_tree_add_51_79_groupi_n_5419);
  and csa_tree_add_51_79_groupi_g40388(csa_tree_add_51_79_groupi_n_5705 ,csa_tree_add_51_79_groupi_n_4980 ,csa_tree_add_51_79_groupi_n_5156);
  or csa_tree_add_51_79_groupi_g40389(csa_tree_add_51_79_groupi_n_5704 ,csa_tree_add_51_79_groupi_n_4970 ,csa_tree_add_51_79_groupi_n_4808);
  or csa_tree_add_51_79_groupi_g40390(csa_tree_add_51_79_groupi_n_5703 ,csa_tree_add_51_79_groupi_n_3240 ,csa_tree_add_51_79_groupi_n_4796);
  or csa_tree_add_51_79_groupi_g40391(csa_tree_add_51_79_groupi_n_5702 ,csa_tree_add_51_79_groupi_n_4894 ,csa_tree_add_51_79_groupi_n_4846);
  and csa_tree_add_51_79_groupi_g40392(csa_tree_add_51_79_groupi_n_5701 ,csa_tree_add_51_79_groupi_n_4894 ,csa_tree_add_51_79_groupi_n_4846);
  and csa_tree_add_51_79_groupi_g40393(csa_tree_add_51_79_groupi_n_5700 ,csa_tree_add_51_79_groupi_n_3814 ,csa_tree_add_51_79_groupi_n_4845);
  or csa_tree_add_51_79_groupi_g40394(csa_tree_add_51_79_groupi_n_5699 ,csa_tree_add_51_79_groupi_n_4847 ,csa_tree_add_51_79_groupi_n_4849);
  or csa_tree_add_51_79_groupi_g40395(csa_tree_add_51_79_groupi_n_5698 ,csa_tree_add_51_79_groupi_n_4893 ,csa_tree_add_51_79_groupi_n_4848);
  or csa_tree_add_51_79_groupi_g40396(csa_tree_add_51_79_groupi_n_5697 ,csa_tree_add_51_79_groupi_n_5238 ,csa_tree_add_51_79_groupi_n_5232);
  or csa_tree_add_51_79_groupi_g40397(csa_tree_add_51_79_groupi_n_5696 ,csa_tree_add_51_79_groupi_n_5293 ,csa_tree_add_51_79_groupi_n_4851);
  and csa_tree_add_51_79_groupi_g40398(csa_tree_add_51_79_groupi_n_5695 ,csa_tree_add_51_79_groupi_n_5293 ,csa_tree_add_51_79_groupi_n_4851);
  or csa_tree_add_51_79_groupi_g40399(csa_tree_add_51_79_groupi_n_5694 ,csa_tree_add_51_79_groupi_n_4890 ,csa_tree_add_51_79_groupi_n_4854);
  and csa_tree_add_51_79_groupi_g40400(csa_tree_add_51_79_groupi_n_5693 ,csa_tree_add_51_79_groupi_n_4847 ,csa_tree_add_51_79_groupi_n_4849);
  or csa_tree_add_51_79_groupi_g40401(csa_tree_add_51_79_groupi_n_5692 ,csa_tree_add_51_79_groupi_n_4856 ,csa_tree_add_51_79_groupi_n_4857);
  and csa_tree_add_51_79_groupi_g40402(csa_tree_add_51_79_groupi_n_5691 ,csa_tree_add_51_79_groupi_n_4890 ,csa_tree_add_51_79_groupi_n_4854);
  and csa_tree_add_51_79_groupi_g40403(csa_tree_add_51_79_groupi_n_5690 ,csa_tree_add_51_79_groupi_n_4973 ,csa_tree_add_51_79_groupi_n_5164);
  or csa_tree_add_51_79_groupi_g40404(csa_tree_add_51_79_groupi_n_5689 ,csa_tree_add_51_79_groupi_n_3291 ,csa_tree_add_51_79_groupi_n_4862);
  and csa_tree_add_51_79_groupi_g40405(csa_tree_add_51_79_groupi_n_5688 ,csa_tree_add_51_79_groupi_n_4814 ,csa_tree_add_51_79_groupi_n_5413);
  or csa_tree_add_51_79_groupi_g40406(csa_tree_add_51_79_groupi_n_5687 ,csa_tree_add_51_79_groupi_n_4814 ,csa_tree_add_51_79_groupi_n_5413);
  nor csa_tree_add_51_79_groupi_g40407(csa_tree_add_51_79_groupi_n_5686 ,csa_tree_add_51_79_groupi_n_4858 ,csa_tree_add_51_79_groupi_n_4855);
  or csa_tree_add_51_79_groupi_g40408(csa_tree_add_51_79_groupi_n_5685 ,csa_tree_add_51_79_groupi_n_3816 ,csa_tree_add_51_79_groupi_n_5211);
  or csa_tree_add_51_79_groupi_g40409(csa_tree_add_51_79_groupi_n_5684 ,csa_tree_add_51_79_groupi_n_3798 ,csa_tree_add_51_79_groupi_n_4866);
  and csa_tree_add_51_79_groupi_g40410(csa_tree_add_51_79_groupi_n_5683 ,csa_tree_add_51_79_groupi_n_5411 ,csa_tree_add_51_79_groupi_n_4836);
  or csa_tree_add_51_79_groupi_g40411(csa_tree_add_51_79_groupi_n_5682 ,csa_tree_add_51_79_groupi_n_4867 ,csa_tree_add_51_79_groupi_n_4868);
  nor csa_tree_add_51_79_groupi_g40412(csa_tree_add_51_79_groupi_n_5681 ,csa_tree_add_51_79_groupi_n_3799 ,csa_tree_add_51_79_groupi_n_4865);
  or csa_tree_add_51_79_groupi_g40413(csa_tree_add_51_79_groupi_n_5680 ,csa_tree_add_51_79_groupi_n_4870 ,csa_tree_add_51_79_groupi_n_4873);
  and csa_tree_add_51_79_groupi_g40414(csa_tree_add_51_79_groupi_n_5679 ,csa_tree_add_51_79_groupi_n_4867 ,csa_tree_add_51_79_groupi_n_4868);
  or csa_tree_add_51_79_groupi_g40415(csa_tree_add_51_79_groupi_n_5678 ,csa_tree_add_51_79_groupi_n_4871 ,csa_tree_add_51_79_groupi_n_4872);
  or csa_tree_add_51_79_groupi_g40416(csa_tree_add_51_79_groupi_n_5677 ,csa_tree_add_51_79_groupi_n_4289 ,csa_tree_add_51_79_groupi_n_4792);
  nor csa_tree_add_51_79_groupi_g40417(csa_tree_add_51_79_groupi_n_5676 ,csa_tree_add_51_79_groupi_n_1210 ,csa_tree_add_51_79_groupi_n_4811);
  and csa_tree_add_51_79_groupi_g40418(csa_tree_add_51_79_groupi_n_5675 ,csa_tree_add_51_79_groupi_n_4871 ,csa_tree_add_51_79_groupi_n_4872);
  or csa_tree_add_51_79_groupi_g40419(csa_tree_add_51_79_groupi_n_5674 ,csa_tree_add_51_79_groupi_n_4875 ,csa_tree_add_51_79_groupi_n_4876);
  or csa_tree_add_51_79_groupi_g40420(csa_tree_add_51_79_groupi_n_5673 ,csa_tree_add_51_79_groupi_n_4288 ,csa_tree_add_51_79_groupi_n_4781);
  and csa_tree_add_51_79_groupi_g40421(csa_tree_add_51_79_groupi_n_5672 ,csa_tree_add_51_79_groupi_n_4875 ,csa_tree_add_51_79_groupi_n_4876);
  nor csa_tree_add_51_79_groupi_g40422(csa_tree_add_51_79_groupi_n_5671 ,csa_tree_add_51_79_groupi_n_4874 ,csa_tree_add_51_79_groupi_n_4869);
  or csa_tree_add_51_79_groupi_g40423(csa_tree_add_51_79_groupi_n_5670 ,csa_tree_add_51_79_groupi_n_4987 ,csa_tree_add_51_79_groupi_n_4877);
  or csa_tree_add_51_79_groupi_g40424(csa_tree_add_51_79_groupi_n_5669 ,csa_tree_add_51_79_groupi_n_4878 ,csa_tree_add_51_79_groupi_n_4879);
  and csa_tree_add_51_79_groupi_g40425(csa_tree_add_51_79_groupi_n_5668 ,csa_tree_add_51_79_groupi_n_3246 ,csa_tree_add_51_79_groupi_n_4887);
  and csa_tree_add_51_79_groupi_g40426(csa_tree_add_51_79_groupi_n_5667 ,csa_tree_add_51_79_groupi_n_4987 ,csa_tree_add_51_79_groupi_n_4877);
  or csa_tree_add_51_79_groupi_g40427(csa_tree_add_51_79_groupi_n_5666 ,csa_tree_add_51_79_groupi_n_4880 ,csa_tree_add_51_79_groupi_n_4883);
  and csa_tree_add_51_79_groupi_g40428(csa_tree_add_51_79_groupi_n_5665 ,csa_tree_add_51_79_groupi_n_4880 ,csa_tree_add_51_79_groupi_n_4883);
  or csa_tree_add_51_79_groupi_g40429(csa_tree_add_51_79_groupi_n_5664 ,csa_tree_add_51_79_groupi_n_4886 ,csa_tree_add_51_79_groupi_n_4888);
  and csa_tree_add_51_79_groupi_g40430(csa_tree_add_51_79_groupi_n_5663 ,csa_tree_add_51_79_groupi_n_4878 ,csa_tree_add_51_79_groupi_n_4879);
  and csa_tree_add_51_79_groupi_g40431(csa_tree_add_51_79_groupi_n_5662 ,csa_tree_add_51_79_groupi_n_4886 ,csa_tree_add_51_79_groupi_n_4888);
  or csa_tree_add_51_79_groupi_g40432(csa_tree_add_51_79_groupi_n_5661 ,csa_tree_add_51_79_groupi_n_4297 ,csa_tree_add_51_79_groupi_n_4786);
  or csa_tree_add_51_79_groupi_g40433(csa_tree_add_51_79_groupi_n_5660 ,csa_tree_add_51_79_groupi_n_4298 ,csa_tree_add_51_79_groupi_n_4769);
  or csa_tree_add_51_79_groupi_g40434(csa_tree_add_51_79_groupi_n_5659 ,csa_tree_add_51_79_groupi_n_4299 ,csa_tree_add_51_79_groupi_n_4767);
  nor csa_tree_add_51_79_groupi_g40435(csa_tree_add_51_79_groupi_n_5658 ,csa_tree_add_51_79_groupi_n_3292 ,csa_tree_add_51_79_groupi_n_4863);
  nor csa_tree_add_51_79_groupi_g40436(csa_tree_add_51_79_groupi_n_5657 ,csa_tree_add_51_79_groupi_n_3246 ,csa_tree_add_51_79_groupi_n_4887);
  and csa_tree_add_51_79_groupi_g40437(csa_tree_add_51_79_groupi_n_5656 ,csa_tree_add_51_79_groupi_n_3204 ,csa_tree_add_51_79_groupi_n_4904);
  or csa_tree_add_51_79_groupi_g40438(csa_tree_add_51_79_groupi_n_5655 ,csa_tree_add_51_79_groupi_n_3930 ,csa_tree_add_51_79_groupi_n_5059);
  or csa_tree_add_51_79_groupi_g40439(csa_tree_add_51_79_groupi_n_5654 ,csa_tree_add_51_79_groupi_n_765 ,csa_tree_add_51_79_groupi_n_4908);
  or csa_tree_add_51_79_groupi_g40440(csa_tree_add_51_79_groupi_n_5653 ,csa_tree_add_51_79_groupi_n_4909 ,csa_tree_add_51_79_groupi_n_4910);
  and csa_tree_add_51_79_groupi_g40441(csa_tree_add_51_79_groupi_n_5652 ,csa_tree_add_51_79_groupi_n_765 ,csa_tree_add_51_79_groupi_n_4908);
  or csa_tree_add_51_79_groupi_g40442(csa_tree_add_51_79_groupi_n_5651 ,csa_tree_add_51_79_groupi_n_4300 ,csa_tree_add_51_79_groupi_n_4761);
  and csa_tree_add_51_79_groupi_g40443(csa_tree_add_51_79_groupi_n_5650 ,csa_tree_add_51_79_groupi_n_4909 ,csa_tree_add_51_79_groupi_n_4910);
  or csa_tree_add_51_79_groupi_g40444(csa_tree_add_51_79_groupi_n_5649 ,csa_tree_add_51_79_groupi_n_4912 ,csa_tree_add_51_79_groupi_n_4914);
  and csa_tree_add_51_79_groupi_g40445(csa_tree_add_51_79_groupi_n_5648 ,csa_tree_add_51_79_groupi_n_4912 ,csa_tree_add_51_79_groupi_n_4914);
  or csa_tree_add_51_79_groupi_g40446(csa_tree_add_51_79_groupi_n_5647 ,csa_tree_add_51_79_groupi_n_4885 ,csa_tree_add_51_79_groupi_n_4920);
  or csa_tree_add_51_79_groupi_g40447(csa_tree_add_51_79_groupi_n_5646 ,csa_tree_add_51_79_groupi_n_3259 ,csa_tree_add_51_79_groupi_n_4922);
  and csa_tree_add_51_79_groupi_g40448(csa_tree_add_51_79_groupi_n_5645 ,csa_tree_add_51_79_groupi_n_4885 ,csa_tree_add_51_79_groupi_n_4920);
  or csa_tree_add_51_79_groupi_g40449(csa_tree_add_51_79_groupi_n_5644 ,csa_tree_add_51_79_groupi_n_4884 ,csa_tree_add_51_79_groupi_n_4926);
  and csa_tree_add_51_79_groupi_g40450(csa_tree_add_51_79_groupi_n_5643 ,csa_tree_add_51_79_groupi_n_4884 ,csa_tree_add_51_79_groupi_n_4926);
  or csa_tree_add_51_79_groupi_g40451(csa_tree_add_51_79_groupi_n_5642 ,csa_tree_add_51_79_groupi_n_4928 ,csa_tree_add_51_79_groupi_n_4930);
  and csa_tree_add_51_79_groupi_g40452(csa_tree_add_51_79_groupi_n_5641 ,csa_tree_add_51_79_groupi_n_3281 ,csa_tree_add_51_79_groupi_n_4941);
  nor csa_tree_add_51_79_groupi_g40453(csa_tree_add_51_79_groupi_n_5640 ,csa_tree_add_51_79_groupi_n_3204 ,csa_tree_add_51_79_groupi_n_4904);
  and csa_tree_add_51_79_groupi_g40454(csa_tree_add_51_79_groupi_n_5639 ,csa_tree_add_51_79_groupi_n_4928 ,csa_tree_add_51_79_groupi_n_4930);
  nor csa_tree_add_51_79_groupi_g40455(csa_tree_add_51_79_groupi_n_5638 ,csa_tree_add_51_79_groupi_n_3260 ,csa_tree_add_51_79_groupi_n_4923);
  or csa_tree_add_51_79_groupi_g40456(csa_tree_add_51_79_groupi_n_5637 ,csa_tree_add_51_79_groupi_n_4889 ,csa_tree_add_51_79_groupi_n_4850);
  or csa_tree_add_51_79_groupi_g40457(csa_tree_add_51_79_groupi_n_5636 ,csa_tree_add_51_79_groupi_n_4936 ,csa_tree_add_51_79_groupi_n_4939);
  nor csa_tree_add_51_79_groupi_g40458(csa_tree_add_51_79_groupi_n_5635 ,csa_tree_add_51_79_groupi_n_3269 ,csa_tree_add_51_79_groupi_n_4860);
  and csa_tree_add_51_79_groupi_g40459(csa_tree_add_51_79_groupi_n_5634 ,csa_tree_add_51_79_groupi_n_3280 ,csa_tree_add_51_79_groupi_n_4942);
  and csa_tree_add_51_79_groupi_g40460(csa_tree_add_51_79_groupi_n_5633 ,csa_tree_add_51_79_groupi_n_4889 ,csa_tree_add_51_79_groupi_n_4850);
  and csa_tree_add_51_79_groupi_g40461(csa_tree_add_51_79_groupi_n_5632 ,csa_tree_add_51_79_groupi_n_4902 ,csa_tree_add_51_79_groupi_n_5173);
  and csa_tree_add_51_79_groupi_g40462(csa_tree_add_51_79_groupi_n_5631 ,csa_tree_add_51_79_groupi_n_4936 ,csa_tree_add_51_79_groupi_n_4939);
  or csa_tree_add_51_79_groupi_g40463(csa_tree_add_51_79_groupi_n_5630 ,csa_tree_add_51_79_groupi_n_5285 ,csa_tree_add_51_79_groupi_n_5284);
  or csa_tree_add_51_79_groupi_g40464(csa_tree_add_51_79_groupi_n_5629 ,csa_tree_add_51_79_groupi_n_4943 ,csa_tree_add_51_79_groupi_n_4949);
  and csa_tree_add_51_79_groupi_g40465(csa_tree_add_51_79_groupi_n_5628 ,csa_tree_add_51_79_groupi_n_4943 ,csa_tree_add_51_79_groupi_n_4949);
  or csa_tree_add_51_79_groupi_g40466(csa_tree_add_51_79_groupi_n_5627 ,csa_tree_add_51_79_groupi_n_5010 ,csa_tree_add_51_79_groupi_n_4950);
  and csa_tree_add_51_79_groupi_g40467(csa_tree_add_51_79_groupi_n_5626 ,csa_tree_add_51_79_groupi_n_5010 ,csa_tree_add_51_79_groupi_n_4950);
  or csa_tree_add_51_79_groupi_g40468(csa_tree_add_51_79_groupi_n_5625 ,csa_tree_add_51_79_groupi_n_4951 ,csa_tree_add_51_79_groupi_n_4954);
  and csa_tree_add_51_79_groupi_g40469(csa_tree_add_51_79_groupi_n_5624 ,csa_tree_add_51_79_groupi_n_4951 ,csa_tree_add_51_79_groupi_n_4954);
  nor csa_tree_add_51_79_groupi_g40470(csa_tree_add_51_79_groupi_n_5623 ,csa_tree_add_51_79_groupi_n_3280 ,csa_tree_add_51_79_groupi_n_4942);
  nor csa_tree_add_51_79_groupi_g40471(csa_tree_add_51_79_groupi_n_5622 ,csa_tree_add_51_79_groupi_n_4957 ,csa_tree_add_51_79_groupi_n_4962);
  or csa_tree_add_51_79_groupi_g40472(csa_tree_add_51_79_groupi_n_5621 ,csa_tree_add_51_79_groupi_n_3272 ,csa_tree_add_51_79_groupi_n_5291);
  or csa_tree_add_51_79_groupi_g40473(csa_tree_add_51_79_groupi_n_5620 ,csa_tree_add_51_79_groupi_n_4882 ,csa_tree_add_51_79_groupi_n_4966);
  nor csa_tree_add_51_79_groupi_g40474(csa_tree_add_51_79_groupi_n_5619 ,csa_tree_add_51_79_groupi_n_3281 ,csa_tree_add_51_79_groupi_n_4941);
  or csa_tree_add_51_79_groupi_g40475(csa_tree_add_51_79_groupi_n_5618 ,csa_tree_add_51_79_groupi_n_4292 ,csa_tree_add_51_79_groupi_n_4757);
  and csa_tree_add_51_79_groupi_g40476(csa_tree_add_51_79_groupi_n_5617 ,csa_tree_add_51_79_groupi_n_4882 ,csa_tree_add_51_79_groupi_n_4966);
  or csa_tree_add_51_79_groupi_g40477(csa_tree_add_51_79_groupi_n_5616 ,csa_tree_add_51_79_groupi_n_4956 ,csa_tree_add_51_79_groupi_n_4961);
  and csa_tree_add_51_79_groupi_g40478(csa_tree_add_51_79_groupi_n_5615 ,csa_tree_add_51_79_groupi_n_5356 ,csa_tree_add_51_79_groupi_n_4852);
  or csa_tree_add_51_79_groupi_g40479(csa_tree_add_51_79_groupi_n_5614 ,csa_tree_add_51_79_groupi_n_3304 ,csa_tree_add_51_79_groupi_n_4958);
  or csa_tree_add_51_79_groupi_g40480(csa_tree_add_51_79_groupi_n_5613 ,csa_tree_add_51_79_groupi_n_4976 ,csa_tree_add_51_79_groupi_n_4977);
  and csa_tree_add_51_79_groupi_g40481(csa_tree_add_51_79_groupi_n_5612 ,csa_tree_add_51_79_groupi_n_3233 ,csa_tree_add_51_79_groupi_n_5362);
  or csa_tree_add_51_79_groupi_g40482(csa_tree_add_51_79_groupi_n_5611 ,csa_tree_add_51_79_groupi_n_4831 ,csa_tree_add_51_79_groupi_n_4832);
  and csa_tree_add_51_79_groupi_g40483(csa_tree_add_51_79_groupi_n_5610 ,csa_tree_add_51_79_groupi_n_4925 ,csa_tree_add_51_79_groupi_n_4924);
  or csa_tree_add_51_79_groupi_g40484(csa_tree_add_51_79_groupi_n_5609 ,csa_tree_add_51_79_groupi_n_4934 ,csa_tree_add_51_79_groupi_n_4933);
  and csa_tree_add_51_79_groupi_g40485(csa_tree_add_51_79_groupi_n_5608 ,csa_tree_add_51_79_groupi_n_4911 ,csa_tree_add_51_79_groupi_n_5009);
  or csa_tree_add_51_79_groupi_g40486(csa_tree_add_51_79_groupi_n_5607 ,csa_tree_add_51_79_groupi_n_4925 ,csa_tree_add_51_79_groupi_n_4924);
  or csa_tree_add_51_79_groupi_g40487(csa_tree_add_51_79_groupi_n_5606 ,csa_tree_add_51_79_groupi_n_4929 ,csa_tree_add_51_79_groupi_n_4927);
  or csa_tree_add_51_79_groupi_g40488(csa_tree_add_51_79_groupi_n_5605 ,csa_tree_add_51_79_groupi_n_4915 ,csa_tree_add_51_79_groupi_n_5005);
  and csa_tree_add_51_79_groupi_g40489(csa_tree_add_51_79_groupi_n_5604 ,csa_tree_add_51_79_groupi_n_4915 ,csa_tree_add_51_79_groupi_n_5005);
  or csa_tree_add_51_79_groupi_g40490(csa_tree_add_51_79_groupi_n_5603 ,csa_tree_add_51_79_groupi_n_4899 ,csa_tree_add_51_79_groupi_n_4913);
  and csa_tree_add_51_79_groupi_g40491(csa_tree_add_51_79_groupi_n_5602 ,csa_tree_add_51_79_groupi_n_4899 ,csa_tree_add_51_79_groupi_n_4913);
  or csa_tree_add_51_79_groupi_g40492(csa_tree_add_51_79_groupi_n_5601 ,csa_tree_add_51_79_groupi_n_4911 ,csa_tree_add_51_79_groupi_n_5009);
  and csa_tree_add_51_79_groupi_g40493(csa_tree_add_51_79_groupi_n_5600 ,csa_tree_add_51_79_groupi_n_4934 ,csa_tree_add_51_79_groupi_n_4933);
  or csa_tree_add_51_79_groupi_g40494(csa_tree_add_51_79_groupi_n_5599 ,csa_tree_add_51_79_groupi_n_4982 ,csa_tree_add_51_79_groupi_n_4907);
  and csa_tree_add_51_79_groupi_g40495(csa_tree_add_51_79_groupi_n_5598 ,csa_tree_add_51_79_groupi_n_4982 ,csa_tree_add_51_79_groupi_n_4907);
  and csa_tree_add_51_79_groupi_g40496(csa_tree_add_51_79_groupi_n_5597 ,csa_tree_add_51_79_groupi_n_4929 ,csa_tree_add_51_79_groupi_n_4927);
  or csa_tree_add_51_79_groupi_g40497(csa_tree_add_51_79_groupi_n_5596 ,csa_tree_add_51_79_groupi_n_4286 ,csa_tree_add_51_79_groupi_n_4755);
  or csa_tree_add_51_79_groupi_g40498(csa_tree_add_51_79_groupi_n_5595 ,csa_tree_add_51_79_groupi_n_4287 ,csa_tree_add_51_79_groupi_n_4762);
  xnor csa_tree_add_51_79_groupi_g40499(csa_tree_add_51_79_groupi_n_5594 ,csa_tree_add_51_79_groupi_n_4251 ,csa_tree_add_51_79_groupi_n_4249);
  xnor csa_tree_add_51_79_groupi_g40500(csa_tree_add_51_79_groupi_n_5593 ,csa_tree_add_51_79_groupi_n_4225 ,csa_tree_add_51_79_groupi_n_4226);
  xnor csa_tree_add_51_79_groupi_g40501(csa_tree_add_51_79_groupi_n_5592 ,csa_tree_add_51_79_groupi_n_4236 ,csa_tree_add_51_79_groupi_n_4267);
  xnor csa_tree_add_51_79_groupi_g40502(csa_tree_add_51_79_groupi_n_5591 ,csa_tree_add_51_79_groupi_n_4234 ,csa_tree_add_51_79_groupi_n_4235);
  xnor csa_tree_add_51_79_groupi_g40503(csa_tree_add_51_79_groupi_n_5590 ,csa_tree_add_51_79_groupi_n_4243 ,csa_tree_add_51_79_groupi_n_4230);
  xnor csa_tree_add_51_79_groupi_g40504(csa_tree_add_51_79_groupi_n_5589 ,csa_tree_add_51_79_groupi_n_4260 ,csa_tree_add_51_79_groupi_n_4231);
  xnor csa_tree_add_51_79_groupi_g40505(csa_tree_add_51_79_groupi_n_5588 ,csa_tree_add_51_79_groupi_n_4238 ,csa_tree_add_51_79_groupi_n_4233);
  xnor csa_tree_add_51_79_groupi_g40506(csa_tree_add_51_79_groupi_n_5587 ,csa_tree_add_51_79_groupi_n_4245 ,csa_tree_add_51_79_groupi_n_4253);
  xnor csa_tree_add_51_79_groupi_g40507(csa_tree_add_51_79_groupi_n_5586 ,csa_tree_add_51_79_groupi_n_4266 ,csa_tree_add_51_79_groupi_n_4264);
  xnor csa_tree_add_51_79_groupi_g40508(csa_tree_add_51_79_groupi_n_5585 ,csa_tree_add_51_79_groupi_n_4255 ,csa_tree_add_51_79_groupi_n_4283);
  xnor csa_tree_add_51_79_groupi_g40509(csa_tree_add_51_79_groupi_n_5584 ,csa_tree_add_51_79_groupi_n_4242 ,csa_tree_add_51_79_groupi_n_4262);
  xnor csa_tree_add_51_79_groupi_g40510(csa_tree_add_51_79_groupi_n_5583 ,csa_tree_add_51_79_groupi_n_4228 ,csa_tree_add_51_79_groupi_n_4275);
  xnor csa_tree_add_51_79_groupi_g40511(csa_tree_add_51_79_groupi_n_5582 ,csa_tree_add_51_79_groupi_n_4269 ,csa_tree_add_51_79_groupi_n_4271);
  xnor csa_tree_add_51_79_groupi_g40512(csa_tree_add_51_79_groupi_n_5581 ,csa_tree_add_51_79_groupi_n_4281 ,csa_tree_add_51_79_groupi_n_4279);
  xnor csa_tree_add_51_79_groupi_g40513(csa_tree_add_51_79_groupi_n_5580 ,csa_tree_add_51_79_groupi_n_4259 ,csa_tree_add_51_79_groupi_n_4240);
  xnor csa_tree_add_51_79_groupi_g40514(csa_tree_add_51_79_groupi_n_5579 ,csa_tree_add_51_79_groupi_n_4247 ,csa_tree_add_51_79_groupi_n_4257);
  xnor csa_tree_add_51_79_groupi_g40515(csa_tree_add_51_79_groupi_n_5578 ,csa_tree_add_51_79_groupi_n_4277 ,csa_tree_add_51_79_groupi_n_4273);
  and csa_tree_add_51_79_groupi_g40516(csa_tree_add_51_79_groupi_n_5868 ,csa_tree_add_51_79_groupi_n_4192 ,csa_tree_add_51_79_groupi_n_5129);
  and csa_tree_add_51_79_groupi_g40517(csa_tree_add_51_79_groupi_n_5867 ,csa_tree_add_51_79_groupi_n_4633 ,csa_tree_add_51_79_groupi_n_4791);
  and csa_tree_add_51_79_groupi_g40518(csa_tree_add_51_79_groupi_n_5866 ,csa_tree_add_51_79_groupi_n_4194 ,csa_tree_add_51_79_groupi_n_5147);
  or csa_tree_add_51_79_groupi_g40519(csa_tree_add_51_79_groupi_n_5865 ,csa_tree_add_51_79_groupi_n_5076 ,csa_tree_add_51_79_groupi_n_5559);
  xnor csa_tree_add_51_79_groupi_g40520(csa_tree_add_51_79_groupi_n_5864 ,csa_tree_add_51_79_groupi_n_2571 ,csa_tree_add_51_79_groupi_n_3880);
  and csa_tree_add_51_79_groupi_g40521(csa_tree_add_51_79_groupi_n_5863 ,csa_tree_add_51_79_groupi_n_4617 ,csa_tree_add_51_79_groupi_n_4752);
  and csa_tree_add_51_79_groupi_g40522(csa_tree_add_51_79_groupi_n_5861 ,csa_tree_add_51_79_groupi_n_4303 ,csa_tree_add_51_79_groupi_n_5126);
  and csa_tree_add_51_79_groupi_g40523(csa_tree_add_51_79_groupi_n_5860 ,csa_tree_add_51_79_groupi_n_4320 ,csa_tree_add_51_79_groupi_n_5134);
  and csa_tree_add_51_79_groupi_g40524(csa_tree_add_51_79_groupi_n_5859 ,csa_tree_add_51_79_groupi_n_4713 ,csa_tree_add_51_79_groupi_n_5141);
  xnor csa_tree_add_51_79_groupi_g40525(csa_tree_add_51_79_groupi_n_5858 ,csa_tree_add_51_79_groupi_n_2567 ,csa_tree_add_51_79_groupi_n_3876);
  xnor csa_tree_add_51_79_groupi_g40526(csa_tree_add_51_79_groupi_n_5856 ,csa_tree_add_51_79_groupi_n_2548 ,csa_tree_add_51_79_groupi_n_3874);
  xnor csa_tree_add_51_79_groupi_g40527(csa_tree_add_51_79_groupi_n_5854 ,csa_tree_add_51_79_groupi_n_2544 ,csa_tree_add_51_79_groupi_n_3875);
  or csa_tree_add_51_79_groupi_g40528(csa_tree_add_51_79_groupi_n_5853 ,csa_tree_add_51_79_groupi_n_3973 ,csa_tree_add_51_79_groupi_n_4758);
  or csa_tree_add_51_79_groupi_g40529(csa_tree_add_51_79_groupi_n_5851 ,csa_tree_add_51_79_groupi_n_3963 ,csa_tree_add_51_79_groupi_n_4751);
  and csa_tree_add_51_79_groupi_g40530(csa_tree_add_51_79_groupi_n_5850 ,csa_tree_add_51_79_groupi_n_3949 ,csa_tree_add_51_79_groupi_n_4754);
  and csa_tree_add_51_79_groupi_g40531(csa_tree_add_51_79_groupi_n_5849 ,csa_tree_add_51_79_groupi_n_3947 ,csa_tree_add_51_79_groupi_n_4753);
  xnor csa_tree_add_51_79_groupi_g40532(csa_tree_add_51_79_groupi_n_5848 ,csa_tree_add_51_79_groupi_n_2543 ,csa_tree_add_51_79_groupi_n_3877);
  xnor csa_tree_add_51_79_groupi_g40533(csa_tree_add_51_79_groupi_n_5846 ,csa_tree_add_51_79_groupi_n_2561 ,csa_tree_add_51_79_groupi_n_3879);
  xnor csa_tree_add_51_79_groupi_g40534(csa_tree_add_51_79_groupi_n_5845 ,csa_tree_add_51_79_groupi_n_2562 ,csa_tree_add_51_79_groupi_n_3878);
  xnor csa_tree_add_51_79_groupi_g40535(csa_tree_add_51_79_groupi_n_5844 ,csa_tree_add_51_79_groupi_n_4229 ,csa_tree_add_51_79_groupi_n_3873);
  and csa_tree_add_51_79_groupi_g40536(csa_tree_add_51_79_groupi_n_5842 ,csa_tree_add_51_79_groupi_n_4302 ,csa_tree_add_51_79_groupi_n_5148);
  or csa_tree_add_51_79_groupi_g40537(csa_tree_add_51_79_groupi_n_5841 ,csa_tree_add_51_79_groupi_n_3935 ,csa_tree_add_51_79_groupi_n_4750);
  not csa_tree_add_51_79_groupi_g40538(csa_tree_add_51_79_groupi_n_5559 ,csa_tree_add_51_79_groupi_n_5558);
  not csa_tree_add_51_79_groupi_g40539(csa_tree_add_51_79_groupi_n_5518 ,csa_tree_add_51_79_groupi_n_5517);
  not csa_tree_add_51_79_groupi_g40540(csa_tree_add_51_79_groupi_n_5454 ,csa_tree_add_51_79_groupi_n_5453);
  not csa_tree_add_51_79_groupi_g40541(csa_tree_add_51_79_groupi_n_5444 ,csa_tree_add_51_79_groupi_n_5443);
  not csa_tree_add_51_79_groupi_g40542(csa_tree_add_51_79_groupi_n_5431 ,csa_tree_add_51_79_groupi_n_5432);
  not csa_tree_add_51_79_groupi_g40543(csa_tree_add_51_79_groupi_n_5425 ,csa_tree_add_51_79_groupi_n_5426);
  not csa_tree_add_51_79_groupi_g40544(csa_tree_add_51_79_groupi_n_5422 ,csa_tree_add_51_79_groupi_n_5423);
  not csa_tree_add_51_79_groupi_g40545(csa_tree_add_51_79_groupi_n_5418 ,csa_tree_add_51_79_groupi_n_5417);
  not csa_tree_add_51_79_groupi_g40546(csa_tree_add_51_79_groupi_n_5415 ,csa_tree_add_51_79_groupi_n_5416);
  not csa_tree_add_51_79_groupi_g40547(csa_tree_add_51_79_groupi_n_5409 ,csa_tree_add_51_79_groupi_n_5410);
  not csa_tree_add_51_79_groupi_g40548(csa_tree_add_51_79_groupi_n_5402 ,csa_tree_add_51_79_groupi_n_5403);
  not csa_tree_add_51_79_groupi_g40549(csa_tree_add_51_79_groupi_n_5400 ,csa_tree_add_51_79_groupi_n_5401);
  not csa_tree_add_51_79_groupi_g40550(csa_tree_add_51_79_groupi_n_5398 ,csa_tree_add_51_79_groupi_n_5399);
  not csa_tree_add_51_79_groupi_g40551(csa_tree_add_51_79_groupi_n_5395 ,csa_tree_add_51_79_groupi_n_5396);
  not csa_tree_add_51_79_groupi_g40552(csa_tree_add_51_79_groupi_n_5389 ,csa_tree_add_51_79_groupi_n_5390);
  not csa_tree_add_51_79_groupi_g40553(csa_tree_add_51_79_groupi_n_5387 ,csa_tree_add_51_79_groupi_n_5388);
  not csa_tree_add_51_79_groupi_g40554(csa_tree_add_51_79_groupi_n_5380 ,csa_tree_add_51_79_groupi_n_5381);
  not csa_tree_add_51_79_groupi_g40555(csa_tree_add_51_79_groupi_n_5374 ,csa_tree_add_51_79_groupi_n_5375);
  not csa_tree_add_51_79_groupi_g40556(csa_tree_add_51_79_groupi_n_5371 ,csa_tree_add_51_79_groupi_n_5372);
  not csa_tree_add_51_79_groupi_g40557(csa_tree_add_51_79_groupi_n_5369 ,csa_tree_add_51_79_groupi_n_5370);
  not csa_tree_add_51_79_groupi_g40558(csa_tree_add_51_79_groupi_n_5366 ,csa_tree_add_51_79_groupi_n_5367);
  not csa_tree_add_51_79_groupi_g40559(csa_tree_add_51_79_groupi_n_5363 ,csa_tree_add_51_79_groupi_n_5364);
  not csa_tree_add_51_79_groupi_g40560(csa_tree_add_51_79_groupi_n_5359 ,csa_tree_add_51_79_groupi_n_5360);
  not csa_tree_add_51_79_groupi_g40561(csa_tree_add_51_79_groupi_n_5354 ,csa_tree_add_51_79_groupi_n_5355);
  not csa_tree_add_51_79_groupi_g40562(csa_tree_add_51_79_groupi_n_5351 ,csa_tree_add_51_79_groupi_n_5352);
  not csa_tree_add_51_79_groupi_g40563(csa_tree_add_51_79_groupi_n_5346 ,csa_tree_add_51_79_groupi_n_5347);
  not csa_tree_add_51_79_groupi_g40564(csa_tree_add_51_79_groupi_n_5342 ,csa_tree_add_51_79_groupi_n_5343);
  not csa_tree_add_51_79_groupi_g40565(csa_tree_add_51_79_groupi_n_5336 ,csa_tree_add_51_79_groupi_n_5337);
  not csa_tree_add_51_79_groupi_g40566(csa_tree_add_51_79_groupi_n_5331 ,csa_tree_add_51_79_groupi_n_5332);
  not csa_tree_add_51_79_groupi_g40567(csa_tree_add_51_79_groupi_n_5327 ,csa_tree_add_51_79_groupi_n_5326);
  not csa_tree_add_51_79_groupi_g40568(csa_tree_add_51_79_groupi_n_5322 ,csa_tree_add_51_79_groupi_n_5323);
  not csa_tree_add_51_79_groupi_g40569(csa_tree_add_51_79_groupi_n_5316 ,csa_tree_add_51_79_groupi_n_5317);
  not csa_tree_add_51_79_groupi_g40570(csa_tree_add_51_79_groupi_n_5313 ,csa_tree_add_51_79_groupi_n_5314);
  not csa_tree_add_51_79_groupi_g40571(csa_tree_add_51_79_groupi_n_5308 ,csa_tree_add_51_79_groupi_n_5309);
  not csa_tree_add_51_79_groupi_g40572(csa_tree_add_51_79_groupi_n_5305 ,csa_tree_add_51_79_groupi_n_5306);
  not csa_tree_add_51_79_groupi_g40573(csa_tree_add_51_79_groupi_n_5302 ,csa_tree_add_51_79_groupi_n_5303);
  not csa_tree_add_51_79_groupi_g40574(csa_tree_add_51_79_groupi_n_5299 ,csa_tree_add_51_79_groupi_n_5300);
  not csa_tree_add_51_79_groupi_g40575(csa_tree_add_51_79_groupi_n_5296 ,csa_tree_add_51_79_groupi_n_5297);
  not csa_tree_add_51_79_groupi_g40576(csa_tree_add_51_79_groupi_n_5291 ,csa_tree_add_51_79_groupi_n_5292);
  not csa_tree_add_51_79_groupi_g40577(csa_tree_add_51_79_groupi_n_5288 ,csa_tree_add_51_79_groupi_n_5289);
  not csa_tree_add_51_79_groupi_g40578(csa_tree_add_51_79_groupi_n_5286 ,csa_tree_add_51_79_groupi_n_5287);
  not csa_tree_add_51_79_groupi_g40579(csa_tree_add_51_79_groupi_n_5280 ,csa_tree_add_51_79_groupi_n_5281);
  not csa_tree_add_51_79_groupi_g40580(csa_tree_add_51_79_groupi_n_5274 ,csa_tree_add_51_79_groupi_n_5275);
  not csa_tree_add_51_79_groupi_g40581(csa_tree_add_51_79_groupi_n_5270 ,csa_tree_add_51_79_groupi_n_5271);
  not csa_tree_add_51_79_groupi_g40582(csa_tree_add_51_79_groupi_n_5267 ,csa_tree_add_51_79_groupi_n_5268);
  not csa_tree_add_51_79_groupi_g40583(csa_tree_add_51_79_groupi_n_5265 ,csa_tree_add_51_79_groupi_n_5266);
  not csa_tree_add_51_79_groupi_g40584(csa_tree_add_51_79_groupi_n_5259 ,csa_tree_add_51_79_groupi_n_5260);
  not csa_tree_add_51_79_groupi_g40585(csa_tree_add_51_79_groupi_n_5257 ,csa_tree_add_51_79_groupi_n_5258);
  not csa_tree_add_51_79_groupi_g40586(csa_tree_add_51_79_groupi_n_5254 ,csa_tree_add_51_79_groupi_n_5255);
  not csa_tree_add_51_79_groupi_g40587(csa_tree_add_51_79_groupi_n_5243 ,csa_tree_add_51_79_groupi_n_5244);
  not csa_tree_add_51_79_groupi_g40588(csa_tree_add_51_79_groupi_n_5240 ,csa_tree_add_51_79_groupi_n_5241);
  not csa_tree_add_51_79_groupi_g40589(csa_tree_add_51_79_groupi_n_5236 ,csa_tree_add_51_79_groupi_n_5237);
  not csa_tree_add_51_79_groupi_g40590(csa_tree_add_51_79_groupi_n_5228 ,csa_tree_add_51_79_groupi_n_5229);
  not csa_tree_add_51_79_groupi_g40591(csa_tree_add_51_79_groupi_n_5217 ,csa_tree_add_51_79_groupi_n_5216);
  not csa_tree_add_51_79_groupi_g40592(csa_tree_add_51_79_groupi_n_5210 ,csa_tree_add_51_79_groupi_n_5211);
  not csa_tree_add_51_79_groupi_g40593(csa_tree_add_51_79_groupi_n_5207 ,csa_tree_add_51_79_groupi_n_5208);
  not csa_tree_add_51_79_groupi_g40594(csa_tree_add_51_79_groupi_n_5200 ,csa_tree_add_51_79_groupi_n_5201);
  not csa_tree_add_51_79_groupi_g40595(csa_tree_add_51_79_groupi_n_5185 ,csa_tree_add_51_79_groupi_n_5184);
  not csa_tree_add_51_79_groupi_g40596(csa_tree_add_51_79_groupi_n_5178 ,csa_tree_add_51_79_groupi_n_5179);
  not csa_tree_add_51_79_groupi_g40597(csa_tree_add_51_79_groupi_n_5162 ,csa_tree_add_51_79_groupi_n_5163);
  not csa_tree_add_51_79_groupi_g40598(csa_tree_add_51_79_groupi_n_5159 ,csa_tree_add_51_79_groupi_n_5160);
  not csa_tree_add_51_79_groupi_g40599(csa_tree_add_51_79_groupi_n_5154 ,csa_tree_add_51_79_groupi_n_5155);
  or csa_tree_add_51_79_groupi_g40600(csa_tree_add_51_79_groupi_n_5152 ,csa_tree_add_51_79_groupi_n_3313 ,csa_tree_add_51_79_groupi_n_4696);
  and csa_tree_add_51_79_groupi_g40601(csa_tree_add_51_79_groupi_n_5151 ,csa_tree_add_51_79_groupi_n_3832 ,csa_tree_add_51_79_groupi_n_3910);
  and csa_tree_add_51_79_groupi_g40602(csa_tree_add_51_79_groupi_n_5150 ,csa_tree_add_51_79_groupi_n_3833 ,csa_tree_add_51_79_groupi_n_4701);
  and csa_tree_add_51_79_groupi_g40603(csa_tree_add_51_79_groupi_n_5149 ,csa_tree_add_51_79_groupi_n_3830 ,csa_tree_add_51_79_groupi_n_4635);
  or csa_tree_add_51_79_groupi_g40604(csa_tree_add_51_79_groupi_n_5148 ,csa_tree_add_51_79_groupi_n_1176 ,csa_tree_add_51_79_groupi_n_4712);
  or csa_tree_add_51_79_groupi_g40605(csa_tree_add_51_79_groupi_n_5147 ,csa_tree_add_51_79_groupi_n_3311 ,csa_tree_add_51_79_groupi_n_3985);
  and csa_tree_add_51_79_groupi_g40606(csa_tree_add_51_79_groupi_n_5146 ,csa_tree_add_51_79_groupi_n_3317 ,csa_tree_add_51_79_groupi_n_4502);
  or csa_tree_add_51_79_groupi_g40607(csa_tree_add_51_79_groupi_n_5145 ,csa_tree_add_51_79_groupi_n_3315 ,csa_tree_add_51_79_groupi_n_4482);
  or csa_tree_add_51_79_groupi_g40608(csa_tree_add_51_79_groupi_n_5144 ,csa_tree_add_51_79_groupi_n_3319 ,csa_tree_add_51_79_groupi_n_4017);
  or csa_tree_add_51_79_groupi_g40609(csa_tree_add_51_79_groupi_n_5143 ,csa_tree_add_51_79_groupi_n_3321 ,csa_tree_add_51_79_groupi_n_4435);
  or csa_tree_add_51_79_groupi_g40610(csa_tree_add_51_79_groupi_n_5142 ,csa_tree_add_51_79_groupi_n_3316 ,csa_tree_add_51_79_groupi_n_4434);
  or csa_tree_add_51_79_groupi_g40611(csa_tree_add_51_79_groupi_n_5141 ,csa_tree_add_51_79_groupi_n_1178 ,csa_tree_add_51_79_groupi_n_4305);
  and csa_tree_add_51_79_groupi_g40612(csa_tree_add_51_79_groupi_n_5140 ,csa_tree_add_51_79_groupi_n_3191 ,csa_tree_add_51_79_groupi_n_4713);
  and csa_tree_add_51_79_groupi_g40613(csa_tree_add_51_79_groupi_n_5139 ,csa_tree_add_51_79_groupi_n_3193 ,csa_tree_add_51_79_groupi_n_4302);
  or csa_tree_add_51_79_groupi_g40614(csa_tree_add_51_79_groupi_n_5138 ,csa_tree_add_51_79_groupi_n_3331 ,csa_tree_add_51_79_groupi_n_3907);
  or csa_tree_add_51_79_groupi_g40615(csa_tree_add_51_79_groupi_n_5137 ,csa_tree_add_51_79_groupi_n_3318 ,csa_tree_add_51_79_groupi_n_4366);
  or csa_tree_add_51_79_groupi_g40616(csa_tree_add_51_79_groupi_n_5136 ,csa_tree_add_51_79_groupi_n_2555 ,csa_tree_add_51_79_groupi_n_4229);
  and csa_tree_add_51_79_groupi_g40617(csa_tree_add_51_79_groupi_n_5135 ,csa_tree_add_51_79_groupi_n_1174 ,csa_tree_add_51_79_groupi_n_4303);
  or csa_tree_add_51_79_groupi_g40618(csa_tree_add_51_79_groupi_n_5134 ,csa_tree_add_51_79_groupi_n_3329 ,csa_tree_add_51_79_groupi_n_4319);
  or csa_tree_add_51_79_groupi_g40619(csa_tree_add_51_79_groupi_n_5133 ,csa_tree_add_51_79_groupi_n_3323 ,csa_tree_add_51_79_groupi_n_4151);
  or csa_tree_add_51_79_groupi_g40620(csa_tree_add_51_79_groupi_n_5132 ,csa_tree_add_51_79_groupi_n_3332 ,csa_tree_add_51_79_groupi_n_4317);
  and csa_tree_add_51_79_groupi_g40621(csa_tree_add_51_79_groupi_n_5131 ,csa_tree_add_51_79_groupi_n_3831 ,csa_tree_add_51_79_groupi_n_4016);
  or csa_tree_add_51_79_groupi_g40622(csa_tree_add_51_79_groupi_n_5130 ,csa_tree_add_51_79_groupi_n_3314 ,csa_tree_add_51_79_groupi_n_4703);
  or csa_tree_add_51_79_groupi_g40623(csa_tree_add_51_79_groupi_n_5129 ,csa_tree_add_51_79_groupi_n_3325 ,csa_tree_add_51_79_groupi_n_4191);
  or csa_tree_add_51_79_groupi_g40624(csa_tree_add_51_79_groupi_n_5128 ,csa_tree_add_51_79_groupi_n_4226 ,csa_tree_add_51_79_groupi_n_4225);
  or csa_tree_add_51_79_groupi_g40625(csa_tree_add_51_79_groupi_n_5127 ,csa_tree_add_51_79_groupi_n_3310 ,csa_tree_add_51_79_groupi_n_4172);
  or csa_tree_add_51_79_groupi_g40626(csa_tree_add_51_79_groupi_n_5126 ,csa_tree_add_51_79_groupi_n_3192 ,csa_tree_add_51_79_groupi_n_4304);
  or csa_tree_add_51_79_groupi_g40627(csa_tree_add_51_79_groupi_n_5577 ,csa_tree_add_51_79_groupi_n_3346 ,csa_tree_add_51_79_groupi_n_4579);
  and csa_tree_add_51_79_groupi_g40628(csa_tree_add_51_79_groupi_n_5576 ,csa_tree_add_51_79_groupi_n_3514 ,csa_tree_add_51_79_groupi_n_4621);
  and csa_tree_add_51_79_groupi_g40629(csa_tree_add_51_79_groupi_n_5575 ,csa_tree_add_51_79_groupi_n_2998 ,csa_tree_add_51_79_groupi_n_4159);
  and csa_tree_add_51_79_groupi_g40630(csa_tree_add_51_79_groupi_n_5574 ,csa_tree_add_51_79_groupi_n_3154 ,csa_tree_add_51_79_groupi_n_4616);
  and csa_tree_add_51_79_groupi_g40631(csa_tree_add_51_79_groupi_n_5573 ,csa_tree_add_51_79_groupi_n_3501 ,csa_tree_add_51_79_groupi_n_4604);
  and csa_tree_add_51_79_groupi_g40632(csa_tree_add_51_79_groupi_n_5572 ,csa_tree_add_51_79_groupi_n_2951 ,csa_tree_add_51_79_groupi_n_4011);
  and csa_tree_add_51_79_groupi_g40633(csa_tree_add_51_79_groupi_n_5571 ,csa_tree_add_51_79_groupi_n_3859 ,csa_tree_add_51_79_groupi_n_4596);
  and csa_tree_add_51_79_groupi_g40634(csa_tree_add_51_79_groupi_n_5570 ,csa_tree_add_51_79_groupi_n_3094 ,csa_tree_add_51_79_groupi_n_4133);
  and csa_tree_add_51_79_groupi_g40635(csa_tree_add_51_79_groupi_n_5569 ,csa_tree_add_51_79_groupi_n_3485 ,csa_tree_add_51_79_groupi_n_4577);
  and csa_tree_add_51_79_groupi_g40636(csa_tree_add_51_79_groupi_n_5568 ,csa_tree_add_51_79_groupi_n_3387 ,csa_tree_add_51_79_groupi_n_4578);
  and csa_tree_add_51_79_groupi_g40637(csa_tree_add_51_79_groupi_n_5567 ,csa_tree_add_51_79_groupi_n_3132 ,csa_tree_add_51_79_groupi_n_4564);
  and csa_tree_add_51_79_groupi_g40638(csa_tree_add_51_79_groupi_n_5566 ,csa_tree_add_51_79_groupi_n_3468 ,csa_tree_add_51_79_groupi_n_4568);
  and csa_tree_add_51_79_groupi_g40639(csa_tree_add_51_79_groupi_n_5565 ,csa_tree_add_51_79_groupi_n_3563 ,csa_tree_add_51_79_groupi_n_4694);
  and csa_tree_add_51_79_groupi_g40640(csa_tree_add_51_79_groupi_n_5564 ,csa_tree_add_51_79_groupi_n_3009 ,csa_tree_add_51_79_groupi_n_4039);
  and csa_tree_add_51_79_groupi_g40641(csa_tree_add_51_79_groupi_n_5563 ,csa_tree_add_51_79_groupi_n_3379 ,csa_tree_add_51_79_groupi_n_4673);
  and csa_tree_add_51_79_groupi_g40642(csa_tree_add_51_79_groupi_n_5562 ,csa_tree_add_51_79_groupi_n_3403 ,csa_tree_add_51_79_groupi_n_4574);
  and csa_tree_add_51_79_groupi_g40643(csa_tree_add_51_79_groupi_n_5561 ,csa_tree_add_51_79_groupi_n_2885 ,csa_tree_add_51_79_groupi_n_4050);
  and csa_tree_add_51_79_groupi_g40644(csa_tree_add_51_79_groupi_n_5560 ,csa_tree_add_51_79_groupi_n_3451 ,csa_tree_add_51_79_groupi_n_4556);
  and csa_tree_add_51_79_groupi_g40645(csa_tree_add_51_79_groupi_n_5558 ,csa_tree_add_51_79_groupi_n_3337 ,csa_tree_add_51_79_groupi_n_4027);
  and csa_tree_add_51_79_groupi_g40646(csa_tree_add_51_79_groupi_n_5557 ,csa_tree_add_51_79_groupi_n_3369 ,csa_tree_add_51_79_groupi_n_4329);
  and csa_tree_add_51_79_groupi_g40647(csa_tree_add_51_79_groupi_n_5556 ,csa_tree_add_51_79_groupi_n_3460 ,csa_tree_add_51_79_groupi_n_4567);
  or csa_tree_add_51_79_groupi_g40648(csa_tree_add_51_79_groupi_n_5555 ,csa_tree_add_51_79_groupi_n_3846 ,csa_tree_add_51_79_groupi_n_4693);
  and csa_tree_add_51_79_groupi_g40649(csa_tree_add_51_79_groupi_n_5554 ,csa_tree_add_51_79_groupi_n_3022 ,csa_tree_add_51_79_groupi_n_4546);
  and csa_tree_add_51_79_groupi_g40650(csa_tree_add_51_79_groupi_n_5553 ,csa_tree_add_51_79_groupi_n_3019 ,csa_tree_add_51_79_groupi_n_4542);
  and csa_tree_add_51_79_groupi_g40651(csa_tree_add_51_79_groupi_n_5552 ,csa_tree_add_51_79_groupi_n_3004 ,csa_tree_add_51_79_groupi_n_4539);
  and csa_tree_add_51_79_groupi_g40652(csa_tree_add_51_79_groupi_n_5551 ,csa_tree_add_51_79_groupi_n_2950 ,csa_tree_add_51_79_groupi_n_4531);
  and csa_tree_add_51_79_groupi_g40653(csa_tree_add_51_79_groupi_n_5550 ,csa_tree_add_51_79_groupi_n_3023 ,csa_tree_add_51_79_groupi_n_4532);
  and csa_tree_add_51_79_groupi_g40654(csa_tree_add_51_79_groupi_n_5549 ,csa_tree_add_51_79_groupi_n_3864 ,csa_tree_add_51_79_groupi_n_4513);
  and csa_tree_add_51_79_groupi_g40655(csa_tree_add_51_79_groupi_n_5548 ,csa_tree_add_51_79_groupi_n_2984 ,csa_tree_add_51_79_groupi_n_4528);
  and csa_tree_add_51_79_groupi_g40656(csa_tree_add_51_79_groupi_n_5547 ,csa_tree_add_51_79_groupi_n_3013 ,csa_tree_add_51_79_groupi_n_4522);
  and csa_tree_add_51_79_groupi_g40657(csa_tree_add_51_79_groupi_n_5546 ,csa_tree_add_51_79_groupi_n_3474 ,csa_tree_add_51_79_groupi_n_4523);
  and csa_tree_add_51_79_groupi_g40658(csa_tree_add_51_79_groupi_n_5545 ,csa_tree_add_51_79_groupi_n_3038 ,csa_tree_add_51_79_groupi_n_4153);
  and csa_tree_add_51_79_groupi_g40659(csa_tree_add_51_79_groupi_n_5544 ,csa_tree_add_51_79_groupi_n_3861 ,csa_tree_add_51_79_groupi_n_4043);
  and csa_tree_add_51_79_groupi_g40660(csa_tree_add_51_79_groupi_n_5543 ,csa_tree_add_51_79_groupi_n_3422 ,csa_tree_add_51_79_groupi_n_4214);
  and csa_tree_add_51_79_groupi_g40661(csa_tree_add_51_79_groupi_n_5542 ,csa_tree_add_51_79_groupi_n_3456 ,csa_tree_add_51_79_groupi_n_4516);
  and csa_tree_add_51_79_groupi_g40662(csa_tree_add_51_79_groupi_n_5541 ,csa_tree_add_51_79_groupi_n_3086 ,csa_tree_add_51_79_groupi_n_4512);
  and csa_tree_add_51_79_groupi_g40663(csa_tree_add_51_79_groupi_n_5540 ,csa_tree_add_51_79_groupi_n_3416 ,csa_tree_add_51_79_groupi_n_4506);
  and csa_tree_add_51_79_groupi_g40664(csa_tree_add_51_79_groupi_n_5539 ,csa_tree_add_51_79_groupi_n_3343 ,csa_tree_add_51_79_groupi_n_4362);
  and csa_tree_add_51_79_groupi_g40665(csa_tree_add_51_79_groupi_n_5538 ,csa_tree_add_51_79_groupi_n_2926 ,csa_tree_add_51_79_groupi_n_4548);
  and csa_tree_add_51_79_groupi_g40666(csa_tree_add_51_79_groupi_n_5537 ,csa_tree_add_51_79_groupi_n_3426 ,csa_tree_add_51_79_groupi_n_4496);
  and csa_tree_add_51_79_groupi_g40667(csa_tree_add_51_79_groupi_n_5536 ,csa_tree_add_51_79_groupi_n_3434 ,csa_tree_add_51_79_groupi_n_4491);
  and csa_tree_add_51_79_groupi_g40668(csa_tree_add_51_79_groupi_n_5535 ,csa_tree_add_51_79_groupi_n_3473 ,csa_tree_add_51_79_groupi_n_4486);
  and csa_tree_add_51_79_groupi_g40669(csa_tree_add_51_79_groupi_n_5534 ,csa_tree_add_51_79_groupi_n_3847 ,csa_tree_add_51_79_groupi_n_4581);
  and csa_tree_add_51_79_groupi_g40670(csa_tree_add_51_79_groupi_n_5533 ,csa_tree_add_51_79_groupi_n_3544 ,csa_tree_add_51_79_groupi_n_4638);
  and csa_tree_add_51_79_groupi_g40671(csa_tree_add_51_79_groupi_n_5532 ,csa_tree_add_51_79_groupi_n_3455 ,csa_tree_add_51_79_groupi_n_4690);
  and csa_tree_add_51_79_groupi_g40672(csa_tree_add_51_79_groupi_n_5531 ,csa_tree_add_51_79_groupi_n_2962 ,csa_tree_add_51_79_groupi_n_4681);
  and csa_tree_add_51_79_groupi_g40673(csa_tree_add_51_79_groupi_n_5530 ,csa_tree_add_51_79_groupi_n_3439 ,csa_tree_add_51_79_groupi_n_4479);
  and csa_tree_add_51_79_groupi_g40674(csa_tree_add_51_79_groupi_n_5529 ,csa_tree_add_51_79_groupi_n_3550 ,csa_tree_add_51_79_groupi_n_4672);
  and csa_tree_add_51_79_groupi_g40675(csa_tree_add_51_79_groupi_n_5528 ,csa_tree_add_51_79_groupi_n_3371 ,csa_tree_add_51_79_groupi_n_4112);
  and csa_tree_add_51_79_groupi_g40676(csa_tree_add_51_79_groupi_n_5527 ,csa_tree_add_51_79_groupi_n_2996 ,csa_tree_add_51_79_groupi_n_4088);
  and csa_tree_add_51_79_groupi_g40677(csa_tree_add_51_79_groupi_n_5526 ,csa_tree_add_51_79_groupi_n_3419 ,csa_tree_add_51_79_groupi_n_4472);
  and csa_tree_add_51_79_groupi_g40678(csa_tree_add_51_79_groupi_n_5525 ,csa_tree_add_51_79_groupi_n_3554 ,csa_tree_add_51_79_groupi_n_4059);
  and csa_tree_add_51_79_groupi_g40679(csa_tree_add_51_79_groupi_n_5524 ,csa_tree_add_51_79_groupi_n_3479 ,csa_tree_add_51_79_groupi_n_4489);
  and csa_tree_add_51_79_groupi_g40680(csa_tree_add_51_79_groupi_n_5523 ,csa_tree_add_51_79_groupi_n_3517 ,csa_tree_add_51_79_groupi_n_3988);
  or csa_tree_add_51_79_groupi_g40681(csa_tree_add_51_79_groupi_n_5522 ,csa_tree_add_51_79_groupi_n_3866 ,csa_tree_add_51_79_groupi_n_4369);
  and csa_tree_add_51_79_groupi_g40682(csa_tree_add_51_79_groupi_n_5521 ,csa_tree_add_51_79_groupi_n_3342 ,csa_tree_add_51_79_groupi_n_4469);
  and csa_tree_add_51_79_groupi_g40683(csa_tree_add_51_79_groupi_n_5520 ,csa_tree_add_51_79_groupi_n_3105 ,csa_tree_add_51_79_groupi_n_4441);
  and csa_tree_add_51_79_groupi_g40684(csa_tree_add_51_79_groupi_n_5519 ,csa_tree_add_51_79_groupi_n_3359 ,csa_tree_add_51_79_groupi_n_4450);
  and csa_tree_add_51_79_groupi_g40685(csa_tree_add_51_79_groupi_n_5517 ,csa_tree_add_51_79_groupi_n_3082 ,csa_tree_add_51_79_groupi_n_4443);
  and csa_tree_add_51_79_groupi_g40686(csa_tree_add_51_79_groupi_n_5516 ,csa_tree_add_51_79_groupi_n_2973 ,csa_tree_add_51_79_groupi_n_4334);
  and csa_tree_add_51_79_groupi_g40687(csa_tree_add_51_79_groupi_n_5515 ,csa_tree_add_51_79_groupi_n_3398 ,csa_tree_add_51_79_groupi_n_4670);
  and csa_tree_add_51_79_groupi_g40688(csa_tree_add_51_79_groupi_n_5514 ,csa_tree_add_51_79_groupi_n_3465 ,csa_tree_add_51_79_groupi_n_4585);
  and csa_tree_add_51_79_groupi_g40689(csa_tree_add_51_79_groupi_n_5513 ,csa_tree_add_51_79_groupi_n_3538 ,csa_tree_add_51_79_groupi_n_4025);
  and csa_tree_add_51_79_groupi_g40690(csa_tree_add_51_79_groupi_n_5512 ,csa_tree_add_51_79_groupi_n_3143 ,csa_tree_add_51_79_groupi_n_4426);
  and csa_tree_add_51_79_groupi_g40691(csa_tree_add_51_79_groupi_n_5511 ,csa_tree_add_51_79_groupi_n_3457 ,csa_tree_add_51_79_groupi_n_4425);
  and csa_tree_add_51_79_groupi_g40692(csa_tree_add_51_79_groupi_n_5510 ,csa_tree_add_51_79_groupi_n_3014 ,csa_tree_add_51_79_groupi_n_4458);
  and csa_tree_add_51_79_groupi_g40693(csa_tree_add_51_79_groupi_n_5509 ,csa_tree_add_51_79_groupi_n_3859 ,csa_tree_add_51_79_groupi_n_4114);
  and csa_tree_add_51_79_groupi_g40694(csa_tree_add_51_79_groupi_n_5508 ,csa_tree_add_51_79_groupi_n_3580 ,csa_tree_add_51_79_groupi_n_4697);
  and csa_tree_add_51_79_groupi_g40695(csa_tree_add_51_79_groupi_n_5507 ,csa_tree_add_51_79_groupi_n_2907 ,csa_tree_add_51_79_groupi_n_4412);
  and csa_tree_add_51_79_groupi_g40696(csa_tree_add_51_79_groupi_n_5506 ,csa_tree_add_51_79_groupi_n_2949 ,csa_tree_add_51_79_groupi_n_4409);
  and csa_tree_add_51_79_groupi_g40697(csa_tree_add_51_79_groupi_n_5505 ,csa_tree_add_51_79_groupi_n_3061 ,csa_tree_add_51_79_groupi_n_4408);
  and csa_tree_add_51_79_groupi_g40698(csa_tree_add_51_79_groupi_n_5504 ,csa_tree_add_51_79_groupi_n_3578 ,csa_tree_add_51_79_groupi_n_4406);
  and csa_tree_add_51_79_groupi_g40699(csa_tree_add_51_79_groupi_n_5503 ,csa_tree_add_51_79_groupi_n_3518 ,csa_tree_add_51_79_groupi_n_4397);
  and csa_tree_add_51_79_groupi_g40700(csa_tree_add_51_79_groupi_n_5502 ,csa_tree_add_51_79_groupi_n_3470 ,csa_tree_add_51_79_groupi_n_4464);
  and csa_tree_add_51_79_groupi_g40701(csa_tree_add_51_79_groupi_n_5501 ,csa_tree_add_51_79_groupi_n_3104 ,csa_tree_add_51_79_groupi_n_4395);
  and csa_tree_add_51_79_groupi_g40702(csa_tree_add_51_79_groupi_n_5500 ,csa_tree_add_51_79_groupi_n_3033 ,csa_tree_add_51_79_groupi_n_4018);
  and csa_tree_add_51_79_groupi_g40703(csa_tree_add_51_79_groupi_n_5499 ,csa_tree_add_51_79_groupi_n_3842 ,csa_tree_add_51_79_groupi_n_3998);
  and csa_tree_add_51_79_groupi_g40704(csa_tree_add_51_79_groupi_n_5498 ,csa_tree_add_51_79_groupi_n_3528 ,csa_tree_add_51_79_groupi_n_4371);
  or csa_tree_add_51_79_groupi_g40705(csa_tree_add_51_79_groupi_n_5497 ,csa_tree_add_51_79_groupi_n_3360 ,csa_tree_add_51_79_groupi_n_3995);
  and csa_tree_add_51_79_groupi_g40706(csa_tree_add_51_79_groupi_n_5496 ,csa_tree_add_51_79_groupi_n_3556 ,csa_tree_add_51_79_groupi_n_4384);
  and csa_tree_add_51_79_groupi_g40707(csa_tree_add_51_79_groupi_n_5495 ,csa_tree_add_51_79_groupi_n_3155 ,csa_tree_add_51_79_groupi_n_4666);
  and csa_tree_add_51_79_groupi_g40708(csa_tree_add_51_79_groupi_n_5494 ,csa_tree_add_51_79_groupi_n_2989 ,csa_tree_add_51_79_groupi_n_4558);
  and csa_tree_add_51_79_groupi_g40709(csa_tree_add_51_79_groupi_n_5493 ,csa_tree_add_51_79_groupi_n_3628 ,csa_tree_add_51_79_groupi_n_4376);
  and csa_tree_add_51_79_groupi_g40710(csa_tree_add_51_79_groupi_n_5492 ,csa_tree_add_51_79_groupi_n_3539 ,csa_tree_add_51_79_groupi_n_4662);
  and csa_tree_add_51_79_groupi_g40711(csa_tree_add_51_79_groupi_n_5491 ,csa_tree_add_51_79_groupi_n_3644 ,csa_tree_add_51_79_groupi_n_4432);
  and csa_tree_add_51_79_groupi_g40712(csa_tree_add_51_79_groupi_n_5490 ,csa_tree_add_51_79_groupi_n_3401 ,csa_tree_add_51_79_groupi_n_4657);
  and csa_tree_add_51_79_groupi_g40713(csa_tree_add_51_79_groupi_n_5489 ,csa_tree_add_51_79_groupi_n_3541 ,csa_tree_add_51_79_groupi_n_4656);
  and csa_tree_add_51_79_groupi_g40714(csa_tree_add_51_79_groupi_n_5488 ,csa_tree_add_51_79_groupi_n_3502 ,csa_tree_add_51_79_groupi_n_4658);
  and csa_tree_add_51_79_groupi_g40715(csa_tree_add_51_79_groupi_n_5487 ,csa_tree_add_51_79_groupi_n_3119 ,csa_tree_add_51_79_groupi_n_4086);
  and csa_tree_add_51_79_groupi_g40716(csa_tree_add_51_79_groupi_n_5486 ,csa_tree_add_51_79_groupi_n_3459 ,csa_tree_add_51_79_groupi_n_4356);
  and csa_tree_add_51_79_groupi_g40717(csa_tree_add_51_79_groupi_n_5485 ,csa_tree_add_51_79_groupi_n_3508 ,csa_tree_add_51_79_groupi_n_4340);
  and csa_tree_add_51_79_groupi_g40718(csa_tree_add_51_79_groupi_n_5484 ,csa_tree_add_51_79_groupi_n_3336 ,csa_tree_add_51_79_groupi_n_4338);
  and csa_tree_add_51_79_groupi_g40719(csa_tree_add_51_79_groupi_n_5483 ,csa_tree_add_51_79_groupi_n_3081 ,csa_tree_add_51_79_groupi_n_4328);
  and csa_tree_add_51_79_groupi_g40720(csa_tree_add_51_79_groupi_n_5482 ,csa_tree_add_51_79_groupi_n_3138 ,csa_tree_add_51_79_groupi_n_4324);
  and csa_tree_add_51_79_groupi_g40721(csa_tree_add_51_79_groupi_n_5481 ,csa_tree_add_51_79_groupi_n_2923 ,csa_tree_add_51_79_groupi_n_4497);
  and csa_tree_add_51_79_groupi_g40722(csa_tree_add_51_79_groupi_n_5480 ,csa_tree_add_51_79_groupi_n_3131 ,csa_tree_add_51_79_groupi_n_4648);
  and csa_tree_add_51_79_groupi_g40723(csa_tree_add_51_79_groupi_n_5479 ,csa_tree_add_51_79_groupi_n_3351 ,csa_tree_add_51_79_groupi_n_4647);
  and csa_tree_add_51_79_groupi_g40724(csa_tree_add_51_79_groupi_n_5478 ,csa_tree_add_51_79_groupi_n_3135 ,csa_tree_add_51_79_groupi_n_4318);
  and csa_tree_add_51_79_groupi_g40725(csa_tree_add_51_79_groupi_n_5477 ,csa_tree_add_51_79_groupi_n_3148 ,csa_tree_add_51_79_groupi_n_4087);
  and csa_tree_add_51_79_groupi_g40726(csa_tree_add_51_79_groupi_n_5476 ,csa_tree_add_51_79_groupi_n_3845 ,csa_tree_add_51_79_groupi_n_4165);
  and csa_tree_add_51_79_groupi_g40727(csa_tree_add_51_79_groupi_n_5475 ,csa_tree_add_51_79_groupi_n_3129 ,csa_tree_add_51_79_groupi_n_4594);
  and csa_tree_add_51_79_groupi_g40728(csa_tree_add_51_79_groupi_n_5474 ,csa_tree_add_51_79_groupi_n_3016 ,csa_tree_add_51_79_groupi_n_4129);
  and csa_tree_add_51_79_groupi_g40729(csa_tree_add_51_79_groupi_n_5473 ,csa_tree_add_51_79_groupi_n_3087 ,csa_tree_add_51_79_groupi_n_4310);
  and csa_tree_add_51_79_groupi_g40730(csa_tree_add_51_79_groupi_n_5472 ,csa_tree_add_51_79_groupi_n_2982 ,csa_tree_add_51_79_groupi_n_4520);
  and csa_tree_add_51_79_groupi_g40731(csa_tree_add_51_79_groupi_n_5471 ,csa_tree_add_51_79_groupi_n_3520 ,csa_tree_add_51_79_groupi_n_4642);
  and csa_tree_add_51_79_groupi_g40732(csa_tree_add_51_79_groupi_n_5470 ,csa_tree_add_51_79_groupi_n_3124 ,csa_tree_add_51_79_groupi_n_4223);
  and csa_tree_add_51_79_groupi_g40733(csa_tree_add_51_79_groupi_n_5469 ,csa_tree_add_51_79_groupi_n_2927 ,csa_tree_add_51_79_groupi_n_4221);
  and csa_tree_add_51_79_groupi_g40734(csa_tree_add_51_79_groupi_n_5468 ,csa_tree_add_51_79_groupi_n_3872 ,csa_tree_add_51_79_groupi_n_3903);
  and csa_tree_add_51_79_groupi_g40735(csa_tree_add_51_79_groupi_n_5467 ,csa_tree_add_51_79_groupi_n_2997 ,csa_tree_add_51_79_groupi_n_4212);
  and csa_tree_add_51_79_groupi_g40736(csa_tree_add_51_79_groupi_n_5466 ,csa_tree_add_51_79_groupi_n_2961 ,csa_tree_add_51_79_groupi_n_4213);
  and csa_tree_add_51_79_groupi_g40737(csa_tree_add_51_79_groupi_n_5465 ,csa_tree_add_51_79_groupi_n_2974 ,csa_tree_add_51_79_groupi_n_4200);
  and csa_tree_add_51_79_groupi_g40738(csa_tree_add_51_79_groupi_n_5464 ,csa_tree_add_51_79_groupi_n_2994 ,csa_tree_add_51_79_groupi_n_3906);
  and csa_tree_add_51_79_groupi_g40739(csa_tree_add_51_79_groupi_n_5463 ,csa_tree_add_51_79_groupi_n_2953 ,csa_tree_add_51_79_groupi_n_4636);
  and csa_tree_add_51_79_groupi_g40740(csa_tree_add_51_79_groupi_n_5462 ,csa_tree_add_51_79_groupi_n_3570 ,csa_tree_add_51_79_groupi_n_4193);
  or csa_tree_add_51_79_groupi_g40741(csa_tree_add_51_79_groupi_n_5461 ,csa_tree_add_51_79_groupi_n_3870 ,csa_tree_add_51_79_groupi_n_4643);
  and csa_tree_add_51_79_groupi_g40742(csa_tree_add_51_79_groupi_n_5460 ,csa_tree_add_51_79_groupi_n_3577 ,csa_tree_add_51_79_groupi_n_4152);
  and csa_tree_add_51_79_groupi_g40743(csa_tree_add_51_79_groupi_n_5459 ,csa_tree_add_51_79_groupi_n_3365 ,csa_tree_add_51_79_groupi_n_4135);
  and csa_tree_add_51_79_groupi_g40744(csa_tree_add_51_79_groupi_n_5458 ,csa_tree_add_51_79_groupi_n_2967 ,csa_tree_add_51_79_groupi_n_4054);
  and csa_tree_add_51_79_groupi_g40745(csa_tree_add_51_79_groupi_n_5457 ,csa_tree_add_51_79_groupi_n_3112 ,csa_tree_add_51_79_groupi_n_4314);
  and csa_tree_add_51_79_groupi_g40746(csa_tree_add_51_79_groupi_n_5456 ,csa_tree_add_51_79_groupi_n_3026 ,csa_tree_add_51_79_groupi_n_4177);
  and csa_tree_add_51_79_groupi_g40747(csa_tree_add_51_79_groupi_n_5455 ,csa_tree_add_51_79_groupi_n_3850 ,csa_tree_add_51_79_groupi_n_4202);
  and csa_tree_add_51_79_groupi_g40748(csa_tree_add_51_79_groupi_n_5453 ,csa_tree_add_51_79_groupi_n_3855 ,csa_tree_add_51_79_groupi_n_4627);
  and csa_tree_add_51_79_groupi_g40749(csa_tree_add_51_79_groupi_n_5452 ,csa_tree_add_51_79_groupi_n_3659 ,csa_tree_add_51_79_groupi_n_4684);
  or csa_tree_add_51_79_groupi_g40750(csa_tree_add_51_79_groupi_n_5451 ,csa_tree_add_51_79_groupi_n_3340 ,csa_tree_add_51_79_groupi_n_4057);
  and csa_tree_add_51_79_groupi_g40751(csa_tree_add_51_79_groupi_n_5450 ,csa_tree_add_51_79_groupi_n_3080 ,csa_tree_add_51_79_groupi_n_4600);
  and csa_tree_add_51_79_groupi_g40752(csa_tree_add_51_79_groupi_n_5449 ,csa_tree_add_51_79_groupi_n_3856 ,csa_tree_add_51_79_groupi_n_4466);
  and csa_tree_add_51_79_groupi_g40753(csa_tree_add_51_79_groupi_n_5448 ,csa_tree_add_51_79_groupi_n_3043 ,csa_tree_add_51_79_groupi_n_4049);
  and csa_tree_add_51_79_groupi_g40754(csa_tree_add_51_79_groupi_n_5447 ,csa_tree_add_51_79_groupi_n_3489 ,csa_tree_add_51_79_groupi_n_4630);
  or csa_tree_add_51_79_groupi_g40755(csa_tree_add_51_79_groupi_n_5446 ,csa_tree_add_51_79_groupi_n_3362 ,csa_tree_add_51_79_groupi_n_4561);
  and csa_tree_add_51_79_groupi_g40756(csa_tree_add_51_79_groupi_n_5445 ,csa_tree_add_51_79_groupi_n_3072 ,csa_tree_add_51_79_groupi_n_4158);
  and csa_tree_add_51_79_groupi_g40757(csa_tree_add_51_79_groupi_n_5443 ,csa_tree_add_51_79_groupi_n_3337 ,csa_tree_add_51_79_groupi_n_4181);
  and csa_tree_add_51_79_groupi_g40758(csa_tree_add_51_79_groupi_n_5442 ,csa_tree_add_51_79_groupi_n_3109 ,csa_tree_add_51_79_groupi_n_4433);
  and csa_tree_add_51_79_groupi_g40759(csa_tree_add_51_79_groupi_n_5441 ,csa_tree_add_51_79_groupi_n_2921 ,csa_tree_add_51_79_groupi_n_3982);
  and csa_tree_add_51_79_groupi_g40760(csa_tree_add_51_79_groupi_n_5440 ,csa_tree_add_51_79_groupi_n_3055 ,csa_tree_add_51_79_groupi_n_4156);
  and csa_tree_add_51_79_groupi_g40761(csa_tree_add_51_79_groupi_n_5439 ,csa_tree_add_51_79_groupi_n_3561 ,csa_tree_add_51_79_groupi_n_4211);
  and csa_tree_add_51_79_groupi_g40762(csa_tree_add_51_79_groupi_n_5438 ,csa_tree_add_51_79_groupi_n_3001 ,csa_tree_add_51_79_groupi_n_4147);
  and csa_tree_add_51_79_groupi_g40763(csa_tree_add_51_79_groupi_n_5437 ,csa_tree_add_51_79_groupi_n_3056 ,csa_tree_add_51_79_groupi_n_3892);
  and csa_tree_add_51_79_groupi_g40764(csa_tree_add_51_79_groupi_n_5436 ,csa_tree_add_51_79_groupi_n_3041 ,csa_tree_add_51_79_groupi_n_4138);
  and csa_tree_add_51_79_groupi_g40765(csa_tree_add_51_79_groupi_n_5435 ,csa_tree_add_51_79_groupi_n_3339 ,csa_tree_add_51_79_groupi_n_4331);
  and csa_tree_add_51_79_groupi_g40766(csa_tree_add_51_79_groupi_n_5434 ,csa_tree_add_51_79_groupi_n_3355 ,csa_tree_add_51_79_groupi_n_4569);
  and csa_tree_add_51_79_groupi_g40767(csa_tree_add_51_79_groupi_n_5433 ,csa_tree_add_51_79_groupi_n_3507 ,csa_tree_add_51_79_groupi_n_4612);
  and csa_tree_add_51_79_groupi_g40768(csa_tree_add_51_79_groupi_n_5432 ,csa_tree_add_51_79_groupi_n_3848 ,csa_tree_add_51_79_groupi_n_4677);
  and csa_tree_add_51_79_groupi_g40769(csa_tree_add_51_79_groupi_n_5430 ,csa_tree_add_51_79_groupi_n_3367 ,csa_tree_add_51_79_groupi_n_4688);
  and csa_tree_add_51_79_groupi_g40770(csa_tree_add_51_79_groupi_n_5429 ,csa_tree_add_51_79_groupi_n_2945 ,csa_tree_add_51_79_groupi_n_3986);
  and csa_tree_add_51_79_groupi_g40771(csa_tree_add_51_79_groupi_n_5428 ,csa_tree_add_51_79_groupi_n_3140 ,csa_tree_add_51_79_groupi_n_4659);
  and csa_tree_add_51_79_groupi_g40772(csa_tree_add_51_79_groupi_n_5427 ,csa_tree_add_51_79_groupi_n_2968 ,csa_tree_add_51_79_groupi_n_4608);
  and csa_tree_add_51_79_groupi_g40773(csa_tree_add_51_79_groupi_n_5426 ,csa_tree_add_51_79_groupi_n_3865 ,csa_tree_add_51_79_groupi_n_4660);
  and csa_tree_add_51_79_groupi_g40774(csa_tree_add_51_79_groupi_n_5424 ,csa_tree_add_51_79_groupi_n_3027 ,csa_tree_add_51_79_groupi_n_4605);
  and csa_tree_add_51_79_groupi_g40775(csa_tree_add_51_79_groupi_n_5423 ,csa_tree_add_51_79_groupi_n_3113 ,csa_tree_add_51_79_groupi_n_4444);
  and csa_tree_add_51_79_groupi_g40776(csa_tree_add_51_79_groupi_n_5421 ,csa_tree_add_51_79_groupi_n_3096 ,csa_tree_add_51_79_groupi_n_4601);
  and csa_tree_add_51_79_groupi_g40777(csa_tree_add_51_79_groupi_n_5420 ,csa_tree_add_51_79_groupi_n_3543 ,csa_tree_add_51_79_groupi_n_4467);
  and csa_tree_add_51_79_groupi_g40778(csa_tree_add_51_79_groupi_n_5419 ,csa_tree_add_51_79_groupi_n_2979 ,csa_tree_add_51_79_groupi_n_4175);
  or csa_tree_add_51_79_groupi_g40779(csa_tree_add_51_79_groupi_n_5417 ,csa_tree_add_51_79_groupi_n_3375 ,csa_tree_add_51_79_groupi_n_4062);
  and csa_tree_add_51_79_groupi_g40780(csa_tree_add_51_79_groupi_n_5416 ,csa_tree_add_51_79_groupi_n_3871 ,csa_tree_add_51_79_groupi_n_4453);
  and csa_tree_add_51_79_groupi_g40781(csa_tree_add_51_79_groupi_n_5414 ,csa_tree_add_51_79_groupi_n_3654 ,csa_tree_add_51_79_groupi_n_4591);
  and csa_tree_add_51_79_groupi_g40782(csa_tree_add_51_79_groupi_n_5413 ,csa_tree_add_51_79_groupi_n_3402 ,csa_tree_add_51_79_groupi_n_4476);
  and csa_tree_add_51_79_groupi_g40783(csa_tree_add_51_79_groupi_n_5412 ,csa_tree_add_51_79_groupi_n_3091 ,csa_tree_add_51_79_groupi_n_4566);
  and csa_tree_add_51_79_groupi_g40784(csa_tree_add_51_79_groupi_n_5411 ,csa_tree_add_51_79_groupi_n_3521 ,csa_tree_add_51_79_groupi_n_4140);
  and csa_tree_add_51_79_groupi_g40785(csa_tree_add_51_79_groupi_n_5410 ,csa_tree_add_51_79_groupi_n_3512 ,csa_tree_add_51_79_groupi_n_4587);
  and csa_tree_add_51_79_groupi_g40786(csa_tree_add_51_79_groupi_n_5408 ,csa_tree_add_51_79_groupi_n_3486 ,csa_tree_add_51_79_groupi_n_4582);
  and csa_tree_add_51_79_groupi_g40787(csa_tree_add_51_79_groupi_n_5407 ,csa_tree_add_51_79_groupi_n_3378 ,csa_tree_add_51_79_groupi_n_4580);
  and csa_tree_add_51_79_groupi_g40788(csa_tree_add_51_79_groupi_n_5406 ,csa_tree_add_51_79_groupi_n_3552 ,csa_tree_add_51_79_groupi_n_4678);
  and csa_tree_add_51_79_groupi_g40789(csa_tree_add_51_79_groupi_n_5405 ,csa_tree_add_51_79_groupi_n_2948 ,csa_tree_add_51_79_groupi_n_4655);
  and csa_tree_add_51_79_groupi_g40790(csa_tree_add_51_79_groupi_n_5404 ,csa_tree_add_51_79_groupi_n_3869 ,csa_tree_add_51_79_groupi_n_4040);
  and csa_tree_add_51_79_groupi_g40791(csa_tree_add_51_79_groupi_n_5403 ,csa_tree_add_51_79_groupi_n_3341 ,csa_tree_add_51_79_groupi_n_4128);
  and csa_tree_add_51_79_groupi_g40792(csa_tree_add_51_79_groupi_n_5401 ,csa_tree_add_51_79_groupi_n_3553 ,csa_tree_add_51_79_groupi_n_4446);
  and csa_tree_add_51_79_groupi_g40793(csa_tree_add_51_79_groupi_n_5399 ,csa_tree_add_51_79_groupi_n_3415 ,csa_tree_add_51_79_groupi_n_4051);
  and csa_tree_add_51_79_groupi_g40794(csa_tree_add_51_79_groupi_n_5397 ,csa_tree_add_51_79_groupi_n_3076 ,csa_tree_add_51_79_groupi_n_4315);
  and csa_tree_add_51_79_groupi_g40795(csa_tree_add_51_79_groupi_n_5396 ,csa_tree_add_51_79_groupi_n_3872 ,csa_tree_add_51_79_groupi_n_4699);
  and csa_tree_add_51_79_groupi_g40796(csa_tree_add_51_79_groupi_n_5394 ,csa_tree_add_51_79_groupi_n_3394 ,csa_tree_add_51_79_groupi_n_4571);
  and csa_tree_add_51_79_groupi_g40797(csa_tree_add_51_79_groupi_n_5393 ,csa_tree_add_51_79_groupi_n_3383 ,csa_tree_add_51_79_groupi_n_4219);
  and csa_tree_add_51_79_groupi_g40798(csa_tree_add_51_79_groupi_n_5392 ,csa_tree_add_51_79_groupi_n_3348 ,csa_tree_add_51_79_groupi_n_4463);
  and csa_tree_add_51_79_groupi_g40799(csa_tree_add_51_79_groupi_n_5391 ,csa_tree_add_51_79_groupi_n_3412 ,csa_tree_add_51_79_groupi_n_4654);
  and csa_tree_add_51_79_groupi_g40800(csa_tree_add_51_79_groupi_n_5390 ,csa_tree_add_51_79_groupi_n_3345 ,csa_tree_add_51_79_groupi_n_4094);
  and csa_tree_add_51_79_groupi_g40801(csa_tree_add_51_79_groupi_n_5388 ,csa_tree_add_51_79_groupi_n_3437 ,csa_tree_add_51_79_groupi_n_4438);
  and csa_tree_add_51_79_groupi_g40802(csa_tree_add_51_79_groupi_n_5386 ,csa_tree_add_51_79_groupi_n_3115 ,csa_tree_add_51_79_groupi_n_4188);
  and csa_tree_add_51_79_groupi_g40803(csa_tree_add_51_79_groupi_n_5385 ,csa_tree_add_51_79_groupi_n_3540 ,csa_tree_add_51_79_groupi_n_4653);
  and csa_tree_add_51_79_groupi_g40804(csa_tree_add_51_79_groupi_n_5384 ,csa_tree_add_51_79_groupi_n_3537 ,csa_tree_add_51_79_groupi_n_4650);
  and csa_tree_add_51_79_groupi_g40805(csa_tree_add_51_79_groupi_n_5383 ,csa_tree_add_51_79_groupi_n_3095 ,csa_tree_add_51_79_groupi_n_4430);
  and csa_tree_add_51_79_groupi_g40806(csa_tree_add_51_79_groupi_n_5382 ,csa_tree_add_51_79_groupi_n_3021 ,csa_tree_add_51_79_groupi_n_4651);
  and csa_tree_add_51_79_groupi_g40807(csa_tree_add_51_79_groupi_n_5381 ,csa_tree_add_51_79_groupi_n_3054 ,csa_tree_add_51_79_groupi_n_4428);
  and csa_tree_add_51_79_groupi_g40808(csa_tree_add_51_79_groupi_n_5379 ,csa_tree_add_51_79_groupi_n_3461 ,csa_tree_add_51_79_groupi_n_4427);
  and csa_tree_add_51_79_groupi_g40809(csa_tree_add_51_79_groupi_n_5378 ,csa_tree_add_51_79_groupi_n_3134 ,csa_tree_add_51_79_groupi_n_4649);
  and csa_tree_add_51_79_groupi_g40810(csa_tree_add_51_79_groupi_n_5377 ,csa_tree_add_51_79_groupi_n_3432 ,csa_tree_add_51_79_groupi_n_4676);
  and csa_tree_add_51_79_groupi_g40811(csa_tree_add_51_79_groupi_n_5376 ,csa_tree_add_51_79_groupi_n_3499 ,csa_tree_add_51_79_groupi_n_4560);
  and csa_tree_add_51_79_groupi_g40812(csa_tree_add_51_79_groupi_n_5375 ,csa_tree_add_51_79_groupi_n_3480 ,csa_tree_add_51_79_groupi_n_4559);
  and csa_tree_add_51_79_groupi_g40813(csa_tree_add_51_79_groupi_n_5373 ,csa_tree_add_51_79_groupi_n_3579 ,csa_tree_add_51_79_groupi_n_4459);
  and csa_tree_add_51_79_groupi_g40814(csa_tree_add_51_79_groupi_n_5372 ,csa_tree_add_51_79_groupi_n_2988 ,csa_tree_add_51_79_groupi_n_4423);
  and csa_tree_add_51_79_groupi_g40815(csa_tree_add_51_79_groupi_n_5370 ,csa_tree_add_51_79_groupi_n_3478 ,csa_tree_add_51_79_groupi_n_4420);
  and csa_tree_add_51_79_groupi_g40816(csa_tree_add_51_79_groupi_n_5368 ,csa_tree_add_51_79_groupi_n_3139 ,csa_tree_add_51_79_groupi_n_4419);
  and csa_tree_add_51_79_groupi_g40817(csa_tree_add_51_79_groupi_n_5367 ,csa_tree_add_51_79_groupi_n_3490 ,csa_tree_add_51_79_groupi_n_4413);
  and csa_tree_add_51_79_groupi_g40818(csa_tree_add_51_79_groupi_n_5365 ,csa_tree_add_51_79_groupi_n_2955 ,csa_tree_add_51_79_groupi_n_4414);
  and csa_tree_add_51_79_groupi_g40819(csa_tree_add_51_79_groupi_n_5364 ,csa_tree_add_51_79_groupi_n_3869 ,csa_tree_add_51_79_groupi_n_4637);
  and csa_tree_add_51_79_groupi_g40820(csa_tree_add_51_79_groupi_n_5362 ,csa_tree_add_51_79_groupi_n_3861 ,csa_tree_add_51_79_groupi_n_4641);
  and csa_tree_add_51_79_groupi_g40821(csa_tree_add_51_79_groupi_n_5361 ,csa_tree_add_51_79_groupi_n_2899 ,csa_tree_add_51_79_groupi_n_4410);
  and csa_tree_add_51_79_groupi_g40822(csa_tree_add_51_79_groupi_n_5360 ,csa_tree_add_51_79_groupi_n_3533 ,csa_tree_add_51_79_groupi_n_4386);
  and csa_tree_add_51_79_groupi_g40823(csa_tree_add_51_79_groupi_n_5358 ,csa_tree_add_51_79_groupi_n_3494 ,csa_tree_add_51_79_groupi_n_3989);
  and csa_tree_add_51_79_groupi_g40824(csa_tree_add_51_79_groupi_n_5357 ,csa_tree_add_51_79_groupi_n_3496 ,csa_tree_add_51_79_groupi_n_4013);
  and csa_tree_add_51_79_groupi_g40825(csa_tree_add_51_79_groupi_n_5356 ,csa_tree_add_51_79_groupi_n_3445 ,csa_tree_add_51_79_groupi_n_4313);
  and csa_tree_add_51_79_groupi_g40826(csa_tree_add_51_79_groupi_n_5355 ,csa_tree_add_51_79_groupi_n_3562 ,csa_tree_add_51_79_groupi_n_4646);
  and csa_tree_add_51_79_groupi_g40827(csa_tree_add_51_79_groupi_n_5353 ,csa_tree_add_51_79_groupi_n_2971 ,csa_tree_add_51_79_groupi_n_4405);
  and csa_tree_add_51_79_groupi_g40828(csa_tree_add_51_79_groupi_n_5352 ,csa_tree_add_51_79_groupi_n_3347 ,csa_tree_add_51_79_groupi_n_4349);
  and csa_tree_add_51_79_groupi_g40829(csa_tree_add_51_79_groupi_n_5350 ,csa_tree_add_51_79_groupi_n_3048 ,csa_tree_add_51_79_groupi_n_4398);
  and csa_tree_add_51_79_groupi_g40830(csa_tree_add_51_79_groupi_n_5349 ,csa_tree_add_51_79_groupi_n_3558 ,csa_tree_add_51_79_groupi_n_4421);
  and csa_tree_add_51_79_groupi_g40831(csa_tree_add_51_79_groupi_n_5348 ,csa_tree_add_51_79_groupi_n_3414 ,csa_tree_add_51_79_groupi_n_4555);
  and csa_tree_add_51_79_groupi_g40832(csa_tree_add_51_79_groupi_n_5347 ,csa_tree_add_51_79_groupi_n_3852 ,csa_tree_add_51_79_groupi_n_4107);
  and csa_tree_add_51_79_groupi_g40833(csa_tree_add_51_79_groupi_n_5345 ,csa_tree_add_51_79_groupi_n_3565 ,csa_tree_add_51_79_groupi_n_4553);
  and csa_tree_add_51_79_groupi_g40834(csa_tree_add_51_79_groupi_n_5344 ,csa_tree_add_51_79_groupi_n_3530 ,csa_tree_add_51_79_groupi_n_4551);
  and csa_tree_add_51_79_groupi_g40835(csa_tree_add_51_79_groupi_n_5343 ,csa_tree_add_51_79_groupi_n_3524 ,csa_tree_add_51_79_groupi_n_4346);
  and csa_tree_add_51_79_groupi_g40836(csa_tree_add_51_79_groupi_n_5341 ,csa_tree_add_51_79_groupi_n_3443 ,csa_tree_add_51_79_groupi_n_4626);
  and csa_tree_add_51_79_groupi_g40837(csa_tree_add_51_79_groupi_n_5340 ,csa_tree_add_51_79_groupi_n_3527 ,csa_tree_add_51_79_groupi_n_4588);
  and csa_tree_add_51_79_groupi_g40838(csa_tree_add_51_79_groupi_n_5339 ,csa_tree_add_51_79_groupi_n_2890 ,csa_tree_add_51_79_groupi_n_4589);
  and csa_tree_add_51_79_groupi_g40839(csa_tree_add_51_79_groupi_n_5338 ,csa_tree_add_51_79_groupi_n_3133 ,csa_tree_add_51_79_groupi_n_4077);
  and csa_tree_add_51_79_groupi_g40840(csa_tree_add_51_79_groupi_n_5337 ,csa_tree_add_51_79_groupi_n_3555 ,csa_tree_add_51_79_groupi_n_4385);
  and csa_tree_add_51_79_groupi_g40841(csa_tree_add_51_79_groupi_n_5335 ,csa_tree_add_51_79_groupi_n_3338 ,csa_tree_add_51_79_groupi_n_4639);
  and csa_tree_add_51_79_groupi_g40842(csa_tree_add_51_79_groupi_n_5334 ,csa_tree_add_51_79_groupi_n_3392 ,csa_tree_add_51_79_groupi_n_4030);
  and csa_tree_add_51_79_groupi_g40843(csa_tree_add_51_79_groupi_n_5333 ,csa_tree_add_51_79_groupi_n_3462 ,csa_tree_add_51_79_groupi_n_4379);
  and csa_tree_add_51_79_groupi_g40844(csa_tree_add_51_79_groupi_n_5332 ,csa_tree_add_51_79_groupi_n_3547 ,csa_tree_add_51_79_groupi_n_4669);
  and csa_tree_add_51_79_groupi_g40845(csa_tree_add_51_79_groupi_n_5330 ,csa_tree_add_51_79_groupi_n_3029 ,csa_tree_add_51_79_groupi_n_4066);
  and csa_tree_add_51_79_groupi_g40846(csa_tree_add_51_79_groupi_n_5329 ,csa_tree_add_51_79_groupi_n_3011 ,csa_tree_add_51_79_groupi_n_4174);
  and csa_tree_add_51_79_groupi_g40847(csa_tree_add_51_79_groupi_n_5328 ,csa_tree_add_51_79_groupi_n_3103 ,csa_tree_add_51_79_groupi_n_4375);
  and csa_tree_add_51_79_groupi_g40848(csa_tree_add_51_79_groupi_n_5326 ,csa_tree_add_51_79_groupi_n_3569 ,csa_tree_add_51_79_groupi_n_4373);
  and csa_tree_add_51_79_groupi_g40849(csa_tree_add_51_79_groupi_n_5325 ,csa_tree_add_51_79_groupi_n_3399 ,csa_tree_add_51_79_groupi_n_4671);
  and csa_tree_add_51_79_groupi_g40850(csa_tree_add_51_79_groupi_n_5324 ,csa_tree_add_51_79_groupi_n_2946 ,csa_tree_add_51_79_groupi_n_4545);
  and csa_tree_add_51_79_groupi_g40851(csa_tree_add_51_79_groupi_n_5323 ,csa_tree_add_51_79_groupi_n_3867 ,csa_tree_add_51_79_groupi_n_4113);
  and csa_tree_add_51_79_groupi_g40852(csa_tree_add_51_79_groupi_n_5321 ,csa_tree_add_51_79_groupi_n_3851 ,csa_tree_add_51_79_groupi_n_4572);
  and csa_tree_add_51_79_groupi_g40853(csa_tree_add_51_79_groupi_n_5320 ,csa_tree_add_51_79_groupi_n_3097 ,csa_tree_add_51_79_groupi_n_4547);
  and csa_tree_add_51_79_groupi_g40854(csa_tree_add_51_79_groupi_n_5319 ,csa_tree_add_51_79_groupi_n_3482 ,csa_tree_add_51_79_groupi_n_4424);
  and csa_tree_add_51_79_groupi_g40855(csa_tree_add_51_79_groupi_n_5318 ,csa_tree_add_51_79_groupi_n_3436 ,csa_tree_add_51_79_groupi_n_4540);
  and csa_tree_add_51_79_groupi_g40856(csa_tree_add_51_79_groupi_n_5317 ,csa_tree_add_51_79_groupi_n_3845 ,csa_tree_add_51_79_groupi_n_4521);
  and csa_tree_add_51_79_groupi_g40857(csa_tree_add_51_79_groupi_n_5315 ,csa_tree_add_51_79_groupi_n_3361 ,csa_tree_add_51_79_groupi_n_3991);
  and csa_tree_add_51_79_groupi_g40858(csa_tree_add_51_79_groupi_n_5314 ,csa_tree_add_51_79_groupi_n_3423 ,csa_tree_add_51_79_groupi_n_4704);
  and csa_tree_add_51_79_groupi_g40859(csa_tree_add_51_79_groupi_n_5312 ,csa_tree_add_51_79_groupi_n_2943 ,csa_tree_add_51_79_groupi_n_4533);
  and csa_tree_add_51_79_groupi_g40860(csa_tree_add_51_79_groupi_n_5311 ,csa_tree_add_51_79_groupi_n_3098 ,csa_tree_add_51_79_groupi_n_4182);
  and csa_tree_add_51_79_groupi_g40861(csa_tree_add_51_79_groupi_n_5310 ,csa_tree_add_51_79_groupi_n_3146 ,csa_tree_add_51_79_groupi_n_4337);
  or csa_tree_add_51_79_groupi_g40862(csa_tree_add_51_79_groupi_n_5309 ,csa_tree_add_51_79_groupi_n_3564 ,csa_tree_add_51_79_groupi_n_4344);
  and csa_tree_add_51_79_groupi_g40863(csa_tree_add_51_79_groupi_n_5307 ,csa_tree_add_51_79_groupi_n_3149 ,csa_tree_add_51_79_groupi_n_4149);
  and csa_tree_add_51_79_groupi_g40864(csa_tree_add_51_79_groupi_n_5306 ,csa_tree_add_51_79_groupi_n_3862 ,csa_tree_add_51_79_groupi_n_4343);
  and csa_tree_add_51_79_groupi_g40865(csa_tree_add_51_79_groupi_n_5304 ,csa_tree_add_51_79_groupi_n_3522 ,csa_tree_add_51_79_groupi_n_4342);
  and csa_tree_add_51_79_groupi_g40866(csa_tree_add_51_79_groupi_n_5303 ,csa_tree_add_51_79_groupi_n_3356 ,csa_tree_add_51_79_groupi_n_4525);
  and csa_tree_add_51_79_groupi_g40867(csa_tree_add_51_79_groupi_n_5301 ,csa_tree_add_51_79_groupi_n_3338 ,csa_tree_add_51_79_groupi_n_4330);
  and csa_tree_add_51_79_groupi_g40868(csa_tree_add_51_79_groupi_n_5300 ,csa_tree_add_51_79_groupi_n_3546 ,csa_tree_add_51_79_groupi_n_4667);
  and csa_tree_add_51_79_groupi_g40869(csa_tree_add_51_79_groupi_n_5298 ,csa_tree_add_51_79_groupi_n_3158 ,csa_tree_add_51_79_groupi_n_4357);
  and csa_tree_add_51_79_groupi_g40870(csa_tree_add_51_79_groupi_n_5297 ,csa_tree_add_51_79_groupi_n_3145 ,csa_tree_add_51_79_groupi_n_4336);
  and csa_tree_add_51_79_groupi_g40871(csa_tree_add_51_79_groupi_n_5295 ,csa_tree_add_51_79_groupi_n_3090 ,csa_tree_add_51_79_groupi_n_4335);
  and csa_tree_add_51_79_groupi_g40872(csa_tree_add_51_79_groupi_n_5294 ,csa_tree_add_51_79_groupi_n_3356 ,csa_tree_add_51_79_groupi_n_4333);
  and csa_tree_add_51_79_groupi_g40873(csa_tree_add_51_79_groupi_n_5293 ,csa_tree_add_51_79_groupi_n_2932 ,csa_tree_add_51_79_groupi_n_3999);
  and csa_tree_add_51_79_groupi_g40874(csa_tree_add_51_79_groupi_n_5292 ,csa_tree_add_51_79_groupi_n_3012 ,csa_tree_add_51_79_groupi_n_4173);
  and csa_tree_add_51_79_groupi_g40875(csa_tree_add_51_79_groupi_n_5290 ,csa_tree_add_51_79_groupi_n_3006 ,csa_tree_add_51_79_groupi_n_4325);
  and csa_tree_add_51_79_groupi_g40876(csa_tree_add_51_79_groupi_n_5289 ,csa_tree_add_51_79_groupi_n_3856 ,csa_tree_add_51_79_groupi_n_4620);
  and csa_tree_add_51_79_groupi_g40877(csa_tree_add_51_79_groupi_n_5287 ,csa_tree_add_51_79_groupi_n_3092 ,csa_tree_add_51_79_groupi_n_4632);
  and csa_tree_add_51_79_groupi_g40878(csa_tree_add_51_79_groupi_n_5285 ,csa_tree_add_51_79_groupi_n_2914 ,csa_tree_add_51_79_groupi_n_3905);
  and csa_tree_add_51_79_groupi_g40879(csa_tree_add_51_79_groupi_n_5284 ,csa_tree_add_51_79_groupi_n_2960 ,csa_tree_add_51_79_groupi_n_4323);
  and csa_tree_add_51_79_groupi_g40880(csa_tree_add_51_79_groupi_n_5283 ,csa_tree_add_51_79_groupi_n_2986 ,csa_tree_add_51_79_groupi_n_4118);
  and csa_tree_add_51_79_groupi_g40881(csa_tree_add_51_79_groupi_n_5282 ,csa_tree_add_51_79_groupi_n_2972 ,csa_tree_add_51_79_groupi_n_4529);
  and csa_tree_add_51_79_groupi_g40882(csa_tree_add_51_79_groupi_n_5281 ,csa_tree_add_51_79_groupi_n_3136 ,csa_tree_add_51_79_groupi_n_4505);
  or csa_tree_add_51_79_groupi_g40883(csa_tree_add_51_79_groupi_n_5279 ,csa_tree_add_51_79_groupi_n_3857 ,csa_tree_add_51_79_groupi_n_4611);
  and csa_tree_add_51_79_groupi_g40884(csa_tree_add_51_79_groupi_n_5278 ,csa_tree_add_51_79_groupi_n_3353 ,csa_tree_add_51_79_groupi_n_4527);
  and csa_tree_add_51_79_groupi_g40885(csa_tree_add_51_79_groupi_n_5277 ,csa_tree_add_51_79_groupi_n_2991 ,csa_tree_add_51_79_groupi_n_4526);
  and csa_tree_add_51_79_groupi_g40886(csa_tree_add_51_79_groupi_n_5276 ,csa_tree_add_51_79_groupi_n_3427 ,csa_tree_add_51_79_groupi_n_4524);
  and csa_tree_add_51_79_groupi_g40887(csa_tree_add_51_79_groupi_n_5275 ,csa_tree_add_51_79_groupi_n_3106 ,csa_tree_add_51_79_groupi_n_4389);
  and csa_tree_add_51_79_groupi_g40888(csa_tree_add_51_79_groupi_n_5273 ,csa_tree_add_51_79_groupi_n_3100 ,csa_tree_add_51_79_groupi_n_4183);
  and csa_tree_add_51_79_groupi_g40889(csa_tree_add_51_79_groupi_n_5272 ,csa_tree_add_51_79_groupi_n_2976 ,csa_tree_add_51_79_groupi_n_3967);
  and csa_tree_add_51_79_groupi_g40890(csa_tree_add_51_79_groupi_n_5271 ,csa_tree_add_51_79_groupi_n_3348 ,csa_tree_add_51_79_groupi_n_4084);
  and csa_tree_add_51_79_groupi_g40891(csa_tree_add_51_79_groupi_n_5269 ,csa_tree_add_51_79_groupi_n_3449 ,csa_tree_add_51_79_groupi_n_4473);
  and csa_tree_add_51_79_groupi_g40892(csa_tree_add_51_79_groupi_n_5268 ,csa_tree_add_51_79_groupi_n_3350 ,csa_tree_add_51_79_groupi_n_4471);
  and csa_tree_add_51_79_groupi_g40893(csa_tree_add_51_79_groupi_n_5266 ,csa_tree_add_51_79_groupi_n_2969 ,csa_tree_add_51_79_groupi_n_4557);
  and csa_tree_add_51_79_groupi_g40894(csa_tree_add_51_79_groupi_n_5264 ,csa_tree_add_51_79_groupi_n_3141 ,csa_tree_add_51_79_groupi_n_4321);
  and csa_tree_add_51_79_groupi_g40895(csa_tree_add_51_79_groupi_n_5263 ,csa_tree_add_51_79_groupi_n_3411 ,csa_tree_add_51_79_groupi_n_4628);
  and csa_tree_add_51_79_groupi_g40896(csa_tree_add_51_79_groupi_n_5262 ,csa_tree_add_51_79_groupi_n_2999 ,csa_tree_add_51_79_groupi_n_4150);
  and csa_tree_add_51_79_groupi_g40897(csa_tree_add_51_79_groupi_n_5261 ,csa_tree_add_51_79_groupi_n_3523 ,csa_tree_add_51_79_groupi_n_4311);
  and csa_tree_add_51_79_groupi_g40898(csa_tree_add_51_79_groupi_n_5260 ,csa_tree_add_51_79_groupi_n_3557 ,csa_tree_add_51_79_groupi_n_4685);
  and csa_tree_add_51_79_groupi_g40899(csa_tree_add_51_79_groupi_n_5258 ,csa_tree_add_51_79_groupi_n_2957 ,csa_tree_add_51_79_groupi_n_4309);
  and csa_tree_add_51_79_groupi_g40900(csa_tree_add_51_79_groupi_n_5256 ,csa_tree_add_51_79_groupi_n_3574 ,csa_tree_add_51_79_groupi_n_4308);
  and csa_tree_add_51_79_groupi_g40901(csa_tree_add_51_79_groupi_n_5255 ,csa_tree_add_51_79_groupi_n_3525 ,csa_tree_add_51_79_groupi_n_4307);
  and csa_tree_add_51_79_groupi_g40902(csa_tree_add_51_79_groupi_n_5253 ,csa_tree_add_51_79_groupi_n_3125 ,csa_tree_add_51_79_groupi_n_4306);
  and csa_tree_add_51_79_groupi_g40903(csa_tree_add_51_79_groupi_n_5252 ,csa_tree_add_51_79_groupi_n_3848 ,csa_tree_add_51_79_groupi_n_4019);
  and csa_tree_add_51_79_groupi_g40904(csa_tree_add_51_79_groupi_n_5251 ,csa_tree_add_51_79_groupi_n_3156 ,csa_tree_add_51_79_groupi_n_4624);
  and csa_tree_add_51_79_groupi_g40905(csa_tree_add_51_79_groupi_n_5250 ,csa_tree_add_51_79_groupi_n_3339 ,csa_tree_add_51_79_groupi_n_4347);
  and csa_tree_add_51_79_groupi_g40906(csa_tree_add_51_79_groupi_n_5249 ,csa_tree_add_51_79_groupi_n_3642 ,csa_tree_add_51_79_groupi_n_4224);
  and csa_tree_add_51_79_groupi_g40907(csa_tree_add_51_79_groupi_n_5248 ,csa_tree_add_51_79_groupi_n_3421 ,csa_tree_add_51_79_groupi_n_4518);
  and csa_tree_add_51_79_groupi_g40908(csa_tree_add_51_79_groupi_n_5247 ,csa_tree_add_51_79_groupi_n_3122 ,csa_tree_add_51_79_groupi_n_4595);
  and csa_tree_add_51_79_groupi_g40909(csa_tree_add_51_79_groupi_n_5246 ,csa_tree_add_51_79_groupi_n_3034 ,csa_tree_add_51_79_groupi_n_4130);
  and csa_tree_add_51_79_groupi_g40910(csa_tree_add_51_79_groupi_n_5245 ,csa_tree_add_51_79_groupi_n_3349 ,csa_tree_add_51_79_groupi_n_4623);
  and csa_tree_add_51_79_groupi_g40911(csa_tree_add_51_79_groupi_n_5244 ,csa_tree_add_51_79_groupi_n_3420 ,csa_tree_add_51_79_groupi_n_4515);
  and csa_tree_add_51_79_groupi_g40912(csa_tree_add_51_79_groupi_n_5242 ,csa_tree_add_51_79_groupi_n_3372 ,csa_tree_add_51_79_groupi_n_4218);
  and csa_tree_add_51_79_groupi_g40913(csa_tree_add_51_79_groupi_n_5241 ,csa_tree_add_51_79_groupi_n_3584 ,csa_tree_add_51_79_groupi_n_4216);
  and csa_tree_add_51_79_groupi_g40914(csa_tree_add_51_79_groupi_n_5239 ,csa_tree_add_51_79_groupi_n_3071 ,csa_tree_add_51_79_groupi_n_4215);
  and csa_tree_add_51_79_groupi_g40915(csa_tree_add_51_79_groupi_n_5238 ,csa_tree_add_51_79_groupi_n_3120 ,csa_tree_add_51_79_groupi_n_4708);
  and csa_tree_add_51_79_groupi_g40916(csa_tree_add_51_79_groupi_n_5237 ,csa_tree_add_51_79_groupi_n_3005 ,csa_tree_add_51_79_groupi_n_4116);
  and csa_tree_add_51_79_groupi_g40917(csa_tree_add_51_79_groupi_n_5235 ,csa_tree_add_51_79_groupi_n_3050 ,csa_tree_add_51_79_groupi_n_4625);
  and csa_tree_add_51_79_groupi_g40918(csa_tree_add_51_79_groupi_n_5234 ,csa_tree_add_51_79_groupi_n_3386 ,csa_tree_add_51_79_groupi_n_4387);
  and csa_tree_add_51_79_groupi_g40919(csa_tree_add_51_79_groupi_n_5233 ,csa_tree_add_51_79_groupi_n_2891 ,csa_tree_add_51_79_groupi_n_3955);
  and csa_tree_add_51_79_groupi_g40920(csa_tree_add_51_79_groupi_n_5232 ,csa_tree_add_51_79_groupi_n_3868 ,csa_tree_add_51_79_groupi_n_4209);
  and csa_tree_add_51_79_groupi_g40921(csa_tree_add_51_79_groupi_n_5231 ,csa_tree_add_51_79_groupi_n_2894 ,csa_tree_add_51_79_groupi_n_4210);
  and csa_tree_add_51_79_groupi_g40922(csa_tree_add_51_79_groupi_n_5230 ,csa_tree_add_51_79_groupi_n_2918 ,csa_tree_add_51_79_groupi_n_4457);
  and csa_tree_add_51_79_groupi_g40923(csa_tree_add_51_79_groupi_n_5229 ,csa_tree_add_51_79_groupi_n_3344 ,csa_tree_add_51_79_groupi_n_4119);
  and csa_tree_add_51_79_groupi_g40924(csa_tree_add_51_79_groupi_n_5227 ,csa_tree_add_51_79_groupi_n_2952 ,csa_tree_add_51_79_groupi_n_4205);
  and csa_tree_add_51_79_groupi_g40925(csa_tree_add_51_79_groupi_n_5226 ,csa_tree_add_51_79_groupi_n_3037 ,csa_tree_add_51_79_groupi_n_4586);
  and csa_tree_add_51_79_groupi_g40926(csa_tree_add_51_79_groupi_n_5225 ,csa_tree_add_51_79_groupi_n_3077 ,csa_tree_add_51_79_groupi_n_4180);
  and csa_tree_add_51_79_groupi_g40927(csa_tree_add_51_79_groupi_n_5224 ,csa_tree_add_51_79_groupi_n_3126 ,csa_tree_add_51_79_groupi_n_4622);
  and csa_tree_add_51_79_groupi_g40928(csa_tree_add_51_79_groupi_n_5223 ,csa_tree_add_51_79_groupi_n_2964 ,csa_tree_add_51_79_groupi_n_4203);
  and csa_tree_add_51_79_groupi_g40929(csa_tree_add_51_79_groupi_n_5222 ,csa_tree_add_51_79_groupi_n_3099 ,csa_tree_add_51_79_groupi_n_4201);
  and csa_tree_add_51_79_groupi_g40930(csa_tree_add_51_79_groupi_n_5221 ,csa_tree_add_51_79_groupi_n_3085 ,csa_tree_add_51_79_groupi_n_4511);
  and csa_tree_add_51_79_groupi_g40931(csa_tree_add_51_79_groupi_n_5220 ,csa_tree_add_51_79_groupi_n_3542 ,csa_tree_add_51_79_groupi_n_4448);
  and csa_tree_add_51_79_groupi_g40932(csa_tree_add_51_79_groupi_n_5219 ,csa_tree_add_51_79_groupi_n_3560 ,csa_tree_add_51_79_groupi_n_4195);
  and csa_tree_add_51_79_groupi_g40933(csa_tree_add_51_79_groupi_n_5218 ,csa_tree_add_51_79_groupi_n_3114 ,csa_tree_add_51_79_groupi_n_4033);
  and csa_tree_add_51_79_groupi_g40934(csa_tree_add_51_79_groupi_n_5216 ,csa_tree_add_51_79_groupi_n_3349 ,csa_tree_add_51_79_groupi_n_4345);
  and csa_tree_add_51_79_groupi_g40935(csa_tree_add_51_79_groupi_n_5215 ,csa_tree_add_51_79_groupi_n_3117 ,csa_tree_add_51_79_groupi_n_4510);
  and csa_tree_add_51_79_groupi_g40936(csa_tree_add_51_79_groupi_n_5214 ,csa_tree_add_51_79_groupi_n_3116 ,csa_tree_add_51_79_groupi_n_4509);
  and csa_tree_add_51_79_groupi_g40937(csa_tree_add_51_79_groupi_n_5213 ,csa_tree_add_51_79_groupi_n_3442 ,csa_tree_add_51_79_groupi_n_4507);
  and csa_tree_add_51_79_groupi_g40938(csa_tree_add_51_79_groupi_n_5212 ,csa_tree_add_51_79_groupi_n_3032 ,csa_tree_add_51_79_groupi_n_4020);
  and csa_tree_add_51_79_groupi_g40939(csa_tree_add_51_79_groupi_n_5211 ,csa_tree_add_51_79_groupi_n_3450 ,csa_tree_add_51_79_groupi_n_4691);
  and csa_tree_add_51_79_groupi_g40940(csa_tree_add_51_79_groupi_n_5209 ,csa_tree_add_51_79_groupi_n_3431 ,csa_tree_add_51_79_groupi_n_4392);
  and csa_tree_add_51_79_groupi_g40941(csa_tree_add_51_79_groupi_n_5208 ,csa_tree_add_51_79_groupi_n_3413 ,csa_tree_add_51_79_groupi_n_4508);
  and csa_tree_add_51_79_groupi_g40942(csa_tree_add_51_79_groupi_n_5206 ,csa_tree_add_51_79_groupi_n_3363 ,csa_tree_add_51_79_groupi_n_4339);
  and csa_tree_add_51_79_groupi_g40943(csa_tree_add_51_79_groupi_n_5205 ,csa_tree_add_51_79_groupi_n_3390 ,csa_tree_add_51_79_groupi_n_4665);
  and csa_tree_add_51_79_groupi_g40944(csa_tree_add_51_79_groupi_n_5204 ,csa_tree_add_51_79_groupi_n_3089 ,csa_tree_add_51_79_groupi_n_4161);
  and csa_tree_add_51_79_groupi_g40945(csa_tree_add_51_79_groupi_n_5203 ,csa_tree_add_51_79_groupi_n_3454 ,csa_tree_add_51_79_groupi_n_4663);
  and csa_tree_add_51_79_groupi_g40946(csa_tree_add_51_79_groupi_n_5202 ,csa_tree_add_51_79_groupi_n_3649 ,csa_tree_add_51_79_groupi_n_4370);
  and csa_tree_add_51_79_groupi_g40947(csa_tree_add_51_79_groupi_n_5201 ,csa_tree_add_51_79_groupi_n_3509 ,csa_tree_add_51_79_groupi_n_4683);
  and csa_tree_add_51_79_groupi_g40948(csa_tree_add_51_79_groupi_n_5199 ,csa_tree_add_51_79_groupi_n_3444 ,csa_tree_add_51_79_groupi_n_4391);
  and csa_tree_add_51_79_groupi_g40949(csa_tree_add_51_79_groupi_n_5198 ,csa_tree_add_51_79_groupi_n_3535 ,csa_tree_add_51_79_groupi_n_4501);
  and csa_tree_add_51_79_groupi_g40950(csa_tree_add_51_79_groupi_n_5197 ,csa_tree_add_51_79_groupi_n_3052 ,csa_tree_add_51_79_groupi_n_4121);
  and csa_tree_add_51_79_groupi_g40951(csa_tree_add_51_79_groupi_n_5196 ,csa_tree_add_51_79_groupi_n_3519 ,csa_tree_add_51_79_groupi_n_4575);
  and csa_tree_add_51_79_groupi_g40952(csa_tree_add_51_79_groupi_n_5195 ,csa_tree_add_51_79_groupi_n_3487 ,csa_tree_add_51_79_groupi_n_4500);
  and csa_tree_add_51_79_groupi_g40953(csa_tree_add_51_79_groupi_n_5194 ,csa_tree_add_51_79_groupi_n_3075 ,csa_tree_add_51_79_groupi_n_4514);
  and csa_tree_add_51_79_groupi_g40954(csa_tree_add_51_79_groupi_n_5193 ,csa_tree_add_51_79_groupi_n_3441 ,csa_tree_add_51_79_groupi_n_4498);
  and csa_tree_add_51_79_groupi_g40955(csa_tree_add_51_79_groupi_n_5192 ,csa_tree_add_51_79_groupi_n_3385 ,csa_tree_add_51_79_groupi_n_4053);
  and csa_tree_add_51_79_groupi_g40956(csa_tree_add_51_79_groupi_n_5191 ,csa_tree_add_51_79_groupi_n_3446 ,csa_tree_add_51_79_groupi_n_4499);
  and csa_tree_add_51_79_groupi_g40957(csa_tree_add_51_79_groupi_n_5190 ,csa_tree_add_51_79_groupi_n_3513 ,csa_tree_add_51_79_groupi_n_4618);
  and csa_tree_add_51_79_groupi_g40958(csa_tree_add_51_79_groupi_n_5189 ,csa_tree_add_51_79_groupi_n_3108 ,csa_tree_add_51_79_groupi_n_4377);
  and csa_tree_add_51_79_groupi_g40959(csa_tree_add_51_79_groupi_n_5188 ,csa_tree_add_51_79_groupi_n_3410 ,csa_tree_add_51_79_groupi_n_4495);
  and csa_tree_add_51_79_groupi_g40960(csa_tree_add_51_79_groupi_n_5187 ,csa_tree_add_51_79_groupi_n_3532 ,csa_tree_add_51_79_groupi_n_4552);
  and csa_tree_add_51_79_groupi_g40961(csa_tree_add_51_79_groupi_n_5186 ,csa_tree_add_51_79_groupi_n_3152 ,csa_tree_add_51_79_groupi_n_4157);
  and csa_tree_add_51_79_groupi_g40962(csa_tree_add_51_79_groupi_n_5184 ,csa_tree_add_51_79_groupi_n_3868 ,csa_tree_add_51_79_groupi_n_4583);
  and csa_tree_add_51_79_groupi_g40963(csa_tree_add_51_79_groupi_n_5183 ,csa_tree_add_51_79_groupi_n_3405 ,csa_tree_add_51_79_groupi_n_4494);
  and csa_tree_add_51_79_groupi_g40964(csa_tree_add_51_79_groupi_n_5182 ,csa_tree_add_51_79_groupi_n_3051 ,csa_tree_add_51_79_groupi_n_4220);
  and csa_tree_add_51_79_groupi_g40965(csa_tree_add_51_79_groupi_n_5181 ,csa_tree_add_51_79_groupi_n_3345 ,csa_tree_add_51_79_groupi_n_4353);
  and csa_tree_add_51_79_groupi_g40966(csa_tree_add_51_79_groupi_n_5180 ,csa_tree_add_51_79_groupi_n_3058 ,csa_tree_add_51_79_groupi_n_4079);
  and csa_tree_add_51_79_groupi_g40967(csa_tree_add_51_79_groupi_n_5179 ,csa_tree_add_51_79_groupi_n_3863 ,csa_tree_add_51_79_groupi_n_4465);
  and csa_tree_add_51_79_groupi_g40968(csa_tree_add_51_79_groupi_n_5177 ,csa_tree_add_51_79_groupi_n_2995 ,csa_tree_add_51_79_groupi_n_4475);
  and csa_tree_add_51_79_groupi_g40969(csa_tree_add_51_79_groupi_n_5176 ,csa_tree_add_51_79_groupi_n_3438 ,csa_tree_add_51_79_groupi_n_4492);
  and csa_tree_add_51_79_groupi_g40970(csa_tree_add_51_79_groupi_n_5175 ,csa_tree_add_51_79_groupi_n_3581 ,csa_tree_add_51_79_groupi_n_4700);
  and csa_tree_add_51_79_groupi_g40971(csa_tree_add_51_79_groupi_n_5174 ,csa_tree_add_51_79_groupi_n_3388 ,csa_tree_add_51_79_groupi_n_4488);
  and csa_tree_add_51_79_groupi_g40972(csa_tree_add_51_79_groupi_n_5173 ,csa_tree_add_51_79_groupi_n_3534 ,csa_tree_add_51_79_groupi_n_4364);
  and csa_tree_add_51_79_groupi_g40973(csa_tree_add_51_79_groupi_n_5172 ,csa_tree_add_51_79_groupi_n_2966 ,csa_tree_add_51_79_groupi_n_4487);
  and csa_tree_add_51_79_groupi_g40974(csa_tree_add_51_79_groupi_n_5171 ,csa_tree_add_51_79_groupi_n_3582 ,csa_tree_add_51_79_groupi_n_4145);
  and csa_tree_add_51_79_groupi_g40975(csa_tree_add_51_79_groupi_n_5170 ,csa_tree_add_51_79_groupi_n_3400 ,csa_tree_add_51_79_groupi_n_4176);
  and csa_tree_add_51_79_groupi_g40976(csa_tree_add_51_79_groupi_n_5169 ,csa_tree_add_51_79_groupi_n_3073 ,csa_tree_add_51_79_groupi_n_4143);
  and csa_tree_add_51_79_groupi_g40977(csa_tree_add_51_79_groupi_n_5168 ,csa_tree_add_51_79_groupi_n_3002 ,csa_tree_add_51_79_groupi_n_4615);
  and csa_tree_add_51_79_groupi_g40978(csa_tree_add_51_79_groupi_n_5167 ,csa_tree_add_51_79_groupi_n_3035 ,csa_tree_add_51_79_groupi_n_4141);
  and csa_tree_add_51_79_groupi_g40979(csa_tree_add_51_79_groupi_n_5166 ,csa_tree_add_51_79_groupi_n_3510 ,csa_tree_add_51_79_groupi_n_4614);
  and csa_tree_add_51_79_groupi_g40980(csa_tree_add_51_79_groupi_n_5165 ,csa_tree_add_51_79_groupi_n_3079 ,csa_tree_add_51_79_groupi_n_4360);
  and csa_tree_add_51_79_groupi_g40981(csa_tree_add_51_79_groupi_n_5164 ,csa_tree_add_51_79_groupi_n_2978 ,csa_tree_add_51_79_groupi_n_4024);
  and csa_tree_add_51_79_groupi_g40982(csa_tree_add_51_79_groupi_n_5163 ,csa_tree_add_51_79_groupi_n_3342 ,csa_tree_add_51_79_groupi_n_4104);
  and csa_tree_add_51_79_groupi_g40983(csa_tree_add_51_79_groupi_n_5161 ,csa_tree_add_51_79_groupi_n_3010 ,csa_tree_add_51_79_groupi_n_4032);
  and csa_tree_add_51_79_groupi_g40984(csa_tree_add_51_79_groupi_n_5160 ,csa_tree_add_51_79_groupi_n_3028 ,csa_tree_add_51_79_groupi_n_4400);
  and csa_tree_add_51_79_groupi_g40985(csa_tree_add_51_79_groupi_n_5158 ,csa_tree_add_51_79_groupi_n_3030 ,csa_tree_add_51_79_groupi_n_4449);
  and csa_tree_add_51_79_groupi_g40986(csa_tree_add_51_79_groupi_n_5157 ,csa_tree_add_51_79_groupi_n_3492 ,csa_tree_add_51_79_groupi_n_4484);
  and csa_tree_add_51_79_groupi_g40987(csa_tree_add_51_79_groupi_n_5156 ,csa_tree_add_51_79_groupi_n_3495 ,csa_tree_add_51_79_groupi_n_4381);
  and csa_tree_add_51_79_groupi_g40988(csa_tree_add_51_79_groupi_n_5155 ,csa_tree_add_51_79_groupi_n_3357 ,csa_tree_add_51_79_groupi_n_4480);
  and csa_tree_add_51_79_groupi_g40989(csa_tree_add_51_79_groupi_n_5153 ,csa_tree_add_51_79_groupi_n_3851 ,csa_tree_add_51_79_groupi_n_4388);
  not csa_tree_add_51_79_groupi_g40992(csa_tree_add_51_79_groupi_n_5035 ,csa_tree_add_51_79_groupi_n_5034);
  not csa_tree_add_51_79_groupi_g40993(csa_tree_add_51_79_groupi_n_4988 ,csa_tree_add_51_79_groupi_n_4989);
  not csa_tree_add_51_79_groupi_g40994(csa_tree_add_51_79_groupi_n_4967 ,csa_tree_add_51_79_groupi_n_4968);
  not csa_tree_add_51_79_groupi_g40995(csa_tree_add_51_79_groupi_n_4963 ,csa_tree_add_51_79_groupi_n_4964);
  not csa_tree_add_51_79_groupi_g40996(csa_tree_add_51_79_groupi_n_4961 ,csa_tree_add_51_79_groupi_n_4962);
  not csa_tree_add_51_79_groupi_g40997(csa_tree_add_51_79_groupi_n_4958 ,csa_tree_add_51_79_groupi_n_4959);
  not csa_tree_add_51_79_groupi_g40998(csa_tree_add_51_79_groupi_n_4956 ,csa_tree_add_51_79_groupi_n_4957);
  not csa_tree_add_51_79_groupi_g40999(csa_tree_add_51_79_groupi_n_4945 ,csa_tree_add_51_79_groupi_n_4946);
  not csa_tree_add_51_79_groupi_g41000(csa_tree_add_51_79_groupi_n_4931 ,csa_tree_add_51_79_groupi_n_4932);
  not csa_tree_add_51_79_groupi_g41001(csa_tree_add_51_79_groupi_n_4923 ,csa_tree_add_51_79_groupi_n_4922);
  not csa_tree_add_51_79_groupi_g41002(csa_tree_add_51_79_groupi_n_4896 ,csa_tree_add_51_79_groupi_n_4897);
  not csa_tree_add_51_79_groupi_g41003(csa_tree_add_51_79_groupi_n_4891 ,csa_tree_add_51_79_groupi_n_4892);
  not csa_tree_add_51_79_groupi_g41004(csa_tree_add_51_79_groupi_n_4874 ,csa_tree_add_51_79_groupi_n_4873);
  not csa_tree_add_51_79_groupi_g41005(csa_tree_add_51_79_groupi_n_4869 ,csa_tree_add_51_79_groupi_n_4870);
  not csa_tree_add_51_79_groupi_g41006(csa_tree_add_51_79_groupi_n_4865 ,csa_tree_add_51_79_groupi_n_4866);
  not csa_tree_add_51_79_groupi_g41007(csa_tree_add_51_79_groupi_n_4863 ,csa_tree_add_51_79_groupi_n_4862);
  not csa_tree_add_51_79_groupi_g41008(csa_tree_add_51_79_groupi_n_4858 ,csa_tree_add_51_79_groupi_n_4857);
  not csa_tree_add_51_79_groupi_g41009(csa_tree_add_51_79_groupi_n_4855 ,csa_tree_add_51_79_groupi_n_4856);
  not csa_tree_add_51_79_groupi_g41010(csa_tree_add_51_79_groupi_n_4839 ,csa_tree_add_51_79_groupi_n_4840);
  not csa_tree_add_51_79_groupi_g41011(csa_tree_add_51_79_groupi_n_4834 ,csa_tree_add_51_79_groupi_n_4833);
  not csa_tree_add_51_79_groupi_g41012(csa_tree_add_51_79_groupi_n_4827 ,csa_tree_add_51_79_groupi_n_4828);
  not csa_tree_add_51_79_groupi_g41013(csa_tree_add_51_79_groupi_n_4825 ,csa_tree_add_51_79_groupi_n_4826);
  not csa_tree_add_51_79_groupi_g41014(csa_tree_add_51_79_groupi_n_4823 ,csa_tree_add_51_79_groupi_n_4824);
  not csa_tree_add_51_79_groupi_g41015(csa_tree_add_51_79_groupi_n_4811 ,csa_tree_add_51_79_groupi_n_11);
  not csa_tree_add_51_79_groupi_g41016(csa_tree_add_51_79_groupi_n_4804 ,csa_tree_add_51_79_groupi_n_4803);
  not csa_tree_add_51_79_groupi_g41017(csa_tree_add_51_79_groupi_n_4795 ,csa_tree_add_51_79_groupi_n_4796);
  nor csa_tree_add_51_79_groupi_g41018(csa_tree_add_51_79_groupi_n_4792 ,csa_tree_add_51_79_groupi_n_4281 ,csa_tree_add_51_79_groupi_n_4278);
  or csa_tree_add_51_79_groupi_g41019(csa_tree_add_51_79_groupi_n_4791 ,csa_tree_add_51_79_groupi_n_3322 ,csa_tree_add_51_79_groupi_n_4707);
  and csa_tree_add_51_79_groupi_g41020(csa_tree_add_51_79_groupi_n_4790 ,csa_tree_add_51_79_groupi_n_2555 ,csa_tree_add_51_79_groupi_n_4229);
  and csa_tree_add_51_79_groupi_g41021(csa_tree_add_51_79_groupi_n_4789 ,csa_tree_add_51_79_groupi_n_4226 ,csa_tree_add_51_79_groupi_n_4225);
  or csa_tree_add_51_79_groupi_g41022(csa_tree_add_51_79_groupi_n_4788 ,csa_tree_add_51_79_groupi_n_3333 ,csa_tree_add_51_79_groupi_n_4644);
  nor csa_tree_add_51_79_groupi_g41023(csa_tree_add_51_79_groupi_n_4787 ,csa_tree_add_51_79_groupi_n_4255 ,csa_tree_add_51_79_groupi_n_4282);
  nor csa_tree_add_51_79_groupi_g41024(csa_tree_add_51_79_groupi_n_4786 ,csa_tree_add_51_79_groupi_n_4238 ,csa_tree_add_51_79_groupi_n_4232);
  or csa_tree_add_51_79_groupi_g41025(csa_tree_add_51_79_groupi_n_4785 ,csa_tree_add_51_79_groupi_n_4241 ,csa_tree_add_51_79_groupi_n_4262);
  or csa_tree_add_51_79_groupi_g41026(csa_tree_add_51_79_groupi_n_4784 ,csa_tree_add_51_79_groupi_n_4246 ,csa_tree_add_51_79_groupi_n_4257);
  or csa_tree_add_51_79_groupi_g41027(csa_tree_add_51_79_groupi_n_4783 ,csa_tree_add_51_79_groupi_n_4280 ,csa_tree_add_51_79_groupi_n_4279);
  nor csa_tree_add_51_79_groupi_g41028(csa_tree_add_51_79_groupi_n_4782 ,csa_tree_add_51_79_groupi_n_4259 ,csa_tree_add_51_79_groupi_n_4239);
  nor csa_tree_add_51_79_groupi_g41029(csa_tree_add_51_79_groupi_n_4781 ,csa_tree_add_51_79_groupi_n_4245 ,csa_tree_add_51_79_groupi_n_4252);
  nor csa_tree_add_51_79_groupi_g41030(csa_tree_add_51_79_groupi_n_4780 ,csa_tree_add_51_79_groupi_n_4277 ,csa_tree_add_51_79_groupi_n_4272);
  nor csa_tree_add_51_79_groupi_g41031(csa_tree_add_51_79_groupi_n_4779 ,csa_tree_add_51_79_groupi_n_4242 ,csa_tree_add_51_79_groupi_n_4261);
  or csa_tree_add_51_79_groupi_g41032(csa_tree_add_51_79_groupi_n_4778 ,csa_tree_add_51_79_groupi_n_4254 ,csa_tree_add_51_79_groupi_n_4283);
  nor csa_tree_add_51_79_groupi_g41033(csa_tree_add_51_79_groupi_n_4777 ,csa_tree_add_51_79_groupi_n_4269 ,csa_tree_add_51_79_groupi_n_4270);
  or csa_tree_add_51_79_groupi_g41034(csa_tree_add_51_79_groupi_n_4776 ,csa_tree_add_51_79_groupi_n_4268 ,csa_tree_add_51_79_groupi_n_4271);
  or csa_tree_add_51_79_groupi_g41035(csa_tree_add_51_79_groupi_n_4775 ,csa_tree_add_51_79_groupi_n_4244 ,csa_tree_add_51_79_groupi_n_4253);
  or csa_tree_add_51_79_groupi_g41036(csa_tree_add_51_79_groupi_n_4774 ,csa_tree_add_51_79_groupi_n_4258 ,csa_tree_add_51_79_groupi_n_4240);
  or csa_tree_add_51_79_groupi_g41037(csa_tree_add_51_79_groupi_n_4773 ,csa_tree_add_51_79_groupi_n_4276 ,csa_tree_add_51_79_groupi_n_4273);
  nor csa_tree_add_51_79_groupi_g41038(csa_tree_add_51_79_groupi_n_4772 ,csa_tree_add_51_79_groupi_n_4247 ,csa_tree_add_51_79_groupi_n_4256);
  or csa_tree_add_51_79_groupi_g41039(csa_tree_add_51_79_groupi_n_4771 ,csa_tree_add_51_79_groupi_n_3312 ,csa_tree_add_51_79_groupi_n_4047);
  or csa_tree_add_51_79_groupi_g41040(csa_tree_add_51_79_groupi_n_4770 ,csa_tree_add_51_79_groupi_n_4227 ,csa_tree_add_51_79_groupi_n_4275);
  nor csa_tree_add_51_79_groupi_g41041(csa_tree_add_51_79_groupi_n_4769 ,csa_tree_add_51_79_groupi_n_4251 ,csa_tree_add_51_79_groupi_n_4248);
  or csa_tree_add_51_79_groupi_g41042(csa_tree_add_51_79_groupi_n_4768 ,csa_tree_add_51_79_groupi_n_4250 ,csa_tree_add_51_79_groupi_n_4249);
  nor csa_tree_add_51_79_groupi_g41043(csa_tree_add_51_79_groupi_n_4767 ,csa_tree_add_51_79_groupi_n_4266 ,csa_tree_add_51_79_groupi_n_4263);
  or csa_tree_add_51_79_groupi_g41044(csa_tree_add_51_79_groupi_n_4766 ,csa_tree_add_51_79_groupi_n_4265 ,csa_tree_add_51_79_groupi_n_4264);
  nor csa_tree_add_51_79_groupi_g41045(csa_tree_add_51_79_groupi_n_4765 ,csa_tree_add_51_79_groupi_n_4228 ,csa_tree_add_51_79_groupi_n_4274);
  or csa_tree_add_51_79_groupi_g41046(csa_tree_add_51_79_groupi_n_4764 ,csa_tree_add_51_79_groupi_n_4237 ,csa_tree_add_51_79_groupi_n_4233);
  or csa_tree_add_51_79_groupi_g41047(csa_tree_add_51_79_groupi_n_4763 ,csa_tree_add_51_79_groupi_n_4234 ,csa_tree_add_51_79_groupi_n_4235);
  and csa_tree_add_51_79_groupi_g41048(csa_tree_add_51_79_groupi_n_4762 ,csa_tree_add_51_79_groupi_n_4236 ,csa_tree_add_51_79_groupi_n_4267);
  and csa_tree_add_51_79_groupi_g41049(csa_tree_add_51_79_groupi_n_4761 ,csa_tree_add_51_79_groupi_n_4243 ,csa_tree_add_51_79_groupi_n_4230);
  or csa_tree_add_51_79_groupi_g41050(csa_tree_add_51_79_groupi_n_4760 ,csa_tree_add_51_79_groupi_n_4243 ,csa_tree_add_51_79_groupi_n_4230);
  or csa_tree_add_51_79_groupi_g41051(csa_tree_add_51_79_groupi_n_4759 ,csa_tree_add_51_79_groupi_n_4236 ,csa_tree_add_51_79_groupi_n_4267);
  and csa_tree_add_51_79_groupi_g41052(csa_tree_add_51_79_groupi_n_4758 ,csa_tree_add_51_79_groupi_n_3334 ,csa_tree_add_51_79_groupi_n_4549);
  and csa_tree_add_51_79_groupi_g41053(csa_tree_add_51_79_groupi_n_4757 ,csa_tree_add_51_79_groupi_n_4234 ,csa_tree_add_51_79_groupi_n_4235);
  or csa_tree_add_51_79_groupi_g41054(csa_tree_add_51_79_groupi_n_4756 ,csa_tree_add_51_79_groupi_n_4260 ,csa_tree_add_51_79_groupi_n_4231);
  and csa_tree_add_51_79_groupi_g41055(csa_tree_add_51_79_groupi_n_4755 ,csa_tree_add_51_79_groupi_n_4260 ,csa_tree_add_51_79_groupi_n_4231);
  or csa_tree_add_51_79_groupi_g41056(csa_tree_add_51_79_groupi_n_4754 ,csa_tree_add_51_79_groupi_n_3328 ,csa_tree_add_51_79_groupi_n_3948);
  or csa_tree_add_51_79_groupi_g41057(csa_tree_add_51_79_groupi_n_4753 ,csa_tree_add_51_79_groupi_n_3324 ,csa_tree_add_51_79_groupi_n_3945);
  or csa_tree_add_51_79_groupi_g41058(csa_tree_add_51_79_groupi_n_4752 ,csa_tree_add_51_79_groupi_n_3326 ,csa_tree_add_51_79_groupi_n_3944);
  and csa_tree_add_51_79_groupi_g41059(csa_tree_add_51_79_groupi_n_4751 ,csa_tree_add_51_79_groupi_n_3327 ,csa_tree_add_51_79_groupi_n_3882);
  and csa_tree_add_51_79_groupi_g41060(csa_tree_add_51_79_groupi_n_4750 ,csa_tree_add_51_79_groupi_n_3330 ,csa_tree_add_51_79_groupi_n_3928);
  xnor csa_tree_add_51_79_groupi_g41061(csa_tree_add_51_79_groupi_n_4749 ,csa_tree_add_51_79_groupi_n_3236 ,csa_tree_add_51_79_groupi_n_3288);
  xnor csa_tree_add_51_79_groupi_g41062(csa_tree_add_51_79_groupi_n_4748 ,csa_tree_add_51_79_groupi_n_3801 ,csa_tree_add_51_79_groupi_n_3800);
  xnor csa_tree_add_51_79_groupi_g41063(csa_tree_add_51_79_groupi_n_4747 ,csa_tree_add_51_79_groupi_n_3242 ,csa_tree_add_51_79_groupi_n_3738);
  xnor csa_tree_add_51_79_groupi_g41064(csa_tree_add_51_79_groupi_n_4746 ,csa_tree_add_51_79_groupi_n_3263 ,csa_tree_add_51_79_groupi_n_3266);
  xnor csa_tree_add_51_79_groupi_g41065(csa_tree_add_51_79_groupi_n_4745 ,csa_tree_add_51_79_groupi_n_3763 ,csa_tree_add_51_79_groupi_n_3245);
  xnor csa_tree_add_51_79_groupi_g41066(csa_tree_add_51_79_groupi_n_4744 ,csa_tree_add_51_79_groupi_n_3815 ,csa_tree_add_51_79_groupi_n_3797);
  xnor csa_tree_add_51_79_groupi_g41067(csa_tree_add_51_79_groupi_n_4743 ,csa_tree_add_51_79_groupi_n_3244 ,csa_tree_add_51_79_groupi_n_3796);
  xnor csa_tree_add_51_79_groupi_g41068(csa_tree_add_51_79_groupi_n_4742 ,csa_tree_add_51_79_groupi_n_3216 ,csa_tree_add_51_79_groupi_n_3795);
  xnor csa_tree_add_51_79_groupi_g41069(csa_tree_add_51_79_groupi_n_4741 ,csa_tree_add_51_79_groupi_n_3252 ,csa_tree_add_51_79_groupi_n_3276);
  xnor csa_tree_add_51_79_groupi_g41070(csa_tree_add_51_79_groupi_n_4740 ,csa_tree_add_51_79_groupi_n_3297 ,csa_tree_add_51_79_groupi_n_3753);
  xnor csa_tree_add_51_79_groupi_g41071(csa_tree_add_51_79_groupi_n_4739 ,csa_tree_add_51_79_groupi_n_3243 ,csa_tree_add_51_79_groupi_n_3737);
  xnor csa_tree_add_51_79_groupi_g41072(csa_tree_add_51_79_groupi_n_4738 ,csa_tree_add_51_79_groupi_n_3249 ,csa_tree_add_51_79_groupi_n_3755);
  xnor csa_tree_add_51_79_groupi_g41073(csa_tree_add_51_79_groupi_n_4737 ,csa_tree_add_51_79_groupi_n_3293 ,csa_tree_add_51_79_groupi_n_3209);
  xnor csa_tree_add_51_79_groupi_g41074(csa_tree_add_51_79_groupi_n_4736 ,csa_tree_add_51_79_groupi_n_3199 ,csa_tree_add_51_79_groupi_n_3311);
  xnor csa_tree_add_51_79_groupi_g41075(csa_tree_add_51_79_groupi_n_4735 ,csa_tree_add_51_79_groupi_n_3207 ,csa_tree_add_51_79_groupi_n_3224);
  xnor csa_tree_add_51_79_groupi_g41076(csa_tree_add_51_79_groupi_n_4734 ,csa_tree_add_51_79_groupi_n_3198 ,csa_tree_add_51_79_groupi_n_3201);
  xnor csa_tree_add_51_79_groupi_g41077(csa_tree_add_51_79_groupi_n_4733 ,csa_tree_add_51_79_groupi_n_3230 ,csa_tree_add_51_79_groupi_n_3325);
  xnor csa_tree_add_51_79_groupi_g41078(csa_tree_add_51_79_groupi_n_4732 ,csa_tree_add_51_79_groupi_n_3277 ,csa_tree_add_51_79_groupi_n_3319);
  xnor csa_tree_add_51_79_groupi_g41079(csa_tree_add_51_79_groupi_n_4731 ,csa_tree_add_51_79_groupi_n_3781 ,csa_tree_add_51_79_groupi_n_3790);
  xnor csa_tree_add_51_79_groupi_g41080(csa_tree_add_51_79_groupi_n_4730 ,csa_tree_add_51_79_groupi_n_3257 ,csa_tree_add_51_79_groupi_n_3294);
  xnor csa_tree_add_51_79_groupi_g41081(csa_tree_add_51_79_groupi_n_4729 ,csa_tree_add_51_79_groupi_n_3195 ,csa_tree_add_51_79_groupi_n_3333);
  xnor csa_tree_add_51_79_groupi_g41082(csa_tree_add_51_79_groupi_n_4728 ,csa_tree_add_51_79_groupi_n_3219 ,csa_tree_add_51_79_groupi_n_3223);
  xnor csa_tree_add_51_79_groupi_g41083(csa_tree_add_51_79_groupi_n_4727 ,csa_tree_add_51_79_groupi_n_3218 ,csa_tree_add_51_79_groupi_n_3315);
  xnor csa_tree_add_51_79_groupi_g41084(csa_tree_add_51_79_groupi_n_4726 ,csa_tree_add_51_79_groupi_n_3208 ,csa_tree_add_51_79_groupi_n_3200);
  xnor csa_tree_add_51_79_groupi_g41085(csa_tree_add_51_79_groupi_n_4725 ,csa_tree_add_51_79_groupi_n_3265 ,csa_tree_add_51_79_groupi_n_3287);
  xnor csa_tree_add_51_79_groupi_g41086(csa_tree_add_51_79_groupi_n_4724 ,csa_tree_add_51_79_groupi_n_3289 ,csa_tree_add_51_79_groupi_n_3202);
  xnor csa_tree_add_51_79_groupi_g41087(csa_tree_add_51_79_groupi_n_4723 ,csa_tree_add_51_79_groupi_n_3222 ,csa_tree_add_51_79_groupi_n_3211);
  xnor csa_tree_add_51_79_groupi_g41088(csa_tree_add_51_79_groupi_n_4722 ,csa_tree_add_51_79_groupi_n_3262 ,csa_tree_add_51_79_groupi_n_3203);
  xnor csa_tree_add_51_79_groupi_g41089(csa_tree_add_51_79_groupi_n_4721 ,csa_tree_add_51_79_groupi_n_3267 ,csa_tree_add_51_79_groupi_n_3221);
  xnor csa_tree_add_51_79_groupi_g41090(csa_tree_add_51_79_groupi_n_4720 ,csa_tree_add_51_79_groupi_n_3258 ,csa_tree_add_51_79_groupi_n_3322);
  xnor csa_tree_add_51_79_groupi_g41091(csa_tree_add_51_79_groupi_n_4719 ,csa_tree_add_51_79_groupi_n_3253 ,csa_tree_add_51_79_groupi_n_3326);
  xnor csa_tree_add_51_79_groupi_g41092(csa_tree_add_51_79_groupi_n_4718 ,csa_tree_add_51_79_groupi_n_3823 ,csa_tree_add_51_79_groupi_n_3255);
  xnor csa_tree_add_51_79_groupi_g41093(csa_tree_add_51_79_groupi_n_4717 ,csa_tree_add_51_79_groupi_n_3307 ,csa_tree_add_51_79_groupi_n_3274);
  xnor csa_tree_add_51_79_groupi_g41094(csa_tree_add_51_79_groupi_n_4716 ,csa_tree_add_51_79_groupi_n_3206 ,csa_tree_add_51_79_groupi_n_3194);
  xnor csa_tree_add_51_79_groupi_g41096(csa_tree_add_51_79_groupi_n_4715 ,csa_tree_add_51_79_groupi_n_3210 ,csa_tree_add_51_79_groupi_n_3804);
  xnor csa_tree_add_51_79_groupi_g41097(csa_tree_add_51_79_groupi_n_4714 ,csa_tree_add_51_79_groupi_n_3787 ,csa_tree_add_51_79_groupi_n_3739);
  and csa_tree_add_51_79_groupi_g41098(csa_tree_add_51_79_groupi_n_5125 ,csa_tree_add_51_79_groupi_n_3504 ,csa_tree_add_51_79_groupi_n_4007);
  and csa_tree_add_51_79_groupi_g41099(csa_tree_add_51_79_groupi_n_5124 ,csa_tree_add_51_79_groupi_n_3497 ,csa_tree_add_51_79_groupi_n_4006);
  and csa_tree_add_51_79_groupi_g41100(csa_tree_add_51_79_groupi_n_5123 ,csa_tree_add_51_79_groupi_n_3491 ,csa_tree_add_51_79_groupi_n_4074);
  and csa_tree_add_51_79_groupi_g41101(csa_tree_add_51_79_groupi_n_5122 ,csa_tree_add_51_79_groupi_n_3384 ,csa_tree_add_51_79_groupi_n_4093);
  and csa_tree_add_51_79_groupi_g41102(csa_tree_add_51_79_groupi_n_5121 ,csa_tree_add_51_79_groupi_n_2992 ,csa_tree_add_51_79_groupi_n_4061);
  and csa_tree_add_51_79_groupi_g41103(csa_tree_add_51_79_groupi_n_5120 ,csa_tree_add_51_79_groupi_n_3448 ,csa_tree_add_51_79_groupi_n_3911);
  and csa_tree_add_51_79_groupi_g41104(csa_tree_add_51_79_groupi_n_5119 ,csa_tree_add_51_79_groupi_n_3464 ,csa_tree_add_51_79_groupi_n_4068);
  and csa_tree_add_51_79_groupi_g41105(csa_tree_add_51_79_groupi_n_5118 ,csa_tree_add_51_79_groupi_n_2931 ,csa_tree_add_51_79_groupi_n_3996);
  and csa_tree_add_51_79_groupi_g41106(csa_tree_add_51_79_groupi_n_5117 ,csa_tree_add_51_79_groupi_n_3144 ,csa_tree_add_51_79_groupi_n_4686);
  and csa_tree_add_51_79_groupi_g41107(csa_tree_add_51_79_groupi_n_5116 ,csa_tree_add_51_79_groupi_n_3017 ,csa_tree_add_51_79_groupi_n_4125);
  and csa_tree_add_51_79_groupi_g41108(csa_tree_add_51_79_groupi_n_5115 ,csa_tree_add_51_79_groupi_n_3500 ,csa_tree_add_51_79_groupi_n_4517);
  and csa_tree_add_51_79_groupi_g41109(csa_tree_add_51_79_groupi_n_5114 ,csa_tree_add_51_79_groupi_n_2913 ,csa_tree_add_51_79_groupi_n_3992);
  and csa_tree_add_51_79_groupi_g41110(csa_tree_add_51_79_groupi_n_5113 ,csa_tree_add_51_79_groupi_n_3549 ,csa_tree_add_51_79_groupi_n_4063);
  and csa_tree_add_51_79_groupi_g41111(csa_tree_add_51_79_groupi_n_5112 ,csa_tree_add_51_79_groupi_n_3863 ,csa_tree_add_51_79_groupi_n_4055);
  and csa_tree_add_51_79_groupi_g41112(csa_tree_add_51_79_groupi_n_5111 ,csa_tree_add_51_79_groupi_n_2993 ,csa_tree_add_51_79_groupi_n_4607);
  and csa_tree_add_51_79_groupi_g41113(csa_tree_add_51_79_groupi_n_5110 ,csa_tree_add_51_79_groupi_n_3418 ,csa_tree_add_51_79_groupi_n_3984);
  and csa_tree_add_51_79_groupi_g41114(csa_tree_add_51_79_groupi_n_5109 ,csa_tree_add_51_79_groupi_n_3842 ,csa_tree_add_51_79_groupi_n_4021);
  and csa_tree_add_51_79_groupi_g41115(csa_tree_add_51_79_groupi_n_5108 ,csa_tree_add_51_79_groupi_n_3397 ,csa_tree_add_51_79_groupi_n_4082);
  or csa_tree_add_51_79_groupi_g41116(csa_tree_add_51_79_groupi_n_5107 ,csa_tree_add_51_79_groupi_n_3354 ,csa_tree_add_51_79_groupi_n_4003);
  and csa_tree_add_51_79_groupi_g41117(csa_tree_add_51_79_groupi_n_5106 ,csa_tree_add_51_79_groupi_n_3425 ,csa_tree_add_51_79_groupi_n_4095);
  and csa_tree_add_51_79_groupi_g41118(csa_tree_add_51_79_groupi_n_5105 ,csa_tree_add_51_79_groupi_n_3000 ,csa_tree_add_51_79_groupi_n_4120);
  and csa_tree_add_51_79_groupi_g41119(csa_tree_add_51_79_groupi_n_5104 ,csa_tree_add_51_79_groupi_n_3127 ,csa_tree_add_51_79_groupi_n_3979);
  and csa_tree_add_51_79_groupi_g41120(csa_tree_add_51_79_groupi_n_5103 ,csa_tree_add_51_79_groupi_n_3864 ,csa_tree_add_51_79_groupi_n_4222);
  and csa_tree_add_51_79_groupi_g41121(csa_tree_add_51_79_groupi_n_5102 ,csa_tree_add_51_79_groupi_n_3024 ,csa_tree_add_51_79_groupi_n_4207);
  and csa_tree_add_51_79_groupi_g41122(csa_tree_add_51_79_groupi_n_5101 ,csa_tree_add_51_79_groupi_n_2942 ,csa_tree_add_51_79_groupi_n_4078);
  and csa_tree_add_51_79_groupi_g41123(csa_tree_add_51_79_groupi_n_5100 ,csa_tree_add_51_79_groupi_n_3060 ,csa_tree_add_51_79_groupi_n_4460);
  and csa_tree_add_51_79_groupi_g41124(csa_tree_add_51_79_groupi_n_5099 ,csa_tree_add_51_79_groupi_n_3531 ,csa_tree_add_51_79_groupi_n_3971);
  and csa_tree_add_51_79_groupi_g41125(csa_tree_add_51_79_groupi_n_5098 ,csa_tree_add_51_79_groupi_n_3428 ,csa_tree_add_51_79_groupi_n_4109);
  or csa_tree_add_51_79_groupi_g41126(csa_tree_add_51_79_groupi_n_5097 ,csa_tree_add_51_79_groupi_n_3854 ,csa_tree_add_51_79_groupi_n_4440);
  and csa_tree_add_51_79_groupi_g41128(csa_tree_add_51_79_groupi_n_5096 ,csa_tree_add_51_79_groupi_n_2977 ,csa_tree_add_51_79_groupi_n_4026);
  and csa_tree_add_51_79_groupi_g41129(csa_tree_add_51_79_groupi_n_5095 ,csa_tree_add_51_79_groupi_n_3380 ,csa_tree_add_51_79_groupi_n_3966);
  and csa_tree_add_51_79_groupi_g41130(csa_tree_add_51_79_groupi_n_5094 ,csa_tree_add_51_79_groupi_n_2912 ,csa_tree_add_51_79_groupi_n_3965);
  and csa_tree_add_51_79_groupi_g41131(csa_tree_add_51_79_groupi_n_5093 ,csa_tree_add_51_79_groupi_n_2929 ,csa_tree_add_51_79_groupi_n_4110);
  and csa_tree_add_51_79_groupi_g41132(csa_tree_add_51_79_groupi_n_5092 ,csa_tree_add_51_79_groupi_n_2970 ,csa_tree_add_51_79_groupi_n_4144);
  and csa_tree_add_51_79_groupi_g41133(csa_tree_add_51_79_groupi_n_5091 ,csa_tree_add_51_79_groupi_n_3865 ,csa_tree_add_51_79_groupi_n_4101);
  and csa_tree_add_51_79_groupi_g41134(csa_tree_add_51_79_groupi_n_5090 ,csa_tree_add_51_79_groupi_n_2910 ,csa_tree_add_51_79_groupi_n_3960);
  and csa_tree_add_51_79_groupi_g41135(csa_tree_add_51_79_groupi_n_5089 ,csa_tree_add_51_79_groupi_n_2944 ,csa_tree_add_51_79_groupi_n_4014);
  and csa_tree_add_51_79_groupi_g41136(csa_tree_add_51_79_groupi_n_5088 ,csa_tree_add_51_79_groupi_n_3590 ,csa_tree_add_51_79_groupi_n_3921);
  and csa_tree_add_51_79_groupi_g41137(csa_tree_add_51_79_groupi_n_5087 ,csa_tree_add_51_79_groupi_n_3595 ,csa_tree_add_51_79_groupi_n_3951);
  or csa_tree_add_51_79_groupi_g41138(csa_tree_add_51_79_groupi_n_5086 ,csa_tree_add_51_79_groupi_n_3370 ,csa_tree_add_51_79_groupi_n_3931);
  and csa_tree_add_51_79_groupi_g41139(csa_tree_add_51_79_groupi_n_5085 ,csa_tree_add_51_79_groupi_n_3488 ,csa_tree_add_51_79_groupi_n_3953);
  and csa_tree_add_51_79_groupi_g41140(csa_tree_add_51_79_groupi_n_5084 ,csa_tree_add_51_79_groupi_n_3568 ,csa_tree_add_51_79_groupi_n_3956);
  and csa_tree_add_51_79_groupi_g41141(csa_tree_add_51_79_groupi_n_5083 ,csa_tree_add_51_79_groupi_n_3648 ,csa_tree_add_51_79_groupi_n_3976);
  and csa_tree_add_51_79_groupi_g41142(csa_tree_add_51_79_groupi_n_5082 ,csa_tree_add_51_79_groupi_n_3596 ,csa_tree_add_51_79_groupi_n_4012);
  and csa_tree_add_51_79_groupi_g41143(csa_tree_add_51_79_groupi_n_5081 ,csa_tree_add_51_79_groupi_n_3599 ,csa_tree_add_51_79_groupi_n_4000);
  and csa_tree_add_51_79_groupi_g41144(csa_tree_add_51_79_groupi_n_5080 ,csa_tree_add_51_79_groupi_n_3506 ,csa_tree_add_51_79_groupi_n_3950);
  and csa_tree_add_51_79_groupi_g41145(csa_tree_add_51_79_groupi_n_5079 ,csa_tree_add_51_79_groupi_n_3836 ,csa_tree_add_51_79_groupi_n_4543);
  and csa_tree_add_51_79_groupi_g41146(csa_tree_add_51_79_groupi_n_5078 ,csa_tree_add_51_79_groupi_n_3453 ,csa_tree_add_51_79_groupi_n_4368);
  and csa_tree_add_51_79_groupi_g41147(csa_tree_add_51_79_groupi_n_5077 ,csa_tree_add_51_79_groupi_n_3068 ,csa_tree_add_51_79_groupi_n_4044);
  and csa_tree_add_51_79_groupi_g41148(csa_tree_add_51_79_groupi_n_5076 ,csa_tree_add_51_79_groupi_n_2987 ,csa_tree_add_51_79_groupi_n_3883);
  and csa_tree_add_51_79_groupi_g41149(csa_tree_add_51_79_groupi_n_5075 ,csa_tree_add_51_79_groupi_n_3093 ,csa_tree_add_51_79_groupi_n_4179);
  and csa_tree_add_51_79_groupi_g41150(csa_tree_add_51_79_groupi_n_5074 ,csa_tree_add_51_79_groupi_n_3065 ,csa_tree_add_51_79_groupi_n_3943);
  and csa_tree_add_51_79_groupi_g41151(csa_tree_add_51_79_groupi_n_5073 ,csa_tree_add_51_79_groupi_n_3603 ,csa_tree_add_51_79_groupi_n_4036);
  and csa_tree_add_51_79_groupi_g41152(csa_tree_add_51_79_groupi_n_5072 ,csa_tree_add_51_79_groupi_n_3606 ,csa_tree_add_51_79_groupi_n_4652);
  and csa_tree_add_51_79_groupi_g41153(csa_tree_add_51_79_groupi_n_5071 ,csa_tree_add_51_79_groupi_n_3844 ,csa_tree_add_51_79_groupi_n_4702);
  and csa_tree_add_51_79_groupi_g41154(csa_tree_add_51_79_groupi_n_5070 ,csa_tree_add_51_79_groupi_n_3608 ,csa_tree_add_51_79_groupi_n_4538);
  and csa_tree_add_51_79_groupi_g41155(csa_tree_add_51_79_groupi_n_5069 ,csa_tree_add_51_79_groupi_n_3645 ,csa_tree_add_51_79_groupi_n_4134);
  and csa_tree_add_51_79_groupi_g41156(csa_tree_add_51_79_groupi_n_5068 ,csa_tree_add_51_79_groupi_n_3682 ,csa_tree_add_51_79_groupi_n_4067);
  and csa_tree_add_51_79_groupi_g41157(csa_tree_add_51_79_groupi_n_5067 ,csa_tree_add_51_79_groupi_n_3680 ,csa_tree_add_51_79_groupi_n_4070);
  and csa_tree_add_51_79_groupi_g41158(csa_tree_add_51_79_groupi_n_5066 ,csa_tree_add_51_79_groupi_n_2937 ,csa_tree_add_51_79_groupi_n_3936);
  and csa_tree_add_51_79_groupi_g41159(csa_tree_add_51_79_groupi_n_5065 ,csa_tree_add_51_79_groupi_n_3447 ,csa_tree_add_51_79_groupi_n_4404);
  and csa_tree_add_51_79_groupi_g41160(csa_tree_add_51_79_groupi_n_5064 ,csa_tree_add_51_79_groupi_n_3623 ,csa_tree_add_51_79_groupi_n_4073);
  and csa_tree_add_51_79_groupi_g41161(csa_tree_add_51_79_groupi_n_5063 ,csa_tree_add_51_79_groupi_n_3834 ,csa_tree_add_51_79_groupi_n_4089);
  and csa_tree_add_51_79_groupi_g41162(csa_tree_add_51_79_groupi_n_5062 ,csa_tree_add_51_79_groupi_n_3440 ,csa_tree_add_51_79_groupi_n_4437);
  and csa_tree_add_51_79_groupi_g41163(csa_tree_add_51_79_groupi_n_5061 ,csa_tree_add_51_79_groupi_n_3123 ,csa_tree_add_51_79_groupi_n_3932);
  and csa_tree_add_51_79_groupi_g41164(csa_tree_add_51_79_groupi_n_5060 ,csa_tree_add_51_79_groupi_n_3650 ,csa_tree_add_51_79_groupi_n_4098);
  and csa_tree_add_51_79_groupi_g41165(csa_tree_add_51_79_groupi_n_5059 ,csa_tree_add_51_79_groupi_n_2892 ,csa_tree_add_51_79_groupi_n_3925);
  or csa_tree_add_51_79_groupi_g41166(csa_tree_add_51_79_groupi_n_5058 ,csa_tree_add_51_79_groupi_n_3335 ,csa_tree_add_51_79_groupi_n_3922);
  and csa_tree_add_51_79_groupi_g41167(csa_tree_add_51_79_groupi_n_5057 ,csa_tree_add_51_79_groupi_n_2920 ,csa_tree_add_51_79_groupi_n_3926);
  and csa_tree_add_51_79_groupi_g41168(csa_tree_add_51_79_groupi_n_5056 ,csa_tree_add_51_79_groupi_n_3646 ,csa_tree_add_51_79_groupi_n_4442);
  and csa_tree_add_51_79_groupi_g41169(csa_tree_add_51_79_groupi_n_5055 ,csa_tree_add_51_79_groupi_n_3839 ,csa_tree_add_51_79_groupi_n_4417);
  and csa_tree_add_51_79_groupi_g41170(csa_tree_add_51_79_groupi_n_5054 ,csa_tree_add_51_79_groupi_n_3699 ,csa_tree_add_51_79_groupi_n_4103);
  and csa_tree_add_51_79_groupi_g41171(csa_tree_add_51_79_groupi_n_5053 ,csa_tree_add_51_79_groupi_n_3701 ,csa_tree_add_51_79_groupi_n_4634);
  and csa_tree_add_51_79_groupi_g41172(csa_tree_add_51_79_groupi_n_5052 ,csa_tree_add_51_79_groupi_n_2886 ,csa_tree_add_51_79_groupi_n_4436);
  and csa_tree_add_51_79_groupi_g41173(csa_tree_add_51_79_groupi_n_5051 ,csa_tree_add_51_79_groupi_n_2922 ,csa_tree_add_51_79_groupi_n_3917);
  and csa_tree_add_51_79_groupi_g41174(csa_tree_add_51_79_groupi_n_5050 ,csa_tree_add_51_79_groupi_n_3664 ,csa_tree_add_51_79_groupi_n_4148);
  and csa_tree_add_51_79_groupi_g41175(csa_tree_add_51_79_groupi_n_5049 ,csa_tree_add_51_79_groupi_n_2940 ,csa_tree_add_51_79_groupi_n_3913);
  and csa_tree_add_51_79_groupi_g41176(csa_tree_add_51_79_groupi_n_5048 ,csa_tree_add_51_79_groupi_n_3618 ,csa_tree_add_51_79_groupi_n_4355);
  and csa_tree_add_51_79_groupi_g41177(csa_tree_add_51_79_groupi_n_5047 ,csa_tree_add_51_79_groupi_n_3653 ,csa_tree_add_51_79_groupi_n_3889);
  and csa_tree_add_51_79_groupi_g41178(csa_tree_add_51_79_groupi_n_5046 ,csa_tree_add_51_79_groupi_n_2904 ,csa_tree_add_51_79_groupi_n_4031);
  and csa_tree_add_51_79_groupi_g41179(csa_tree_add_51_79_groupi_n_5045 ,csa_tree_add_51_79_groupi_n_3835 ,csa_tree_add_51_79_groupi_n_4137);
  and csa_tree_add_51_79_groupi_g41180(csa_tree_add_51_79_groupi_n_5044 ,csa_tree_add_51_79_groupi_n_3374 ,csa_tree_add_51_79_groupi_n_4354);
  and csa_tree_add_51_79_groupi_g41181(csa_tree_add_51_79_groupi_n_5043 ,csa_tree_add_51_79_groupi_n_3624 ,csa_tree_add_51_79_groupi_n_4197);
  or csa_tree_add_51_79_groupi_g41182(csa_tree_add_51_79_groupi_n_5042 ,csa_tree_add_51_79_groupi_n_3849 ,csa_tree_add_51_79_groupi_n_3893);
  and csa_tree_add_51_79_groupi_g41183(csa_tree_add_51_79_groupi_n_5041 ,csa_tree_add_51_79_groupi_n_3663 ,csa_tree_add_51_79_groupi_n_4196);
  and csa_tree_add_51_79_groupi_g41184(csa_tree_add_51_79_groupi_n_5040 ,csa_tree_add_51_79_groupi_n_3015 ,csa_tree_add_51_79_groupi_n_3898);
  and csa_tree_add_51_79_groupi_g41185(csa_tree_add_51_79_groupi_n_5039 ,csa_tree_add_51_79_groupi_n_3626 ,csa_tree_add_51_79_groupi_n_4204);
  and csa_tree_add_51_79_groupi_g41186(csa_tree_add_51_79_groupi_n_5038 ,csa_tree_add_51_79_groupi_n_3025 ,csa_tree_add_51_79_groupi_n_3895);
  and csa_tree_add_51_79_groupi_g41187(csa_tree_add_51_79_groupi_n_5037 ,csa_tree_add_51_79_groupi_n_3601 ,csa_tree_add_51_79_groupi_n_4208);
  and csa_tree_add_51_79_groupi_g41188(csa_tree_add_51_79_groupi_n_5036 ,csa_tree_add_51_79_groupi_n_3694 ,csa_tree_add_51_79_groupi_n_4695);
  and csa_tree_add_51_79_groupi_g41189(csa_tree_add_51_79_groupi_n_5034 ,csa_tree_add_51_79_groupi_n_3137 ,csa_tree_add_51_79_groupi_n_4322);
  and csa_tree_add_51_79_groupi_g41190(csa_tree_add_51_79_groupi_n_5033 ,csa_tree_add_51_79_groupi_n_3853 ,csa_tree_add_51_79_groupi_n_4710);
  and csa_tree_add_51_79_groupi_g41191(csa_tree_add_51_79_groupi_n_5032 ,csa_tree_add_51_79_groupi_n_3667 ,csa_tree_add_51_79_groupi_n_4184);
  and csa_tree_add_51_79_groupi_g41192(csa_tree_add_51_79_groupi_n_5031 ,csa_tree_add_51_79_groupi_n_3838 ,csa_tree_add_51_79_groupi_n_4326);
  and csa_tree_add_51_79_groupi_g41193(csa_tree_add_51_79_groupi_n_5030 ,csa_tree_add_51_79_groupi_n_2983 ,csa_tree_add_51_79_groupi_n_3886);
  and csa_tree_add_51_79_groupi_g41194(csa_tree_add_51_79_groupi_n_5029 ,csa_tree_add_51_79_groupi_n_3351 ,csa_tree_add_51_79_groupi_n_3884);
  and csa_tree_add_51_79_groupi_g41195(csa_tree_add_51_79_groupi_n_5028 ,csa_tree_add_51_79_groupi_n_3702 ,csa_tree_add_51_79_groupi_n_4111);
  and csa_tree_add_51_79_groupi_g41196(csa_tree_add_51_79_groupi_n_5027 ,csa_tree_add_51_79_groupi_n_3350 ,csa_tree_add_51_79_groupi_n_3881);
  and csa_tree_add_51_79_groupi_g41197(csa_tree_add_51_79_groupi_n_5026 ,csa_tree_add_51_79_groupi_n_3121 ,csa_tree_add_51_79_groupi_n_3885);
  and csa_tree_add_51_79_groupi_g41198(csa_tree_add_51_79_groupi_n_5025 ,csa_tree_add_51_79_groupi_n_3655 ,csa_tree_add_51_79_groupi_n_4374);
  and csa_tree_add_51_79_groupi_g41199(csa_tree_add_51_79_groupi_n_5024 ,csa_tree_add_51_79_groupi_n_3695 ,csa_tree_add_51_79_groupi_n_4378);
  and csa_tree_add_51_79_groupi_g41200(csa_tree_add_51_79_groupi_n_5023 ,csa_tree_add_51_79_groupi_n_3844 ,csa_tree_add_51_79_groupi_n_4383);
  and csa_tree_add_51_79_groupi_g41201(csa_tree_add_51_79_groupi_n_5022 ,csa_tree_add_51_79_groupi_n_3843 ,csa_tree_add_51_79_groupi_n_4139);
  and csa_tree_add_51_79_groupi_g41202(csa_tree_add_51_79_groupi_n_5021 ,csa_tree_add_51_79_groupi_n_3652 ,csa_tree_add_51_79_groupi_n_4123);
  and csa_tree_add_51_79_groupi_g41203(csa_tree_add_51_79_groupi_n_5020 ,csa_tree_add_51_79_groupi_n_3670 ,csa_tree_add_51_79_groupi_n_4418);
  and csa_tree_add_51_79_groupi_g41204(csa_tree_add_51_79_groupi_n_5019 ,csa_tree_add_51_79_groupi_n_3611 ,csa_tree_add_51_79_groupi_n_4422);
  and csa_tree_add_51_79_groupi_g41205(csa_tree_add_51_79_groupi_n_5018 ,csa_tree_add_51_79_groupi_n_3665 ,csa_tree_add_51_79_groupi_n_4682);
  and csa_tree_add_51_79_groupi_g41206(csa_tree_add_51_79_groupi_n_5017 ,csa_tree_add_51_79_groupi_n_3677 ,csa_tree_add_51_79_groupi_n_4477);
  and csa_tree_add_51_79_groupi_g41207(csa_tree_add_51_79_groupi_n_5016 ,csa_tree_add_51_79_groupi_n_3668 ,csa_tree_add_51_79_groupi_n_4468);
  and csa_tree_add_51_79_groupi_g41208(csa_tree_add_51_79_groupi_n_5015 ,csa_tree_add_51_79_groupi_n_3636 ,csa_tree_add_51_79_groupi_n_4185);
  and csa_tree_add_51_79_groupi_g41209(csa_tree_add_51_79_groupi_n_5014 ,csa_tree_add_51_79_groupi_n_3835 ,csa_tree_add_51_79_groupi_n_4565);
  and csa_tree_add_51_79_groupi_g41210(csa_tree_add_51_79_groupi_n_5013 ,csa_tree_add_51_79_groupi_n_3662 ,csa_tree_add_51_79_groupi_n_4590);
  and csa_tree_add_51_79_groupi_g41211(csa_tree_add_51_79_groupi_n_5012 ,csa_tree_add_51_79_groupi_n_3684 ,csa_tree_add_51_79_groupi_n_4613);
  and csa_tree_add_51_79_groupi_g41212(csa_tree_add_51_79_groupi_n_5011 ,csa_tree_add_51_79_groupi_n_3679 ,csa_tree_add_51_79_groupi_n_4631);
  and csa_tree_add_51_79_groupi_g41213(csa_tree_add_51_79_groupi_n_5010 ,csa_tree_add_51_79_groupi_n_2938 ,csa_tree_add_51_79_groupi_n_3897);
  and csa_tree_add_51_79_groupi_g41214(csa_tree_add_51_79_groupi_n_5009 ,csa_tree_add_51_79_groupi_n_3614 ,csa_tree_add_51_79_groupi_n_4606);
  and csa_tree_add_51_79_groupi_g41215(csa_tree_add_51_79_groupi_n_5008 ,csa_tree_add_51_79_groupi_n_3625 ,csa_tree_add_51_79_groupi_n_4602);
  and csa_tree_add_51_79_groupi_g41216(csa_tree_add_51_79_groupi_n_5007 ,csa_tree_add_51_79_groupi_n_3678 ,csa_tree_add_51_79_groupi_n_4592);
  and csa_tree_add_51_79_groupi_g41217(csa_tree_add_51_79_groupi_n_5006 ,csa_tree_add_51_79_groupi_n_3683 ,csa_tree_add_51_79_groupi_n_4609);
  and csa_tree_add_51_79_groupi_g41218(csa_tree_add_51_79_groupi_n_5005 ,csa_tree_add_51_79_groupi_n_3676 ,csa_tree_add_51_79_groupi_n_4075);
  and csa_tree_add_51_79_groupi_g41219(csa_tree_add_51_79_groupi_n_5004 ,csa_tree_add_51_79_groupi_n_3860 ,csa_tree_add_51_79_groupi_n_4689);
  and csa_tree_add_51_79_groupi_g41220(csa_tree_add_51_79_groupi_n_5003 ,csa_tree_add_51_79_groupi_n_3604 ,csa_tree_add_51_79_groupi_n_4563);
  and csa_tree_add_51_79_groupi_g41221(csa_tree_add_51_79_groupi_n_5002 ,csa_tree_add_51_79_groupi_n_3686 ,csa_tree_add_51_79_groupi_n_4619);
  and csa_tree_add_51_79_groupi_g41222(csa_tree_add_51_79_groupi_n_5001 ,csa_tree_add_51_79_groupi_n_3600 ,csa_tree_add_51_79_groupi_n_4535);
  and csa_tree_add_51_79_groupi_g41223(csa_tree_add_51_79_groupi_n_5000 ,csa_tree_add_51_79_groupi_n_3635 ,csa_tree_add_51_79_groupi_n_4519);
  and csa_tree_add_51_79_groupi_g41224(csa_tree_add_51_79_groupi_n_4999 ,csa_tree_add_51_79_groupi_n_3687 ,csa_tree_add_51_79_groupi_n_4629);
  and csa_tree_add_51_79_groupi_g41225(csa_tree_add_51_79_groupi_n_4998 ,csa_tree_add_51_79_groupi_n_3673 ,csa_tree_add_51_79_groupi_n_4504);
  and csa_tree_add_51_79_groupi_g41226(csa_tree_add_51_79_groupi_n_4997 ,csa_tree_add_51_79_groupi_n_3692 ,csa_tree_add_51_79_groupi_n_4661);
  and csa_tree_add_51_79_groupi_g41227(csa_tree_add_51_79_groupi_n_4996 ,csa_tree_add_51_79_groupi_n_3621 ,csa_tree_add_51_79_groupi_n_4167);
  and csa_tree_add_51_79_groupi_g41228(csa_tree_add_51_79_groupi_n_4995 ,csa_tree_add_51_79_groupi_n_3671 ,csa_tree_add_51_79_groupi_n_4485);
  and csa_tree_add_51_79_groupi_g41229(csa_tree_add_51_79_groupi_n_4994 ,csa_tree_add_51_79_groupi_n_3675 ,csa_tree_add_51_79_groupi_n_4198);
  and csa_tree_add_51_79_groupi_g41230(csa_tree_add_51_79_groupi_n_4993 ,csa_tree_add_51_79_groupi_n_3672 ,csa_tree_add_51_79_groupi_n_4493);
  and csa_tree_add_51_79_groupi_g41231(csa_tree_add_51_79_groupi_n_4992 ,csa_tree_add_51_79_groupi_n_3700 ,csa_tree_add_51_79_groupi_n_4664);
  and csa_tree_add_51_79_groupi_g41232(csa_tree_add_51_79_groupi_n_4991 ,csa_tree_add_51_79_groupi_n_3640 ,csa_tree_add_51_79_groupi_n_4199);
  and csa_tree_add_51_79_groupi_g41233(csa_tree_add_51_79_groupi_n_4990 ,csa_tree_add_51_79_groupi_n_3632 ,csa_tree_add_51_79_groupi_n_4124);
  and csa_tree_add_51_79_groupi_g41234(csa_tree_add_51_79_groupi_n_4989 ,csa_tree_add_51_79_groupi_n_3860 ,csa_tree_add_51_79_groupi_n_4166);
  and csa_tree_add_51_79_groupi_g41235(csa_tree_add_51_79_groupi_n_4987 ,csa_tree_add_51_79_groupi_n_3669 ,csa_tree_add_51_79_groupi_n_3964);
  and csa_tree_add_51_79_groupi_g41236(csa_tree_add_51_79_groupi_n_4986 ,csa_tree_add_51_79_groupi_n_3697 ,csa_tree_add_51_79_groupi_n_4115);
  and csa_tree_add_51_79_groupi_g41237(csa_tree_add_51_79_groupi_n_4985 ,csa_tree_add_51_79_groupi_n_3843 ,csa_tree_add_51_79_groupi_n_4451);
  and csa_tree_add_51_79_groupi_g41238(csa_tree_add_51_79_groupi_n_4984 ,csa_tree_add_51_79_groupi_n_3661 ,csa_tree_add_51_79_groupi_n_4431);
  and csa_tree_add_51_79_groupi_g41239(csa_tree_add_51_79_groupi_n_4983 ,csa_tree_add_51_79_groupi_n_3651 ,csa_tree_add_51_79_groupi_n_4429);
  and csa_tree_add_51_79_groupi_g41240(csa_tree_add_51_79_groupi_n_4982 ,csa_tree_add_51_79_groupi_n_3690 ,csa_tree_add_51_79_groupi_n_4028);
  and csa_tree_add_51_79_groupi_g41241(csa_tree_add_51_79_groupi_n_4981 ,csa_tree_add_51_79_groupi_n_3696 ,csa_tree_add_51_79_groupi_n_4680);
  and csa_tree_add_51_79_groupi_g41242(csa_tree_add_51_79_groupi_n_4980 ,csa_tree_add_51_79_groupi_n_3637 ,csa_tree_add_51_79_groupi_n_4155);
  and csa_tree_add_51_79_groupi_g41243(csa_tree_add_51_79_groupi_n_4979 ,csa_tree_add_51_79_groupi_n_3585 ,csa_tree_add_51_79_groupi_n_4416);
  and csa_tree_add_51_79_groupi_g41244(csa_tree_add_51_79_groupi_n_4978 ,csa_tree_add_51_79_groupi_n_3834 ,csa_tree_add_51_79_groupi_n_4351);
  and csa_tree_add_51_79_groupi_g41245(csa_tree_add_51_79_groupi_n_4977 ,csa_tree_add_51_79_groupi_n_3147 ,csa_tree_add_51_79_groupi_n_4160);
  and csa_tree_add_51_79_groupi_g41246(csa_tree_add_51_79_groupi_n_4976 ,csa_tree_add_51_79_groupi_n_3647 ,csa_tree_add_51_79_groupi_n_4052);
  and csa_tree_add_51_79_groupi_g41247(csa_tree_add_51_79_groupi_n_4975 ,csa_tree_add_51_79_groupi_n_3617 ,csa_tree_add_51_79_groupi_n_4380);
  and csa_tree_add_51_79_groupi_g41248(csa_tree_add_51_79_groupi_n_4974 ,csa_tree_add_51_79_groupi_n_3838 ,csa_tree_add_51_79_groupi_n_4645);
  and csa_tree_add_51_79_groupi_g41249(csa_tree_add_51_79_groupi_n_4973 ,csa_tree_add_51_79_groupi_n_3853 ,csa_tree_add_51_79_groupi_n_4170);
  and csa_tree_add_51_79_groupi_g41250(csa_tree_add_51_79_groupi_n_4972 ,csa_tree_add_51_79_groupi_n_3620 ,csa_tree_add_51_79_groupi_n_4122);
  and csa_tree_add_51_79_groupi_g41251(csa_tree_add_51_79_groupi_n_4971 ,csa_tree_add_51_79_groupi_n_3629 ,csa_tree_add_51_79_groupi_n_4359);
  and csa_tree_add_51_79_groupi_g41252(csa_tree_add_51_79_groupi_n_4970 ,csa_tree_add_51_79_groupi_n_3837 ,csa_tree_add_51_79_groupi_n_4038);
  and csa_tree_add_51_79_groupi_g41253(csa_tree_add_51_79_groupi_n_4969 ,csa_tree_add_51_79_groupi_n_3150 ,csa_tree_add_51_79_groupi_n_4022);
  and csa_tree_add_51_79_groupi_g41254(csa_tree_add_51_79_groupi_n_4968 ,csa_tree_add_51_79_groupi_n_3837 ,csa_tree_add_51_79_groupi_n_4034);
  and csa_tree_add_51_79_groupi_g41255(csa_tree_add_51_79_groupi_n_4966 ,csa_tree_add_51_79_groupi_n_3118 ,csa_tree_add_51_79_groupi_n_3887);
  and csa_tree_add_51_79_groupi_g41256(csa_tree_add_51_79_groupi_n_4965 ,csa_tree_add_51_79_groupi_n_3685 ,csa_tree_add_51_79_groupi_n_4327);
  and csa_tree_add_51_79_groupi_g41257(csa_tree_add_51_79_groupi_n_4964 ,csa_tree_add_51_79_groupi_n_3839 ,csa_tree_add_51_79_groupi_n_4503);
  and csa_tree_add_51_79_groupi_g41258(csa_tree_add_51_79_groupi_n_4962 ,csa_tree_add_51_79_groupi_n_3102 ,csa_tree_add_51_79_groupi_n_4178);
  and csa_tree_add_51_79_groupi_g41259(csa_tree_add_51_79_groupi_n_4960 ,csa_tree_add_51_79_groupi_n_3630 ,csa_tree_add_51_79_groupi_n_4312);
  and csa_tree_add_51_79_groupi_g41260(csa_tree_add_51_79_groupi_n_4959 ,csa_tree_add_51_79_groupi_n_2959 ,csa_tree_add_51_79_groupi_n_4169);
  and csa_tree_add_51_79_groupi_g41261(csa_tree_add_51_79_groupi_n_4957 ,csa_tree_add_51_79_groupi_n_3083 ,csa_tree_add_51_79_groupi_n_3891);
  and csa_tree_add_51_79_groupi_g41262(csa_tree_add_51_79_groupi_n_4955 ,csa_tree_add_51_79_groupi_n_3698 ,csa_tree_add_51_79_groupi_n_4217);
  and csa_tree_add_51_79_groupi_g41263(csa_tree_add_51_79_groupi_n_4954 ,csa_tree_add_51_79_groupi_n_3063 ,csa_tree_add_51_79_groupi_n_4142);
  and csa_tree_add_51_79_groupi_g41264(csa_tree_add_51_79_groupi_n_4953 ,csa_tree_add_51_79_groupi_n_3639 ,csa_tree_add_51_79_groupi_n_4597);
  and csa_tree_add_51_79_groupi_g41265(csa_tree_add_51_79_groupi_n_4952 ,csa_tree_add_51_79_groupi_n_3622 ,csa_tree_add_51_79_groupi_n_4206);
  and csa_tree_add_51_79_groupi_g41266(csa_tree_add_51_79_groupi_n_4951 ,csa_tree_add_51_79_groupi_n_3064 ,csa_tree_add_51_79_groupi_n_3894);
  and csa_tree_add_51_79_groupi_g41267(csa_tree_add_51_79_groupi_n_4950 ,csa_tree_add_51_79_groupi_n_3020 ,csa_tree_add_51_79_groupi_n_3896);
  and csa_tree_add_51_79_groupi_g41268(csa_tree_add_51_79_groupi_n_4949 ,csa_tree_add_51_79_groupi_n_2933 ,csa_tree_add_51_79_groupi_n_3901);
  and csa_tree_add_51_79_groupi_g41269(csa_tree_add_51_79_groupi_n_4948 ,csa_tree_add_51_79_groupi_n_3689 ,csa_tree_add_51_79_groupi_n_4332);
  and csa_tree_add_51_79_groupi_g41270(csa_tree_add_51_79_groupi_n_4947 ,csa_tree_add_51_79_groupi_n_3666 ,csa_tree_add_51_79_groupi_n_4190);
  and csa_tree_add_51_79_groupi_g41271(csa_tree_add_51_79_groupi_n_4946 ,csa_tree_add_51_79_groupi_n_3836 ,csa_tree_add_51_79_groupi_n_4189);
  and csa_tree_add_51_79_groupi_g41272(csa_tree_add_51_79_groupi_n_4944 ,csa_tree_add_51_79_groupi_n_3631 ,csa_tree_add_51_79_groupi_n_4162);
  and csa_tree_add_51_79_groupi_g41273(csa_tree_add_51_79_groupi_n_4943 ,csa_tree_add_51_79_groupi_n_3551 ,csa_tree_add_51_79_groupi_n_3902);
  and csa_tree_add_51_79_groupi_g41274(csa_tree_add_51_79_groupi_n_4942 ,csa_tree_add_51_79_groupi_n_3344 ,csa_tree_add_51_79_groupi_n_3904);
  and csa_tree_add_51_79_groupi_g41275(csa_tree_add_51_79_groupi_n_4941 ,csa_tree_add_51_79_groupi_n_3373 ,csa_tree_add_51_79_groupi_n_3900);
  and csa_tree_add_51_79_groupi_g41276(csa_tree_add_51_79_groupi_n_4940 ,csa_tree_add_51_79_groupi_n_3619 ,csa_tree_add_51_79_groupi_n_4154);
  and csa_tree_add_51_79_groupi_g41277(csa_tree_add_51_79_groupi_n_4939 ,csa_tree_add_51_79_groupi_n_2947 ,csa_tree_add_51_79_groupi_n_3912);
  and csa_tree_add_51_79_groupi_g41278(csa_tree_add_51_79_groupi_n_4938 ,csa_tree_add_51_79_groupi_n_3602 ,csa_tree_add_51_79_groupi_n_4168);
  and csa_tree_add_51_79_groupi_g41279(csa_tree_add_51_79_groupi_n_4937 ,csa_tree_add_51_79_groupi_n_3643 ,csa_tree_add_51_79_groupi_n_4474);
  and csa_tree_add_51_79_groupi_g41280(csa_tree_add_51_79_groupi_n_4936 ,csa_tree_add_51_79_groupi_n_2939 ,csa_tree_add_51_79_groupi_n_3914);
  and csa_tree_add_51_79_groupi_g41281(csa_tree_add_51_79_groupi_n_4935 ,csa_tree_add_51_79_groupi_n_3841 ,csa_tree_add_51_79_groupi_n_4462);
  and csa_tree_add_51_79_groupi_g41282(csa_tree_add_51_79_groupi_n_4934 ,csa_tree_add_51_79_groupi_n_3607 ,csa_tree_add_51_79_groupi_n_4132);
  and csa_tree_add_51_79_groupi_g41283(csa_tree_add_51_79_groupi_n_4933 ,csa_tree_add_51_79_groupi_n_3586 ,csa_tree_add_51_79_groupi_n_4108);
  and csa_tree_add_51_79_groupi_g41284(csa_tree_add_51_79_groupi_n_4932 ,csa_tree_add_51_79_groupi_n_3658 ,csa_tree_add_51_79_groupi_n_4105);
  and csa_tree_add_51_79_groupi_g41285(csa_tree_add_51_79_groupi_n_4930 ,csa_tree_add_51_79_groupi_n_2887 ,csa_tree_add_51_79_groupi_n_3918);
  and csa_tree_add_51_79_groupi_g41286(csa_tree_add_51_79_groupi_n_4929 ,csa_tree_add_51_79_groupi_n_3633 ,csa_tree_add_51_79_groupi_n_4415);
  and csa_tree_add_51_79_groupi_g41287(csa_tree_add_51_79_groupi_n_4928 ,csa_tree_add_51_79_groupi_n_2888 ,csa_tree_add_51_79_groupi_n_3919);
  and csa_tree_add_51_79_groupi_g41288(csa_tree_add_51_79_groupi_n_4927 ,csa_tree_add_51_79_groupi_n_3660 ,csa_tree_add_51_79_groupi_n_4102);
  and csa_tree_add_51_79_groupi_g41289(csa_tree_add_51_79_groupi_n_4926 ,csa_tree_add_51_79_groupi_n_2889 ,csa_tree_add_51_79_groupi_n_3923);
  and csa_tree_add_51_79_groupi_g41290(csa_tree_add_51_79_groupi_n_4925 ,csa_tree_add_51_79_groupi_n_3609 ,csa_tree_add_51_79_groupi_n_4100);
  and csa_tree_add_51_79_groupi_g41291(csa_tree_add_51_79_groupi_n_4924 ,csa_tree_add_51_79_groupi_n_3641 ,csa_tree_add_51_79_groupi_n_4099);
  or csa_tree_add_51_79_groupi_g41292(csa_tree_add_51_79_groupi_n_4922 ,csa_tree_add_51_79_groupi_n_3366 ,csa_tree_add_51_79_groupi_n_3920);
  and csa_tree_add_51_79_groupi_g41293(csa_tree_add_51_79_groupi_n_4921 ,csa_tree_add_51_79_groupi_n_3840 ,csa_tree_add_51_79_groupi_n_4187);
  and csa_tree_add_51_79_groupi_g41294(csa_tree_add_51_79_groupi_n_4920 ,csa_tree_add_51_79_groupi_n_2954 ,csa_tree_add_51_79_groupi_n_3927);
  and csa_tree_add_51_79_groupi_g41295(csa_tree_add_51_79_groupi_n_4919 ,csa_tree_add_51_79_groupi_n_3638 ,csa_tree_add_51_79_groupi_n_4454);
  and csa_tree_add_51_79_groupi_g41296(csa_tree_add_51_79_groupi_n_4918 ,csa_tree_add_51_79_groupi_n_3627 ,csa_tree_add_51_79_groupi_n_4599);
  and csa_tree_add_51_79_groupi_g41297(csa_tree_add_51_79_groupi_n_4917 ,csa_tree_add_51_79_groupi_n_3674 ,csa_tree_add_51_79_groupi_n_4083);
  and csa_tree_add_51_79_groupi_g41298(csa_tree_add_51_79_groupi_n_4916 ,csa_tree_add_51_79_groupi_n_3588 ,csa_tree_add_51_79_groupi_n_4126);
  and csa_tree_add_51_79_groupi_g41299(csa_tree_add_51_79_groupi_n_4915 ,csa_tree_add_51_79_groupi_n_3612 ,csa_tree_add_51_79_groupi_n_4584);
  and csa_tree_add_51_79_groupi_g41300(csa_tree_add_51_79_groupi_n_4914 ,csa_tree_add_51_79_groupi_n_2893 ,csa_tree_add_51_79_groupi_n_3933);
  and csa_tree_add_51_79_groupi_g41301(csa_tree_add_51_79_groupi_n_4913 ,csa_tree_add_51_79_groupi_n_3589 ,csa_tree_add_51_79_groupi_n_4593);
  and csa_tree_add_51_79_groupi_g41302(csa_tree_add_51_79_groupi_n_4912 ,csa_tree_add_51_79_groupi_n_3430 ,csa_tree_add_51_79_groupi_n_3934);
  and csa_tree_add_51_79_groupi_g41303(csa_tree_add_51_79_groupi_n_4911 ,csa_tree_add_51_79_groupi_n_3634 ,csa_tree_add_51_79_groupi_n_4069);
  and csa_tree_add_51_79_groupi_g41304(csa_tree_add_51_79_groupi_n_4910 ,csa_tree_add_51_79_groupi_n_3567 ,csa_tree_add_51_79_groupi_n_3938);
  and csa_tree_add_51_79_groupi_g41305(csa_tree_add_51_79_groupi_n_4909 ,csa_tree_add_51_79_groupi_n_3452 ,csa_tree_add_51_79_groupi_n_3939);
  and csa_tree_add_51_79_groupi_g41306(csa_tree_add_51_79_groupi_n_4908 ,csa_tree_add_51_79_groupi_n_2895 ,csa_tree_add_51_79_groupi_n_3940);
  and csa_tree_add_51_79_groupi_g41307(csa_tree_add_51_79_groupi_n_4907 ,csa_tree_add_51_79_groupi_n_3703 ,csa_tree_add_51_79_groupi_n_4048);
  and csa_tree_add_51_79_groupi_g41308(csa_tree_add_51_79_groupi_n_4906 ,csa_tree_add_51_79_groupi_n_3616 ,csa_tree_add_51_79_groupi_n_4127);
  and csa_tree_add_51_79_groupi_g41309(csa_tree_add_51_79_groupi_n_4905 ,csa_tree_add_51_79_groupi_n_3691 ,csa_tree_add_51_79_groupi_n_4674);
  and csa_tree_add_51_79_groupi_g41310(csa_tree_add_51_79_groupi_n_4904 ,csa_tree_add_51_79_groupi_n_3862 ,csa_tree_add_51_79_groupi_n_3937);
  and csa_tree_add_51_79_groupi_g41311(csa_tree_add_51_79_groupi_n_4903 ,csa_tree_add_51_79_groupi_n_3597 ,csa_tree_add_51_79_groupi_n_4146);
  and csa_tree_add_51_79_groupi_g41312(csa_tree_add_51_79_groupi_n_4902 ,csa_tree_add_51_79_groupi_n_3615 ,csa_tree_add_51_79_groupi_n_4445);
  and csa_tree_add_51_79_groupi_g41313(csa_tree_add_51_79_groupi_n_4901 ,csa_tree_add_51_79_groupi_n_3605 ,csa_tree_add_51_79_groupi_n_4407);
  and csa_tree_add_51_79_groupi_g41314(csa_tree_add_51_79_groupi_n_4900 ,csa_tree_add_51_79_groupi_n_2985 ,csa_tree_add_51_79_groupi_n_4382);
  and csa_tree_add_51_79_groupi_g41315(csa_tree_add_51_79_groupi_n_4899 ,csa_tree_add_51_79_groupi_n_3681 ,csa_tree_add_51_79_groupi_n_4072);
  and csa_tree_add_51_79_groupi_g41316(csa_tree_add_51_79_groupi_n_4898 ,csa_tree_add_51_79_groupi_n_3840 ,csa_tree_add_51_79_groupi_n_4439);
  and csa_tree_add_51_79_groupi_g41317(csa_tree_add_51_79_groupi_n_4897 ,csa_tree_add_51_79_groupi_n_3841 ,csa_tree_add_51_79_groupi_n_4394);
  and csa_tree_add_51_79_groupi_g41318(csa_tree_add_51_79_groupi_n_4895 ,csa_tree_add_51_79_groupi_n_3376 ,csa_tree_add_51_79_groupi_n_4461);
  and csa_tree_add_51_79_groupi_g41319(csa_tree_add_51_79_groupi_n_4894 ,csa_tree_add_51_79_groupi_n_3656 ,csa_tree_add_51_79_groupi_n_4009);
  and csa_tree_add_51_79_groupi_g41320(csa_tree_add_51_79_groupi_n_4893 ,csa_tree_add_51_79_groupi_n_3594 ,csa_tree_add_51_79_groupi_n_4004);
  and csa_tree_add_51_79_groupi_g41321(csa_tree_add_51_79_groupi_n_4892 ,csa_tree_add_51_79_groupi_n_3433 ,csa_tree_add_51_79_groupi_n_4536);
  and csa_tree_add_51_79_groupi_g41322(csa_tree_add_51_79_groupi_n_4890 ,csa_tree_add_51_79_groupi_n_3591 ,csa_tree_add_51_79_groupi_n_3994);
  and csa_tree_add_51_79_groupi_g41323(csa_tree_add_51_79_groupi_n_4889 ,csa_tree_add_51_79_groupi_n_3598 ,csa_tree_add_51_79_groupi_n_3916);
  and csa_tree_add_51_79_groupi_g41324(csa_tree_add_51_79_groupi_n_4888 ,csa_tree_add_51_79_groupi_n_2905 ,csa_tree_add_51_79_groupi_n_3952);
  and csa_tree_add_51_79_groupi_g41325(csa_tree_add_51_79_groupi_n_4887 ,csa_tree_add_51_79_groupi_n_3372 ,csa_tree_add_51_79_groupi_n_3946);
  and csa_tree_add_51_79_groupi_g41326(csa_tree_add_51_79_groupi_n_4886 ,csa_tree_add_51_79_groupi_n_2906 ,csa_tree_add_51_79_groupi_n_3954);
  and csa_tree_add_51_79_groupi_g41327(csa_tree_add_51_79_groupi_n_4885 ,csa_tree_add_51_79_groupi_n_3593 ,csa_tree_add_51_79_groupi_n_3929);
  and csa_tree_add_51_79_groupi_g41328(csa_tree_add_51_79_groupi_n_4884 ,csa_tree_add_51_79_groupi_n_3592 ,csa_tree_add_51_79_groupi_n_3924);
  and csa_tree_add_51_79_groupi_g41329(csa_tree_add_51_79_groupi_n_4883 ,csa_tree_add_51_79_groupi_n_2908 ,csa_tree_add_51_79_groupi_n_3957);
  and csa_tree_add_51_79_groupi_g41330(csa_tree_add_51_79_groupi_n_4882 ,csa_tree_add_51_79_groupi_n_3613 ,csa_tree_add_51_79_groupi_n_3888);
  and csa_tree_add_51_79_groupi_g41331(csa_tree_add_51_79_groupi_n_4881 ,csa_tree_add_51_79_groupi_n_3587 ,csa_tree_add_51_79_groupi_n_4544);
  and csa_tree_add_51_79_groupi_g41332(csa_tree_add_51_79_groupi_n_4880 ,csa_tree_add_51_79_groupi_n_3429 ,csa_tree_add_51_79_groupi_n_3958);
  and csa_tree_add_51_79_groupi_g41333(csa_tree_add_51_79_groupi_n_4879 ,csa_tree_add_51_79_groupi_n_2909 ,csa_tree_add_51_79_groupi_n_3959);
  and csa_tree_add_51_79_groupi_g41334(csa_tree_add_51_79_groupi_n_4878 ,csa_tree_add_51_79_groupi_n_2911 ,csa_tree_add_51_79_groupi_n_3961);
  and csa_tree_add_51_79_groupi_g41335(csa_tree_add_51_79_groupi_n_4877 ,csa_tree_add_51_79_groupi_n_3395 ,csa_tree_add_51_79_groupi_n_3962);
  and csa_tree_add_51_79_groupi_g41336(csa_tree_add_51_79_groupi_n_4876 ,csa_tree_add_51_79_groupi_n_3409 ,csa_tree_add_51_79_groupi_n_3968);
  and csa_tree_add_51_79_groupi_g41337(csa_tree_add_51_79_groupi_n_4875 ,csa_tree_add_51_79_groupi_n_3483 ,csa_tree_add_51_79_groupi_n_3970);
  or csa_tree_add_51_79_groupi_g41338(csa_tree_add_51_79_groupi_n_4873 ,csa_tree_add_51_79_groupi_n_3368 ,csa_tree_add_51_79_groupi_n_3969);
  and csa_tree_add_51_79_groupi_g41339(csa_tree_add_51_79_groupi_n_4872 ,csa_tree_add_51_79_groupi_n_3498 ,csa_tree_add_51_79_groupi_n_3972);
  and csa_tree_add_51_79_groupi_g41340(csa_tree_add_51_79_groupi_n_4871 ,csa_tree_add_51_79_groupi_n_3657 ,csa_tree_add_51_79_groupi_n_3974);
  and csa_tree_add_51_79_groupi_g41341(csa_tree_add_51_79_groupi_n_4870 ,csa_tree_add_51_79_groupi_n_2915 ,csa_tree_add_51_79_groupi_n_3975);
  and csa_tree_add_51_79_groupi_g41342(csa_tree_add_51_79_groupi_n_4868 ,csa_tree_add_51_79_groupi_n_2917 ,csa_tree_add_51_79_groupi_n_3977);
  and csa_tree_add_51_79_groupi_g41343(csa_tree_add_51_79_groupi_n_4867 ,csa_tree_add_51_79_groupi_n_3128 ,csa_tree_add_51_79_groupi_n_3978);
  and csa_tree_add_51_79_groupi_g41344(csa_tree_add_51_79_groupi_n_4866 ,csa_tree_add_51_79_groupi_n_3101 ,csa_tree_add_51_79_groupi_n_3981);
  and csa_tree_add_51_79_groupi_g41345(csa_tree_add_51_79_groupi_n_4864 ,csa_tree_add_51_79_groupi_n_3343 ,csa_tree_add_51_79_groupi_n_4023);
  or csa_tree_add_51_79_groupi_g41346(csa_tree_add_51_79_groupi_n_4862 ,csa_tree_add_51_79_groupi_n_3364 ,csa_tree_add_51_79_groupi_n_4481);
  and csa_tree_add_51_79_groupi_g41347(csa_tree_add_51_79_groupi_n_4861 ,csa_tree_add_51_79_groupi_n_2900 ,csa_tree_add_51_79_groupi_n_4537);
  and csa_tree_add_51_79_groupi_g41348(csa_tree_add_51_79_groupi_n_4860 ,csa_tree_add_51_79_groupi_n_3357 ,csa_tree_add_51_79_groupi_n_3980);
  and csa_tree_add_51_79_groupi_g41349(csa_tree_add_51_79_groupi_n_4859 ,csa_tree_add_51_79_groupi_n_3573 ,csa_tree_add_51_79_groupi_n_3899);
  or csa_tree_add_51_79_groupi_g41350(csa_tree_add_51_79_groupi_n_4857 ,csa_tree_add_51_79_groupi_n_3358 ,csa_tree_add_51_79_groupi_n_3987);
  and csa_tree_add_51_79_groupi_g41351(csa_tree_add_51_79_groupi_n_4856 ,csa_tree_add_51_79_groupi_n_2928 ,csa_tree_add_51_79_groupi_n_3990);
  and csa_tree_add_51_79_groupi_g41352(csa_tree_add_51_79_groupi_n_4854 ,csa_tree_add_51_79_groupi_n_2902 ,csa_tree_add_51_79_groupi_n_3993);
  and csa_tree_add_51_79_groupi_g41353(csa_tree_add_51_79_groupi_n_4853 ,csa_tree_add_51_79_groupi_n_2901 ,csa_tree_add_51_79_groupi_n_4411);
  and csa_tree_add_51_79_groupi_g41354(csa_tree_add_51_79_groupi_n_4852 ,csa_tree_add_51_79_groupi_n_3576 ,csa_tree_add_51_79_groupi_n_4041);
  and csa_tree_add_51_79_groupi_g41355(csa_tree_add_51_79_groupi_n_4851 ,csa_tree_add_51_79_groupi_n_3151 ,csa_tree_add_51_79_groupi_n_3997);
  and csa_tree_add_51_79_groupi_g41356(csa_tree_add_51_79_groupi_n_4850 ,csa_tree_add_51_79_groupi_n_2930 ,csa_tree_add_51_79_groupi_n_3915);
  and csa_tree_add_51_79_groupi_g41357(csa_tree_add_51_79_groupi_n_4849 ,csa_tree_add_51_79_groupi_n_2934 ,csa_tree_add_51_79_groupi_n_4001);
  and csa_tree_add_51_79_groupi_g41358(csa_tree_add_51_79_groupi_n_4848 ,csa_tree_add_51_79_groupi_n_2935 ,csa_tree_add_51_79_groupi_n_4002);
  and csa_tree_add_51_79_groupi_g41359(csa_tree_add_51_79_groupi_n_4847 ,csa_tree_add_51_79_groupi_n_2936 ,csa_tree_add_51_79_groupi_n_4005);
  and csa_tree_add_51_79_groupi_g41360(csa_tree_add_51_79_groupi_n_4846 ,csa_tree_add_51_79_groupi_n_2941 ,csa_tree_add_51_79_groupi_n_4008);
  and csa_tree_add_51_79_groupi_g41361(csa_tree_add_51_79_groupi_n_4845 ,csa_tree_add_51_79_groupi_n_3107 ,csa_tree_add_51_79_groupi_n_4010);
  and csa_tree_add_51_79_groupi_g41362(csa_tree_add_51_79_groupi_n_4844 ,csa_tree_add_51_79_groupi_n_2924 ,csa_tree_add_51_79_groupi_n_4679);
  and csa_tree_add_51_79_groupi_g41363(csa_tree_add_51_79_groupi_n_4843 ,csa_tree_add_51_79_groupi_n_3526 ,csa_tree_add_51_79_groupi_n_4675);
  and csa_tree_add_51_79_groupi_g41364(csa_tree_add_51_79_groupi_n_4842 ,csa_tree_add_51_79_groupi_n_3153 ,csa_tree_add_51_79_groupi_n_4350);
  and csa_tree_add_51_79_groupi_g41367(csa_tree_add_51_79_groupi_n_4841 ,csa_tree_add_51_79_groupi_n_2958 ,csa_tree_add_51_79_groupi_n_4530);
  and csa_tree_add_51_79_groupi_g41368(csa_tree_add_51_79_groupi_n_4840 ,csa_tree_add_51_79_groupi_n_2956 ,csa_tree_add_51_79_groupi_n_4562);
  and csa_tree_add_51_79_groupi_g41369(csa_tree_add_51_79_groupi_n_4838 ,csa_tree_add_51_79_groupi_n_2981 ,csa_tree_add_51_79_groupi_n_4171);
  and csa_tree_add_51_79_groupi_g41370(csa_tree_add_51_79_groupi_n_4837 ,csa_tree_add_51_79_groupi_n_3503 ,csa_tree_add_51_79_groupi_n_4046);
  and csa_tree_add_51_79_groupi_g41371(csa_tree_add_51_79_groupi_n_4836 ,csa_tree_add_51_79_groupi_n_3529 ,csa_tree_add_51_79_groupi_n_4692);
  and csa_tree_add_51_79_groupi_g41372(csa_tree_add_51_79_groupi_n_4835 ,csa_tree_add_51_79_groupi_n_3435 ,csa_tree_add_51_79_groupi_n_4106);
  or csa_tree_add_51_79_groupi_g41373(csa_tree_add_51_79_groupi_n_4833 ,csa_tree_add_51_79_groupi_n_3352 ,csa_tree_add_51_79_groupi_n_3983);
  and csa_tree_add_51_79_groupi_g41374(csa_tree_add_51_79_groupi_n_4832 ,csa_tree_add_51_79_groupi_n_3044 ,csa_tree_add_51_79_groupi_n_4064);
  and csa_tree_add_51_79_groupi_g41375(csa_tree_add_51_79_groupi_n_4831 ,csa_tree_add_51_79_groupi_n_3516 ,csa_tree_add_51_79_groupi_n_4035);
  and csa_tree_add_51_79_groupi_g41376(csa_tree_add_51_79_groupi_n_4830 ,csa_tree_add_51_79_groupi_n_3047 ,csa_tree_add_51_79_groupi_n_4598);
  and csa_tree_add_51_79_groupi_g41377(csa_tree_add_51_79_groupi_n_4829 ,csa_tree_add_51_79_groupi_n_3111 ,csa_tree_add_51_79_groupi_n_4071);
  and csa_tree_add_51_79_groupi_g41378(csa_tree_add_51_79_groupi_n_4828 ,csa_tree_add_51_79_groupi_n_3396 ,csa_tree_add_51_79_groupi_n_4455);
  and csa_tree_add_51_79_groupi_g41379(csa_tree_add_51_79_groupi_n_4826 ,csa_tree_add_51_79_groupi_n_3484 ,csa_tree_add_51_79_groupi_n_4348);
  and csa_tree_add_51_79_groupi_g41380(csa_tree_add_51_79_groupi_n_4824 ,csa_tree_add_51_79_groupi_n_3373 ,csa_tree_add_51_79_groupi_n_4372);
  and csa_tree_add_51_79_groupi_g41381(csa_tree_add_51_79_groupi_n_4822 ,csa_tree_add_51_79_groupi_n_3505 ,csa_tree_add_51_79_groupi_n_4452);
  and csa_tree_add_51_79_groupi_g41382(csa_tree_add_51_79_groupi_n_4821 ,csa_tree_add_51_79_groupi_n_3545 ,csa_tree_add_51_79_groupi_n_4570);
  and csa_tree_add_51_79_groupi_g41383(csa_tree_add_51_79_groupi_n_4820 ,csa_tree_add_51_79_groupi_n_3610 ,csa_tree_add_51_79_groupi_n_4709);
  and csa_tree_add_51_79_groupi_g41384(csa_tree_add_51_79_groupi_n_4819 ,csa_tree_add_51_79_groupi_n_3515 ,csa_tree_add_51_79_groupi_n_4541);
  and csa_tree_add_51_79_groupi_g41385(csa_tree_add_51_79_groupi_n_4818 ,csa_tree_add_51_79_groupi_n_3084 ,csa_tree_add_51_79_groupi_n_4081);
  and csa_tree_add_51_79_groupi_g41386(csa_tree_add_51_79_groupi_n_4817 ,csa_tree_add_51_79_groupi_n_3417 ,csa_tree_add_51_79_groupi_n_4085);
  and csa_tree_add_51_79_groupi_g41387(csa_tree_add_51_79_groupi_n_4816 ,csa_tree_add_51_79_groupi_n_3018 ,csa_tree_add_51_79_groupi_n_3908);
  and csa_tree_add_51_79_groupi_g41388(csa_tree_add_51_79_groupi_n_4815 ,csa_tree_add_51_79_groupi_n_3404 ,csa_tree_add_51_79_groupi_n_4706);
  and csa_tree_add_51_79_groupi_g41389(csa_tree_add_51_79_groupi_n_4814 ,csa_tree_add_51_79_groupi_n_3467 ,csa_tree_add_51_79_groupi_n_4056);
  and csa_tree_add_51_79_groupi_g41390(csa_tree_add_51_79_groupi_n_4813 ,csa_tree_add_51_79_groupi_n_3377 ,csa_tree_add_51_79_groupi_n_4091);
  and csa_tree_add_51_79_groupi_g41391(csa_tree_add_51_79_groupi_n_4812 ,csa_tree_add_51_79_groupi_n_3008 ,csa_tree_add_51_79_groupi_n_4092);
  and csa_tree_add_51_79_groupi_g41393(csa_tree_add_51_79_groupi_n_4810 ,csa_tree_add_51_79_groupi_n_2975 ,csa_tree_add_51_79_groupi_n_4065);
  and csa_tree_add_51_79_groupi_g41394(csa_tree_add_51_79_groupi_n_4809 ,csa_tree_add_51_79_groupi_n_3583 ,csa_tree_add_51_79_groupi_n_4096);
  and csa_tree_add_51_79_groupi_g41395(csa_tree_add_51_79_groupi_n_4808 ,csa_tree_add_51_79_groupi_n_2919 ,csa_tree_add_51_79_groupi_n_4097);
  xnor csa_tree_add_51_79_groupi_g41396(csa_tree_add_51_79_groupi_n_4807 ,csa_tree_add_51_79_groupi_n_3743 ,csa_tree_add_51_79_groupi_n_3247);
  xnor csa_tree_add_51_79_groupi_g41397(csa_tree_add_51_79_groupi_n_4806 ,csa_tree_add_51_79_groupi_n_3786 ,csa_tree_add_51_79_groupi_n_3250);
  and csa_tree_add_51_79_groupi_g41398(csa_tree_add_51_79_groupi_n_4805 ,csa_tree_add_51_79_groupi_n_3059 ,csa_tree_add_51_79_groupi_n_4363);
  and csa_tree_add_51_79_groupi_g41399(csa_tree_add_51_79_groupi_n_4803 ,csa_tree_add_51_79_groupi_n_3858 ,csa_tree_add_51_79_groupi_n_4164);
  and csa_tree_add_51_79_groupi_g41400(csa_tree_add_51_79_groupi_n_4802 ,csa_tree_add_51_79_groupi_n_2903 ,csa_tree_add_51_79_groupi_n_4470);
  and csa_tree_add_51_79_groupi_g41401(csa_tree_add_51_79_groupi_n_4801 ,csa_tree_add_51_79_groupi_n_3458 ,csa_tree_add_51_79_groupi_n_4341);
  xnor csa_tree_add_51_79_groupi_g41402(csa_tree_add_51_79_groupi_n_4800 ,csa_tree_add_51_79_groupi_n_3744 ,csa_tree_add_51_79_groupi_n_3776);
  and csa_tree_add_51_79_groupi_g41403(csa_tree_add_51_79_groupi_n_4799 ,csa_tree_add_51_79_groupi_n_2963 ,csa_tree_add_51_79_groupi_n_4037);
  and csa_tree_add_51_79_groupi_g41404(csa_tree_add_51_79_groupi_n_4798 ,csa_tree_add_51_79_groupi_n_3391 ,csa_tree_add_51_79_groupi_n_4705);
  and csa_tree_add_51_79_groupi_g41405(csa_tree_add_51_79_groupi_n_4797 ,csa_tree_add_51_79_groupi_n_3852 ,csa_tree_add_51_79_groupi_n_4403);
  and csa_tree_add_51_79_groupi_g41406(csa_tree_add_51_79_groupi_n_4796 ,csa_tree_add_51_79_groupi_n_3078 ,csa_tree_add_51_79_groupi_n_4163);
  and csa_tree_add_51_79_groupi_g41407(csa_tree_add_51_79_groupi_n_4794 ,csa_tree_add_51_79_groupi_n_2925 ,csa_tree_add_51_79_groupi_n_3909);
  and csa_tree_add_51_79_groupi_g41408(csa_tree_add_51_79_groupi_n_4793 ,csa_tree_add_51_79_groupi_n_3040 ,csa_tree_add_51_79_groupi_n_3941);
  or csa_tree_add_51_79_groupi_g41409(csa_tree_add_51_79_groupi_n_4710 ,csa_tree_add_51_79_groupi_n_2759 ,csa_tree_add_51_79_groupi_n_927);
  or csa_tree_add_51_79_groupi_g41410(csa_tree_add_51_79_groupi_n_4709 ,csa_tree_add_51_79_groupi_n_2227 ,csa_tree_add_51_79_groupi_n_426);
  or csa_tree_add_51_79_groupi_g41411(csa_tree_add_51_79_groupi_n_4708 ,csa_tree_add_51_79_groupi_n_2184 ,csa_tree_add_51_79_groupi_n_1008);
  and csa_tree_add_51_79_groupi_g41412(csa_tree_add_51_79_groupi_n_4707 ,csa_tree_add_51_79_groupi_n_3220 ,csa_tree_add_51_79_groupi_n_3258);
  or csa_tree_add_51_79_groupi_g41413(csa_tree_add_51_79_groupi_n_4706 ,csa_tree_add_51_79_groupi_n_2271 ,csa_tree_add_51_79_groupi_n_1068);
  or csa_tree_add_51_79_groupi_g41414(csa_tree_add_51_79_groupi_n_4705 ,csa_tree_add_51_79_groupi_n_2159 ,csa_tree_add_51_79_groupi_n_426);
  or csa_tree_add_51_79_groupi_g41415(csa_tree_add_51_79_groupi_n_4704 ,csa_tree_add_51_79_groupi_n_2057 ,csa_tree_add_51_79_groupi_n_921);
  and csa_tree_add_51_79_groupi_g41416(csa_tree_add_51_79_groupi_n_4703 ,csa_tree_add_51_79_groupi_n_3219 ,csa_tree_add_51_79_groupi_n_3223);
  or csa_tree_add_51_79_groupi_g41417(csa_tree_add_51_79_groupi_n_4702 ,csa_tree_add_51_79_groupi_n_2713 ,csa_tree_add_51_79_groupi_n_942);
  or csa_tree_add_51_79_groupi_g41418(csa_tree_add_51_79_groupi_n_4701 ,csa_tree_add_51_79_groupi_n_3804 ,csa_tree_add_51_79_groupi_n_3210);
  or csa_tree_add_51_79_groupi_g41419(csa_tree_add_51_79_groupi_n_4700 ,csa_tree_add_51_79_groupi_n_2715 ,csa_tree_add_51_79_groupi_n_1002);
  or csa_tree_add_51_79_groupi_g41420(csa_tree_add_51_79_groupi_n_4699 ,csa_tree_add_51_79_groupi_n_2757 ,csa_tree_add_51_79_groupi_n_446);
  or csa_tree_add_51_79_groupi_g41421(csa_tree_add_51_79_groupi_n_4698 ,csa_tree_add_51_79_groupi_n_3222 ,csa_tree_add_51_79_groupi_n_3211);
  or csa_tree_add_51_79_groupi_g41422(csa_tree_add_51_79_groupi_n_4697 ,csa_tree_add_51_79_groupi_n_2137 ,csa_tree_add_51_79_groupi_n_424);
  and csa_tree_add_51_79_groupi_g41423(csa_tree_add_51_79_groupi_n_4696 ,csa_tree_add_51_79_groupi_n_3222 ,csa_tree_add_51_79_groupi_n_3211);
  or csa_tree_add_51_79_groupi_g41424(csa_tree_add_51_79_groupi_n_4695 ,csa_tree_add_51_79_groupi_n_2574 ,csa_tree_add_51_79_groupi_n_936);
  or csa_tree_add_51_79_groupi_g41425(csa_tree_add_51_79_groupi_n_4694 ,csa_tree_add_51_79_groupi_n_2801 ,csa_tree_add_51_79_groupi_n_969);
  nor csa_tree_add_51_79_groupi_g41426(csa_tree_add_51_79_groupi_n_4693 ,csa_tree_add_51_79_groupi_n_2795 ,csa_tree_add_51_79_groupi_n_1038);
  or csa_tree_add_51_79_groupi_g41427(csa_tree_add_51_79_groupi_n_4692 ,csa_tree_add_51_79_groupi_n_2092 ,csa_tree_add_51_79_groupi_n_404);
  or csa_tree_add_51_79_groupi_g41428(csa_tree_add_51_79_groupi_n_4691 ,csa_tree_add_51_79_groupi_n_2658 ,csa_tree_add_51_79_groupi_n_1017);
  or csa_tree_add_51_79_groupi_g41429(csa_tree_add_51_79_groupi_n_4690 ,csa_tree_add_51_79_groupi_n_2268 ,csa_tree_add_51_79_groupi_n_1059);
  or csa_tree_add_51_79_groupi_g41430(csa_tree_add_51_79_groupi_n_4689 ,csa_tree_add_51_79_groupi_n_2047 ,csa_tree_add_51_79_groupi_n_933);
  or csa_tree_add_51_79_groupi_g41431(csa_tree_add_51_79_groupi_n_4688 ,csa_tree_add_51_79_groupi_n_2643 ,csa_tree_add_51_79_groupi_n_1023);
  or csa_tree_add_51_79_groupi_g41432(csa_tree_add_51_79_groupi_n_4687 ,csa_tree_add_51_79_groupi_n_3205 ,csa_tree_add_51_79_groupi_n_3277);
  or csa_tree_add_51_79_groupi_g41433(csa_tree_add_51_79_groupi_n_4686 ,csa_tree_add_51_79_groupi_n_2231 ,csa_tree_add_51_79_groupi_n_1041);
  or csa_tree_add_51_79_groupi_g41434(csa_tree_add_51_79_groupi_n_4685 ,csa_tree_add_51_79_groupi_n_2829 ,csa_tree_add_51_79_groupi_n_966);
  or csa_tree_add_51_79_groupi_g41435(csa_tree_add_51_79_groupi_n_4684 ,csa_tree_add_51_79_groupi_n_2244 ,csa_tree_add_51_79_groupi_n_897);
  or csa_tree_add_51_79_groupi_g41436(csa_tree_add_51_79_groupi_n_4683 ,csa_tree_add_51_79_groupi_n_2266 ,csa_tree_add_51_79_groupi_n_424);
  or csa_tree_add_51_79_groupi_g41437(csa_tree_add_51_79_groupi_n_4682 ,csa_tree_add_51_79_groupi_n_2625 ,csa_tree_add_51_79_groupi_n_490);
  or csa_tree_add_51_79_groupi_g41438(csa_tree_add_51_79_groupi_n_4681 ,csa_tree_add_51_79_groupi_n_2290 ,csa_tree_add_51_79_groupi_n_981);
  or csa_tree_add_51_79_groupi_g41439(csa_tree_add_51_79_groupi_n_4680 ,csa_tree_add_51_79_groupi_n_2113 ,csa_tree_add_51_79_groupi_n_909);
  or csa_tree_add_51_79_groupi_g41440(csa_tree_add_51_79_groupi_n_4679 ,csa_tree_add_51_79_groupi_n_2156 ,csa_tree_add_51_79_groupi_n_1053);
  or csa_tree_add_51_79_groupi_g41441(csa_tree_add_51_79_groupi_n_4678 ,csa_tree_add_51_79_groupi_n_2823 ,csa_tree_add_51_79_groupi_n_975);
  or csa_tree_add_51_79_groupi_g41442(csa_tree_add_51_79_groupi_n_4677 ,csa_tree_add_51_79_groupi_n_2286 ,csa_tree_add_51_79_groupi_n_978);
  or csa_tree_add_51_79_groupi_g41443(csa_tree_add_51_79_groupi_n_4676 ,csa_tree_add_51_79_groupi_n_2128 ,csa_tree_add_51_79_groupi_n_1005);
  or csa_tree_add_51_79_groupi_g41444(csa_tree_add_51_79_groupi_n_4675 ,csa_tree_add_51_79_groupi_n_2850 ,csa_tree_add_51_79_groupi_n_903);
  or csa_tree_add_51_79_groupi_g41445(csa_tree_add_51_79_groupi_n_4674 ,csa_tree_add_51_79_groupi_n_2870 ,csa_tree_add_51_79_groupi_n_924);
  or csa_tree_add_51_79_groupi_g41446(csa_tree_add_51_79_groupi_n_4673 ,csa_tree_add_51_79_groupi_n_2679 ,csa_tree_add_51_79_groupi_n_512);
  or csa_tree_add_51_79_groupi_g41447(csa_tree_add_51_79_groupi_n_4672 ,csa_tree_add_51_79_groupi_n_2860 ,csa_tree_add_51_79_groupi_n_954);
  or csa_tree_add_51_79_groupi_g41448(csa_tree_add_51_79_groupi_n_4671 ,csa_tree_add_51_79_groupi_n_2212 ,csa_tree_add_51_79_groupi_n_1044);
  or csa_tree_add_51_79_groupi_g41449(csa_tree_add_51_79_groupi_n_4670 ,csa_tree_add_51_79_groupi_n_2207 ,csa_tree_add_51_79_groupi_n_1011);
  or csa_tree_add_51_79_groupi_g41450(csa_tree_add_51_79_groupi_n_4669 ,csa_tree_add_51_79_groupi_n_2165 ,csa_tree_add_51_79_groupi_n_1032);
  or csa_tree_add_51_79_groupi_g41451(csa_tree_add_51_79_groupi_n_4668 ,csa_tree_add_51_79_groupi_n_3207 ,csa_tree_add_51_79_groupi_n_3224);
  or csa_tree_add_51_79_groupi_g41452(csa_tree_add_51_79_groupi_n_4667 ,csa_tree_add_51_79_groupi_n_2233 ,csa_tree_add_51_79_groupi_n_1035);
  or csa_tree_add_51_79_groupi_g41453(csa_tree_add_51_79_groupi_n_4666 ,csa_tree_add_51_79_groupi_n_2280 ,csa_tree_add_51_79_groupi_n_930);
  or csa_tree_add_51_79_groupi_g41454(csa_tree_add_51_79_groupi_n_4665 ,csa_tree_add_51_79_groupi_n_2239 ,csa_tree_add_51_79_groupi_n_408);
  or csa_tree_add_51_79_groupi_g41455(csa_tree_add_51_79_groupi_n_4664 ,csa_tree_add_51_79_groupi_n_2880 ,csa_tree_add_51_79_groupi_n_498);
  or csa_tree_add_51_79_groupi_g41456(csa_tree_add_51_79_groupi_n_4663 ,csa_tree_add_51_79_groupi_n_2802 ,csa_tree_add_51_79_groupi_n_422);
  or csa_tree_add_51_79_groupi_g41457(csa_tree_add_51_79_groupi_n_4662 ,csa_tree_add_51_79_groupi_n_2878 ,csa_tree_add_51_79_groupi_n_996);
  or csa_tree_add_51_79_groupi_g41458(csa_tree_add_51_79_groupi_n_4661 ,csa_tree_add_51_79_groupi_n_2877 ,csa_tree_add_51_79_groupi_n_894);
  or csa_tree_add_51_79_groupi_g41459(csa_tree_add_51_79_groupi_n_4660 ,csa_tree_add_51_79_groupi_n_2145 ,csa_tree_add_51_79_groupi_n_960);
  or csa_tree_add_51_79_groupi_g41460(csa_tree_add_51_79_groupi_n_4659 ,csa_tree_add_51_79_groupi_n_2876 ,csa_tree_add_51_79_groupi_n_948);
  or csa_tree_add_51_79_groupi_g41461(csa_tree_add_51_79_groupi_n_4658 ,csa_tree_add_51_79_groupi_n_2729 ,csa_tree_add_51_79_groupi_n_1020);
  or csa_tree_add_51_79_groupi_g41462(csa_tree_add_51_79_groupi_n_4657 ,csa_tree_add_51_79_groupi_n_2169 ,csa_tree_add_51_79_groupi_n_516);
  or csa_tree_add_51_79_groupi_g41463(csa_tree_add_51_79_groupi_n_4656 ,csa_tree_add_51_79_groupi_n_2160 ,csa_tree_add_51_79_groupi_n_420);
  or csa_tree_add_51_79_groupi_g41464(csa_tree_add_51_79_groupi_n_4655 ,csa_tree_add_51_79_groupi_n_2872 ,csa_tree_add_51_79_groupi_n_462);
  or csa_tree_add_51_79_groupi_g41465(csa_tree_add_51_79_groupi_n_4654 ,csa_tree_add_51_79_groupi_n_2871 ,csa_tree_add_51_79_groupi_n_1056);
  or csa_tree_add_51_79_groupi_g41466(csa_tree_add_51_79_groupi_n_4653 ,csa_tree_add_51_79_groupi_n_2868 ,csa_tree_add_51_79_groupi_n_993);
  or csa_tree_add_51_79_groupi_g41467(csa_tree_add_51_79_groupi_n_4652 ,csa_tree_add_51_79_groupi_n_2035 ,csa_tree_add_51_79_groupi_n_900);
  or csa_tree_add_51_79_groupi_g41468(csa_tree_add_51_79_groupi_n_4651 ,csa_tree_add_51_79_groupi_n_2020 ,csa_tree_add_51_79_groupi_n_999);
  or csa_tree_add_51_79_groupi_g41469(csa_tree_add_51_79_groupi_n_4650 ,csa_tree_add_51_79_groupi_n_2867 ,csa_tree_add_51_79_groupi_n_434);
  or csa_tree_add_51_79_groupi_g41470(csa_tree_add_51_79_groupi_n_4649 ,csa_tree_add_51_79_groupi_n_2103 ,csa_tree_add_51_79_groupi_n_990);
  or csa_tree_add_51_79_groupi_g41471(csa_tree_add_51_79_groupi_n_4648 ,csa_tree_add_51_79_groupi_n_2690 ,csa_tree_add_51_79_groupi_n_460);
  or csa_tree_add_51_79_groupi_g41472(csa_tree_add_51_79_groupi_n_4647 ,csa_tree_add_51_79_groupi_n_2647 ,csa_tree_add_51_79_groupi_n_891);
  or csa_tree_add_51_79_groupi_g41473(csa_tree_add_51_79_groupi_n_4646 ,csa_tree_add_51_79_groupi_n_2161 ,csa_tree_add_51_79_groupi_n_420);
  or csa_tree_add_51_79_groupi_g41474(csa_tree_add_51_79_groupi_n_4645 ,csa_tree_add_51_79_groupi_n_2022 ,csa_tree_add_51_79_groupi_n_514);
  and csa_tree_add_51_79_groupi_g41475(csa_tree_add_51_79_groupi_n_4644 ,csa_tree_add_51_79_groupi_n_3261 ,csa_tree_add_51_79_groupi_n_3195);
  nor csa_tree_add_51_79_groupi_g41476(csa_tree_add_51_79_groupi_n_4643 ,csa_tree_add_51_79_groupi_n_2229 ,csa_tree_add_51_79_groupi_n_1068);
  or csa_tree_add_51_79_groupi_g41477(csa_tree_add_51_79_groupi_n_4642 ,csa_tree_add_51_79_groupi_n_2325 ,csa_tree_add_51_79_groupi_n_903);
  or csa_tree_add_51_79_groupi_g41478(csa_tree_add_51_79_groupi_n_4641 ,csa_tree_add_51_79_groupi_n_2267 ,csa_tree_add_51_79_groupi_n_444);
  and csa_tree_add_51_79_groupi_g41479(csa_tree_add_51_79_groupi_n_4640 ,csa_tree_add_51_79_groupi_n_3739 ,csa_tree_add_51_79_groupi_n_3787);
  or csa_tree_add_51_79_groupi_g41480(csa_tree_add_51_79_groupi_n_4639 ,csa_tree_add_51_79_groupi_n_2652 ,csa_tree_add_51_79_groupi_n_452);
  or csa_tree_add_51_79_groupi_g41481(csa_tree_add_51_79_groupi_n_4638 ,csa_tree_add_51_79_groupi_n_2857 ,csa_tree_add_51_79_groupi_n_1062);
  or csa_tree_add_51_79_groupi_g41482(csa_tree_add_51_79_groupi_n_4637 ,csa_tree_add_51_79_groupi_n_2790 ,csa_tree_add_51_79_groupi_n_482);
  or csa_tree_add_51_79_groupi_g41483(csa_tree_add_51_79_groupi_n_4636 ,csa_tree_add_51_79_groupi_n_2854 ,csa_tree_add_51_79_groupi_n_972);
  or csa_tree_add_51_79_groupi_g41484(csa_tree_add_51_79_groupi_n_4635 ,csa_tree_add_51_79_groupi_n_3739 ,csa_tree_add_51_79_groupi_n_3787);
  or csa_tree_add_51_79_groupi_g41485(csa_tree_add_51_79_groupi_n_4634 ,csa_tree_add_51_79_groupi_n_2812 ,csa_tree_add_51_79_groupi_n_492);
  or csa_tree_add_51_79_groupi_g41486(csa_tree_add_51_79_groupi_n_4633 ,csa_tree_add_51_79_groupi_n_3220 ,csa_tree_add_51_79_groupi_n_3258);
  or csa_tree_add_51_79_groupi_g41487(csa_tree_add_51_79_groupi_n_4632 ,csa_tree_add_51_79_groupi_n_2188 ,csa_tree_add_51_79_groupi_n_412);
  or csa_tree_add_51_79_groupi_g41488(csa_tree_add_51_79_groupi_n_4631 ,csa_tree_add_51_79_groupi_n_2048 ,csa_tree_add_51_79_groupi_n_496);
  or csa_tree_add_51_79_groupi_g41489(csa_tree_add_51_79_groupi_n_4630 ,csa_tree_add_51_79_groupi_n_2846 ,csa_tree_add_51_79_groupi_n_1050);
  or csa_tree_add_51_79_groupi_g41490(csa_tree_add_51_79_groupi_n_4629 ,csa_tree_add_51_79_groupi_n_2848 ,csa_tree_add_51_79_groupi_n_918);
  or csa_tree_add_51_79_groupi_g41491(csa_tree_add_51_79_groupi_n_4628 ,csa_tree_add_51_79_groupi_n_2845 ,csa_tree_add_51_79_groupi_n_951);
  or csa_tree_add_51_79_groupi_g41492(csa_tree_add_51_79_groupi_n_4627 ,csa_tree_add_51_79_groupi_n_2773 ,csa_tree_add_51_79_groupi_n_428);
  or csa_tree_add_51_79_groupi_g41493(csa_tree_add_51_79_groupi_n_4626 ,csa_tree_add_51_79_groupi_n_2246 ,csa_tree_add_51_79_groupi_n_897);
  or csa_tree_add_51_79_groupi_g41494(csa_tree_add_51_79_groupi_n_4625 ,csa_tree_add_51_79_groupi_n_2844 ,csa_tree_add_51_79_groupi_n_468);
  or csa_tree_add_51_79_groupi_g41495(csa_tree_add_51_79_groupi_n_4624 ,csa_tree_add_51_79_groupi_n_2236 ,csa_tree_add_51_79_groupi_n_939);
  or csa_tree_add_51_79_groupi_g41496(csa_tree_add_51_79_groupi_n_4623 ,csa_tree_add_51_79_groupi_n_2842 ,csa_tree_add_51_79_groupi_n_912);
  or csa_tree_add_51_79_groupi_g41497(csa_tree_add_51_79_groupi_n_4622 ,csa_tree_add_51_79_groupi_n_2768 ,csa_tree_add_51_79_groupi_n_1014);
  or csa_tree_add_51_79_groupi_g41498(csa_tree_add_51_79_groupi_n_4621 ,csa_tree_add_51_79_groupi_n_2039 ,csa_tree_add_51_79_groupi_n_1002);
  or csa_tree_add_51_79_groupi_g41499(csa_tree_add_51_79_groupi_n_4620 ,csa_tree_add_51_79_groupi_n_2617 ,csa_tree_add_51_79_groupi_n_478);
  or csa_tree_add_51_79_groupi_g41500(csa_tree_add_51_79_groupi_n_4619 ,csa_tree_add_51_79_groupi_n_2312 ,csa_tree_add_51_79_groupi_n_906);
  or csa_tree_add_51_79_groupi_g41501(csa_tree_add_51_79_groupi_n_4618 ,csa_tree_add_51_79_groupi_n_2840 ,csa_tree_add_51_79_groupi_n_1047);
  or csa_tree_add_51_79_groupi_g41502(csa_tree_add_51_79_groupi_n_4617 ,csa_tree_add_51_79_groupi_n_3225 ,csa_tree_add_51_79_groupi_n_3253);
  or csa_tree_add_51_79_groupi_g41503(csa_tree_add_51_79_groupi_n_4616 ,csa_tree_add_51_79_groupi_n_2839 ,csa_tree_add_51_79_groupi_n_436);
  or csa_tree_add_51_79_groupi_g41504(csa_tree_add_51_79_groupi_n_4615 ,csa_tree_add_51_79_groupi_n_2056 ,csa_tree_add_51_79_groupi_n_466);
  or csa_tree_add_51_79_groupi_g41505(csa_tree_add_51_79_groupi_n_4614 ,csa_tree_add_51_79_groupi_n_2837 ,csa_tree_add_51_79_groupi_n_428);
  or csa_tree_add_51_79_groupi_g41506(csa_tree_add_51_79_groupi_n_4613 ,csa_tree_add_51_79_groupi_n_2683 ,csa_tree_add_51_79_groupi_n_936);
  or csa_tree_add_51_79_groupi_g41507(csa_tree_add_51_79_groupi_n_4612 ,csa_tree_add_51_79_groupi_n_2833 ,csa_tree_add_51_79_groupi_n_984);
  nor csa_tree_add_51_79_groupi_g41508(csa_tree_add_51_79_groupi_n_4611 ,csa_tree_add_51_79_groupi_n_2167 ,csa_tree_add_51_79_groupi_n_1053);
  and csa_tree_add_51_79_groupi_g41509(csa_tree_add_51_79_groupi_n_4610 ,csa_tree_add_51_79_groupi_n_3800 ,csa_tree_add_51_79_groupi_n_3801);
  or csa_tree_add_51_79_groupi_g41510(csa_tree_add_51_79_groupi_n_4609 ,csa_tree_add_51_79_groupi_n_2073 ,csa_tree_add_51_79_groupi_n_927);
  or csa_tree_add_51_79_groupi_g41511(csa_tree_add_51_79_groupi_n_4608 ,csa_tree_add_51_79_groupi_n_2069 ,csa_tree_add_51_79_groupi_n_494);
  or csa_tree_add_51_79_groupi_g41512(csa_tree_add_51_79_groupi_n_4607 ,csa_tree_add_51_79_groupi_n_2055 ,csa_tree_add_51_79_groupi_n_954);
  or csa_tree_add_51_79_groupi_g41513(csa_tree_add_51_79_groupi_n_4606 ,csa_tree_add_51_79_groupi_n_2346 ,csa_tree_add_51_79_groupi_n_502);
  or csa_tree_add_51_79_groupi_g41514(csa_tree_add_51_79_groupi_n_4605 ,csa_tree_add_51_79_groupi_n_2828 ,csa_tree_add_51_79_groupi_n_987);
  or csa_tree_add_51_79_groupi_g41515(csa_tree_add_51_79_groupi_n_4604 ,csa_tree_add_51_79_groupi_n_2190 ,csa_tree_add_51_79_groupi_n_1005);
  or csa_tree_add_51_79_groupi_g41516(csa_tree_add_51_79_groupi_n_4603 ,csa_tree_add_51_79_groupi_n_3800 ,csa_tree_add_51_79_groupi_n_3801);
  or csa_tree_add_51_79_groupi_g41517(csa_tree_add_51_79_groupi_n_4602 ,csa_tree_add_51_79_groupi_n_2038 ,csa_tree_add_51_79_groupi_n_945);
  or csa_tree_add_51_79_groupi_g41518(csa_tree_add_51_79_groupi_n_4601 ,csa_tree_add_51_79_groupi_n_2094 ,csa_tree_add_51_79_groupi_n_993);
  or csa_tree_add_51_79_groupi_g41519(csa_tree_add_51_79_groupi_n_4600 ,csa_tree_add_51_79_groupi_n_2753 ,csa_tree_add_51_79_groupi_n_406);
  or csa_tree_add_51_79_groupi_g41520(csa_tree_add_51_79_groupi_n_4599 ,csa_tree_add_51_79_groupi_n_2576 ,csa_tree_add_51_79_groupi_n_484);
  or csa_tree_add_51_79_groupi_g41521(csa_tree_add_51_79_groupi_n_4598 ,csa_tree_add_51_79_groupi_n_2863 ,csa_tree_add_51_79_groupi_n_954);
  or csa_tree_add_51_79_groupi_g41522(csa_tree_add_51_79_groupi_n_4597 ,csa_tree_add_51_79_groupi_n_2824 ,csa_tree_add_51_79_groupi_n_508);
  or csa_tree_add_51_79_groupi_g41523(csa_tree_add_51_79_groupi_n_4596 ,csa_tree_add_51_79_groupi_n_2607 ,csa_tree_add_51_79_groupi_n_450);
  or csa_tree_add_51_79_groupi_g41524(csa_tree_add_51_79_groupi_n_4595 ,csa_tree_add_51_79_groupi_n_2586 ,csa_tree_add_51_79_groupi_n_470);
  or csa_tree_add_51_79_groupi_g41525(csa_tree_add_51_79_groupi_n_4594 ,csa_tree_add_51_79_groupi_n_2593 ,csa_tree_add_51_79_groupi_n_957);
  or csa_tree_add_51_79_groupi_g41526(csa_tree_add_51_79_groupi_n_4593 ,csa_tree_add_51_79_groupi_n_2337 ,csa_tree_add_51_79_groupi_n_900);
  or csa_tree_add_51_79_groupi_g41527(csa_tree_add_51_79_groupi_n_4592 ,csa_tree_add_51_79_groupi_n_2298 ,csa_tree_add_51_79_groupi_n_486);
  or csa_tree_add_51_79_groupi_g41528(csa_tree_add_51_79_groupi_n_4591 ,csa_tree_add_51_79_groupi_n_2819 ,csa_tree_add_51_79_groupi_n_432);
  or csa_tree_add_51_79_groupi_g41529(csa_tree_add_51_79_groupi_n_4590 ,csa_tree_add_51_79_groupi_n_2651 ,csa_tree_add_51_79_groupi_n_915);
  or csa_tree_add_51_79_groupi_g41530(csa_tree_add_51_79_groupi_n_4589 ,csa_tree_add_51_79_groupi_n_2660 ,csa_tree_add_51_79_groupi_n_963);
  or csa_tree_add_51_79_groupi_g41531(csa_tree_add_51_79_groupi_n_4588 ,csa_tree_add_51_79_groupi_n_2664 ,csa_tree_add_51_79_groupi_n_903);
  or csa_tree_add_51_79_groupi_g41532(csa_tree_add_51_79_groupi_n_4587 ,csa_tree_add_51_79_groupi_n_2181 ,csa_tree_add_51_79_groupi_n_418);
  or csa_tree_add_51_79_groupi_g41533(csa_tree_add_51_79_groupi_n_4586 ,csa_tree_add_51_79_groupi_n_2573 ,csa_tree_add_51_79_groupi_n_384);
  or csa_tree_add_51_79_groupi_g41534(csa_tree_add_51_79_groupi_n_4585 ,csa_tree_add_51_79_groupi_n_2816 ,csa_tree_add_51_79_groupi_n_414);
  or csa_tree_add_51_79_groupi_g41535(csa_tree_add_51_79_groupi_n_4584 ,csa_tree_add_51_79_groupi_n_1953 ,csa_tree_add_51_79_groupi_n_518);
  or csa_tree_add_51_79_groupi_g41536(csa_tree_add_51_79_groupi_n_4583 ,csa_tree_add_51_79_groupi_n_2762 ,csa_tree_add_51_79_groupi_n_472);
  or csa_tree_add_51_79_groupi_g41537(csa_tree_add_51_79_groupi_n_4582 ,csa_tree_add_51_79_groupi_n_2284 ,csa_tree_add_51_79_groupi_n_464);
  or csa_tree_add_51_79_groupi_g41538(csa_tree_add_51_79_groupi_n_4581 ,csa_tree_add_51_79_groupi_n_2725 ,csa_tree_add_51_79_groupi_n_48);
  or csa_tree_add_51_79_groupi_g41539(csa_tree_add_51_79_groupi_n_4580 ,csa_tree_add_51_79_groupi_n_2720 ,csa_tree_add_51_79_groupi_n_500);
  nor csa_tree_add_51_79_groupi_g41540(csa_tree_add_51_79_groupi_n_4579 ,csa_tree_add_51_79_groupi_n_2175 ,csa_tree_add_51_79_groupi_n_1041);
  or csa_tree_add_51_79_groupi_g41541(csa_tree_add_51_79_groupi_n_4578 ,csa_tree_add_51_79_groupi_n_2861 ,csa_tree_add_51_79_groupi_n_1026);
  or csa_tree_add_51_79_groupi_g41542(csa_tree_add_51_79_groupi_n_4577 ,csa_tree_add_51_79_groupi_n_2813 ,csa_tree_add_51_79_groupi_n_948);
  and csa_tree_add_51_79_groupi_g41543(csa_tree_add_51_79_groupi_n_4576 ,csa_tree_add_51_79_groupi_n_1071 ,csa_tree_add_51_79_groupi_n_3282);
  or csa_tree_add_51_79_groupi_g41544(csa_tree_add_51_79_groupi_n_4575 ,csa_tree_add_51_79_groupi_n_2746 ,csa_tree_add_51_79_groupi_n_520);
  or csa_tree_add_51_79_groupi_g41545(csa_tree_add_51_79_groupi_n_4574 ,csa_tree_add_51_79_groupi_n_2259 ,csa_tree_add_51_79_groupi_n_108);
  nor csa_tree_add_51_79_groupi_g41546(csa_tree_add_51_79_groupi_n_4573 ,csa_tree_add_51_79_groupi_n_3797 ,csa_tree_add_51_79_groupi_n_3815);
  or csa_tree_add_51_79_groupi_g41547(csa_tree_add_51_79_groupi_n_4572 ,csa_tree_add_51_79_groupi_n_2693 ,csa_tree_add_51_79_groupi_n_930);
  or csa_tree_add_51_79_groupi_g41548(csa_tree_add_51_79_groupi_n_4571 ,csa_tree_add_51_79_groupi_n_2253 ,csa_tree_add_51_79_groupi_n_1032);
  or csa_tree_add_51_79_groupi_g41549(csa_tree_add_51_79_groupi_n_4570 ,csa_tree_add_51_79_groupi_n_2571 ,csa_tree_add_51_79_groupi_n_2916);
  or csa_tree_add_51_79_groupi_g41550(csa_tree_add_51_79_groupi_n_4569 ,csa_tree_add_51_79_groupi_n_2124 ,csa_tree_add_51_79_groupi_n_246);
  or csa_tree_add_51_79_groupi_g41551(csa_tree_add_51_79_groupi_n_4568 ,csa_tree_add_51_79_groupi_n_2277 ,csa_tree_add_51_79_groupi_n_930);
  or csa_tree_add_51_79_groupi_g41552(csa_tree_add_51_79_groupi_n_4567 ,csa_tree_add_51_79_groupi_n_2237 ,csa_tree_add_51_79_groupi_n_156);
  or csa_tree_add_51_79_groupi_g41553(csa_tree_add_51_79_groupi_n_4566 ,csa_tree_add_51_79_groupi_n_2719 ,csa_tree_add_51_79_groupi_n_432);
  or csa_tree_add_51_79_groupi_g41554(csa_tree_add_51_79_groupi_n_4565 ,csa_tree_add_51_79_groupi_n_2168 ,csa_tree_add_51_79_groupi_n_894);
  or csa_tree_add_51_79_groupi_g41555(csa_tree_add_51_79_groupi_n_4564 ,csa_tree_add_51_79_groupi_n_2158 ,csa_tree_add_51_79_groupi_n_1032);
  or csa_tree_add_51_79_groupi_g41556(csa_tree_add_51_79_groupi_n_4563 ,csa_tree_add_51_79_groupi_n_2851 ,csa_tree_add_51_79_groupi_n_945);
  or csa_tree_add_51_79_groupi_g41557(csa_tree_add_51_79_groupi_n_4562 ,csa_tree_add_51_79_groupi_n_2856 ,csa_tree_add_51_79_groupi_n_963);
  nor csa_tree_add_51_79_groupi_g41558(csa_tree_add_51_79_groupi_n_4561 ,csa_tree_add_51_79_groupi_n_2655 ,csa_tree_add_51_79_groupi_n_1047);
  or csa_tree_add_51_79_groupi_g41559(csa_tree_add_51_79_groupi_n_4560 ,csa_tree_add_51_79_groupi_n_2245 ,csa_tree_add_51_79_groupi_n_442);
  or csa_tree_add_51_79_groupi_g41560(csa_tree_add_51_79_groupi_n_4559 ,csa_tree_add_51_79_groupi_n_2796 ,csa_tree_add_51_79_groupi_n_963);
  or csa_tree_add_51_79_groupi_g41561(csa_tree_add_51_79_groupi_n_4558 ,csa_tree_add_51_79_groupi_n_2591 ,csa_tree_add_51_79_groupi_n_198);
  or csa_tree_add_51_79_groupi_g41562(csa_tree_add_51_79_groupi_n_4557 ,csa_tree_add_51_79_groupi_n_2176 ,csa_tree_add_51_79_groupi_n_1041);
  or csa_tree_add_51_79_groupi_g41563(csa_tree_add_51_79_groupi_n_4556 ,csa_tree_add_51_79_groupi_n_2182 ,csa_tree_add_51_79_groupi_n_1008);
  or csa_tree_add_51_79_groupi_g41564(csa_tree_add_51_79_groupi_n_4555 ,csa_tree_add_51_79_groupi_n_2822 ,csa_tree_add_51_79_groupi_n_921);
  and csa_tree_add_51_79_groupi_g41565(csa_tree_add_51_79_groupi_n_4554 ,csa_tree_add_51_79_groupi_n_3795 ,csa_tree_add_51_79_groupi_n_3216);
  or csa_tree_add_51_79_groupi_g41566(csa_tree_add_51_79_groupi_n_4553 ,csa_tree_add_51_79_groupi_n_2820 ,csa_tree_add_51_79_groupi_n_948);
  or csa_tree_add_51_79_groupi_g41567(csa_tree_add_51_79_groupi_n_4552 ,csa_tree_add_51_79_groupi_n_2310 ,csa_tree_add_51_79_groupi_n_506);
  or csa_tree_add_51_79_groupi_g41568(csa_tree_add_51_79_groupi_n_4551 ,csa_tree_add_51_79_groupi_n_2070 ,csa_tree_add_51_79_groupi_n_996);
  and csa_tree_add_51_79_groupi_g41569(csa_tree_add_51_79_groupi_n_4550 ,csa_tree_add_51_79_groupi_n_3738 ,csa_tree_add_51_79_groupi_n_3242);
  or csa_tree_add_51_79_groupi_g41570(csa_tree_add_51_79_groupi_n_4549 ,csa_tree_add_51_79_groupi_n_3266 ,csa_tree_add_51_79_groupi_n_3263);
  or csa_tree_add_51_79_groupi_g41571(csa_tree_add_51_79_groupi_n_4548 ,csa_tree_add_51_79_groupi_n_2196 ,csa_tree_add_51_79_groupi_n_253);
  or csa_tree_add_51_79_groupi_g41572(csa_tree_add_51_79_groupi_n_4547 ,csa_tree_add_51_79_groupi_n_2242 ,csa_tree_add_51_79_groupi_n_408);
  or csa_tree_add_51_79_groupi_g41573(csa_tree_add_51_79_groupi_n_4546 ,csa_tree_add_51_79_groupi_n_2122 ,csa_tree_add_51_79_groupi_n_1068);
  or csa_tree_add_51_79_groupi_g41574(csa_tree_add_51_79_groupi_n_4545 ,csa_tree_add_51_79_groupi_n_2194 ,csa_tree_add_51_79_groupi_n_1059);
  or csa_tree_add_51_79_groupi_g41575(csa_tree_add_51_79_groupi_n_4544 ,csa_tree_add_51_79_groupi_n_2771 ,csa_tree_add_51_79_groupi_n_924);
  or csa_tree_add_51_79_groupi_g41576(csa_tree_add_51_79_groupi_n_4543 ,csa_tree_add_51_79_groupi_n_2061 ,csa_tree_add_51_79_groupi_n_936);
  or csa_tree_add_51_79_groupi_g41577(csa_tree_add_51_79_groupi_n_4542 ,csa_tree_add_51_79_groupi_n_2026 ,csa_tree_add_51_79_groupi_n_978);
  or csa_tree_add_51_79_groupi_g41578(csa_tree_add_51_79_groupi_n_4541 ,csa_tree_add_51_79_groupi_n_2082 ,csa_tree_add_51_79_groupi_n_975);
  or csa_tree_add_51_79_groupi_g41579(csa_tree_add_51_79_groupi_n_4540 ,csa_tree_add_51_79_groupi_n_2769 ,csa_tree_add_51_79_groupi_n_422);
  or csa_tree_add_51_79_groupi_g41580(csa_tree_add_51_79_groupi_n_4539 ,csa_tree_add_51_79_groupi_n_2597 ,csa_tree_add_51_79_groupi_n_996);
  or csa_tree_add_51_79_groupi_g41581(csa_tree_add_51_79_groupi_n_4538 ,csa_tree_add_51_79_groupi_n_2108 ,csa_tree_add_51_79_groupi_n_504);
  or csa_tree_add_51_79_groupi_g41582(csa_tree_add_51_79_groupi_n_4537 ,csa_tree_add_51_79_groupi_n_2150 ,csa_tree_add_51_79_groupi_n_972);
  or csa_tree_add_51_79_groupi_g41583(csa_tree_add_51_79_groupi_n_4536 ,csa_tree_add_51_79_groupi_n_2149 ,csa_tree_add_51_79_groupi_n_488);
  or csa_tree_add_51_79_groupi_g41584(csa_tree_add_51_79_groupi_n_4535 ,csa_tree_add_51_79_groupi_n_2767 ,csa_tree_add_51_79_groupi_n_933);
  or csa_tree_add_51_79_groupi_g41585(csa_tree_add_51_79_groupi_n_4534 ,csa_tree_add_51_79_groupi_n_3738 ,csa_tree_add_51_79_groupi_n_3242);
  or csa_tree_add_51_79_groupi_g41586(csa_tree_add_51_79_groupi_n_4533 ,csa_tree_add_51_79_groupi_n_2766 ,csa_tree_add_51_79_groupi_n_456);
  or csa_tree_add_51_79_groupi_g41587(csa_tree_add_51_79_groupi_n_4532 ,csa_tree_add_51_79_groupi_n_2019 ,csa_tree_add_51_79_groupi_n_912);
  or csa_tree_add_51_79_groupi_g41588(csa_tree_add_51_79_groupi_n_4531 ,csa_tree_add_51_79_groupi_n_2765 ,csa_tree_add_51_79_groupi_n_438);
  or csa_tree_add_51_79_groupi_g41589(csa_tree_add_51_79_groupi_n_4530 ,csa_tree_add_51_79_groupi_n_2764 ,csa_tree_add_51_79_groupi_n_975);
  or csa_tree_add_51_79_groupi_g41590(csa_tree_add_51_79_groupi_n_4529 ,csa_tree_add_51_79_groupi_n_2269 ,csa_tree_add_51_79_groupi_n_897);
  or csa_tree_add_51_79_groupi_g41591(csa_tree_add_51_79_groupi_n_4528 ,csa_tree_add_51_79_groupi_n_2066 ,csa_tree_add_51_79_groupi_n_430);
  or csa_tree_add_51_79_groupi_g41592(csa_tree_add_51_79_groupi_n_4527 ,csa_tree_add_51_79_groupi_n_2761 ,csa_tree_add_51_79_groupi_n_102);
  or csa_tree_add_51_79_groupi_g41593(csa_tree_add_51_79_groupi_n_4526 ,csa_tree_add_51_79_groupi_n_1899 ,csa_tree_add_51_79_groupi_n_472);
  or csa_tree_add_51_79_groupi_g41594(csa_tree_add_51_79_groupi_n_4525 ,csa_tree_add_51_79_groupi_n_2080 ,csa_tree_add_51_79_groupi_n_512);
  or csa_tree_add_51_79_groupi_g41595(csa_tree_add_51_79_groupi_n_4524 ,csa_tree_add_51_79_groupi_n_2036 ,csa_tree_add_51_79_groupi_n_903);
  or csa_tree_add_51_79_groupi_g41596(csa_tree_add_51_79_groupi_n_4523 ,csa_tree_add_51_79_groupi_n_2704 ,csa_tree_add_51_79_groupi_n_454);
  or csa_tree_add_51_79_groupi_g41597(csa_tree_add_51_79_groupi_n_4522 ,csa_tree_add_51_79_groupi_n_1933 ,csa_tree_add_51_79_groupi_n_414);
  or csa_tree_add_51_79_groupi_g41598(csa_tree_add_51_79_groupi_n_4521 ,csa_tree_add_51_79_groupi_n_2575 ,csa_tree_add_51_79_groupi_n_1014);
  or csa_tree_add_51_79_groupi_g41599(csa_tree_add_51_79_groupi_n_4520 ,csa_tree_add_51_79_groupi_n_2216 ,csa_tree_add_51_79_groupi_n_440);
  or csa_tree_add_51_79_groupi_g41600(csa_tree_add_51_79_groupi_n_4519 ,csa_tree_add_51_79_groupi_n_2758 ,csa_tree_add_51_79_groupi_n_927);
  or csa_tree_add_51_79_groupi_g41601(csa_tree_add_51_79_groupi_n_4518 ,csa_tree_add_51_79_groupi_n_2348 ,csa_tree_add_51_79_groupi_n_494);
  or csa_tree_add_51_79_groupi_g41602(csa_tree_add_51_79_groupi_n_4517 ,csa_tree_add_51_79_groupi_n_2711 ,csa_tree_add_51_79_groupi_n_464);
  or csa_tree_add_51_79_groupi_g41603(csa_tree_add_51_79_groupi_n_4516 ,csa_tree_add_51_79_groupi_n_2358 ,csa_tree_add_51_79_groupi_n_478);
  or csa_tree_add_51_79_groupi_g41604(csa_tree_add_51_79_groupi_n_4515 ,csa_tree_add_51_79_groupi_n_2232 ,csa_tree_add_51_79_groupi_n_1011);
  or csa_tree_add_51_79_groupi_g41605(csa_tree_add_51_79_groupi_n_4514 ,csa_tree_add_51_79_groupi_n_2353 ,csa_tree_add_51_79_groupi_n_972);
  or csa_tree_add_51_79_groupi_g41606(csa_tree_add_51_79_groupi_n_4513 ,csa_tree_add_51_79_groupi_n_2046 ,csa_tree_add_51_79_groupi_n_921);
  or csa_tree_add_51_79_groupi_g41607(csa_tree_add_51_79_groupi_n_4512 ,csa_tree_add_51_79_groupi_n_2754 ,csa_tree_add_51_79_groupi_n_969);
  or csa_tree_add_51_79_groupi_g41608(csa_tree_add_51_79_groupi_n_4511 ,csa_tree_add_51_79_groupi_n_2755 ,csa_tree_add_51_79_groupi_n_1029);
  or csa_tree_add_51_79_groupi_g41609(csa_tree_add_51_79_groupi_n_4510 ,csa_tree_add_51_79_groupi_n_2752 ,csa_tree_add_51_79_groupi_n_66);
  or csa_tree_add_51_79_groupi_g41610(csa_tree_add_51_79_groupi_n_4509 ,csa_tree_add_51_79_groupi_n_1908 ,csa_tree_add_51_79_groupi_n_448);
  or csa_tree_add_51_79_groupi_g41611(csa_tree_add_51_79_groupi_n_4508 ,csa_tree_add_51_79_groupi_n_2623 ,csa_tree_add_51_79_groupi_n_466);
  or csa_tree_add_51_79_groupi_g41612(csa_tree_add_51_79_groupi_n_4507 ,csa_tree_add_51_79_groupi_n_2626 ,csa_tree_add_51_79_groupi_n_990);
  or csa_tree_add_51_79_groupi_g41613(csa_tree_add_51_79_groupi_n_4506 ,csa_tree_add_51_79_groupi_n_2750 ,csa_tree_add_51_79_groupi_n_981);
  or csa_tree_add_51_79_groupi_g41614(csa_tree_add_51_79_groupi_n_4505 ,csa_tree_add_51_79_groupi_n_2731 ,csa_tree_add_51_79_groupi_n_60);
  or csa_tree_add_51_79_groupi_g41615(csa_tree_add_51_79_groupi_n_4504 ,csa_tree_add_51_79_groupi_n_2748 ,csa_tree_add_51_79_groupi_n_894);
  or csa_tree_add_51_79_groupi_g41616(csa_tree_add_51_79_groupi_n_4503 ,csa_tree_add_51_79_groupi_n_2601 ,csa_tree_add_51_79_groupi_n_945);
  or csa_tree_add_51_79_groupi_g41617(csa_tree_add_51_79_groupi_n_4502 ,csa_tree_add_51_79_groupi_n_3795 ,csa_tree_add_51_79_groupi_n_3216);
  or csa_tree_add_51_79_groupi_g41618(csa_tree_add_51_79_groupi_n_4501 ,csa_tree_add_51_79_groupi_n_2662 ,csa_tree_add_51_79_groupi_n_480);
  or csa_tree_add_51_79_groupi_g41619(csa_tree_add_51_79_groupi_n_4500 ,csa_tree_add_51_79_groupi_n_2350 ,csa_tree_add_51_79_groupi_n_969);
  or csa_tree_add_51_79_groupi_g41620(csa_tree_add_51_79_groupi_n_4499 ,csa_tree_add_51_79_groupi_n_2708 ,csa_tree_add_51_79_groupi_n_1014);
  or csa_tree_add_51_79_groupi_g41621(csa_tree_add_51_79_groupi_n_4498 ,csa_tree_add_51_79_groupi_n_2742 ,csa_tree_add_51_79_groupi_n_966);
  or csa_tree_add_51_79_groupi_g41622(csa_tree_add_51_79_groupi_n_4497 ,csa_tree_add_51_79_groupi_n_2741 ,csa_tree_add_51_79_groupi_n_410);
  or csa_tree_add_51_79_groupi_g41623(csa_tree_add_51_79_groupi_n_4496 ,csa_tree_add_51_79_groupi_n_2359 ,csa_tree_add_51_79_groupi_n_1002);
  or csa_tree_add_51_79_groupi_g41624(csa_tree_add_51_79_groupi_n_4495 ,csa_tree_add_51_79_groupi_n_2705 ,csa_tree_add_51_79_groupi_n_978);
  or csa_tree_add_51_79_groupi_g41625(csa_tree_add_51_79_groupi_n_4494 ,csa_tree_add_51_79_groupi_n_2710 ,csa_tree_add_51_79_groupi_n_150);
  or csa_tree_add_51_79_groupi_g41626(csa_tree_add_51_79_groupi_n_4493 ,csa_tree_add_51_79_groupi_n_2734 ,csa_tree_add_51_79_groupi_n_909);
  or csa_tree_add_51_79_groupi_g41627(csa_tree_add_51_79_groupi_n_4492 ,csa_tree_add_51_79_groupi_n_2370 ,csa_tree_add_51_79_groupi_n_966);
  or csa_tree_add_51_79_groupi_g41628(csa_tree_add_51_79_groupi_n_4491 ,csa_tree_add_51_79_groupi_n_2786 ,csa_tree_add_51_79_groupi_n_476);
  and csa_tree_add_51_79_groupi_g41629(csa_tree_add_51_79_groupi_n_4490 ,csa_tree_add_51_79_groupi_n_3797 ,csa_tree_add_51_79_groupi_n_3815);
  or csa_tree_add_51_79_groupi_g41630(csa_tree_add_51_79_groupi_n_4489 ,csa_tree_add_51_79_groupi_n_2770 ,csa_tree_add_51_79_groupi_n_981);
  or csa_tree_add_51_79_groupi_g41631(csa_tree_add_51_79_groupi_n_4488 ,csa_tree_add_51_79_groupi_n_2724 ,csa_tree_add_51_79_groupi_n_458);
  or csa_tree_add_51_79_groupi_g41632(csa_tree_add_51_79_groupi_n_4487 ,csa_tree_add_51_79_groupi_n_2800 ,csa_tree_add_51_79_groupi_n_891);
  or csa_tree_add_51_79_groupi_g41633(csa_tree_add_51_79_groupi_n_4486 ,csa_tree_add_51_79_groupi_n_2808 ,csa_tree_add_51_79_groupi_n_474);
  or csa_tree_add_51_79_groupi_g41634(csa_tree_add_51_79_groupi_n_4485 ,csa_tree_add_51_79_groupi_n_2735 ,csa_tree_add_51_79_groupi_n_484);
  or csa_tree_add_51_79_groupi_g41635(csa_tree_add_51_79_groupi_n_4484 ,csa_tree_add_51_79_groupi_n_2335 ,csa_tree_add_51_79_groupi_n_993);
  or csa_tree_add_51_79_groupi_g41636(csa_tree_add_51_79_groupi_n_4483 ,csa_tree_add_51_79_groupi_n_3217 ,csa_tree_add_51_79_groupi_n_3218);
  and csa_tree_add_51_79_groupi_g41637(csa_tree_add_51_79_groupi_n_4482 ,csa_tree_add_51_79_groupi_n_3217 ,csa_tree_add_51_79_groupi_n_3218);
  nor csa_tree_add_51_79_groupi_g41638(csa_tree_add_51_79_groupi_n_4481 ,csa_tree_add_51_79_groupi_n_2118 ,csa_tree_add_51_79_groupi_n_1050);
  or csa_tree_add_51_79_groupi_g41639(csa_tree_add_51_79_groupi_n_4480 ,csa_tree_add_51_79_groupi_n_2260 ,csa_tree_add_51_79_groupi_n_1011);
  or csa_tree_add_51_79_groupi_g41640(csa_tree_add_51_79_groupi_n_4479 ,csa_tree_add_51_79_groupi_n_2051 ,csa_tree_add_51_79_groupi_n_1029);
  or csa_tree_add_51_79_groupi_g41641(csa_tree_add_51_79_groupi_n_4478 ,csa_tree_add_51_79_groupi_n_3267 ,csa_tree_add_51_79_groupi_n_3221);
  or csa_tree_add_51_79_groupi_g41642(csa_tree_add_51_79_groupi_n_4477 ,csa_tree_add_51_79_groupi_n_2083 ,csa_tree_add_51_79_groupi_n_915);
  or csa_tree_add_51_79_groupi_g41643(csa_tree_add_51_79_groupi_n_4476 ,csa_tree_add_51_79_groupi_n_2164 ,csa_tree_add_51_79_groupi_n_1041);
  or csa_tree_add_51_79_groupi_g41644(csa_tree_add_51_79_groupi_n_4475 ,csa_tree_add_51_79_groupi_n_2079 ,csa_tree_add_51_79_groupi_n_416);
  or csa_tree_add_51_79_groupi_g41645(csa_tree_add_51_79_groupi_n_4474 ,csa_tree_add_51_79_groupi_n_2630 ,csa_tree_add_51_79_groupi_n_510);
  or csa_tree_add_51_79_groupi_g41646(csa_tree_add_51_79_groupi_n_4473 ,csa_tree_add_51_79_groupi_n_2637 ,csa_tree_add_51_79_groupi_n_951);
  or csa_tree_add_51_79_groupi_g41647(csa_tree_add_51_79_groupi_n_4472 ,csa_tree_add_51_79_groupi_n_2722 ,csa_tree_add_51_79_groupi_n_404);
  or csa_tree_add_51_79_groupi_g41648(csa_tree_add_51_79_groupi_n_4471 ,csa_tree_add_51_79_groupi_n_2279 ,csa_tree_add_51_79_groupi_n_990);
  or csa_tree_add_51_79_groupi_g41649(csa_tree_add_51_79_groupi_n_4470 ,csa_tree_add_51_79_groupi_n_2582 ,csa_tree_add_51_79_groupi_n_957);
  or csa_tree_add_51_79_groupi_g41650(csa_tree_add_51_79_groupi_n_4469 ,csa_tree_add_51_79_groupi_n_2251 ,csa_tree_add_51_79_groupi_n_939);
  or csa_tree_add_51_79_groupi_g41651(csa_tree_add_51_79_groupi_n_4468 ,csa_tree_add_51_79_groupi_n_2875 ,csa_tree_add_51_79_groupi_n_900);
  or csa_tree_add_51_79_groupi_g41652(csa_tree_add_51_79_groupi_n_4467 ,csa_tree_add_51_79_groupi_n_2641 ,csa_tree_add_51_79_groupi_n_960);
  or csa_tree_add_51_79_groupi_g41653(csa_tree_add_51_79_groupi_n_4466 ,csa_tree_add_51_79_groupi_n_2054 ,csa_tree_add_51_79_groupi_n_954);
  or csa_tree_add_51_79_groupi_g41654(csa_tree_add_51_79_groupi_n_4465 ,csa_tree_add_51_79_groupi_n_2234 ,csa_tree_add_51_79_groupi_n_516);
  or csa_tree_add_51_79_groupi_g41655(csa_tree_add_51_79_groupi_n_4464 ,csa_tree_add_51_79_groupi_n_2561 ,csa_tree_add_51_79_groupi_n_2990);
  or csa_tree_add_51_79_groupi_g41656(csa_tree_add_51_79_groupi_n_4463 ,csa_tree_add_51_79_groupi_n_2789 ,csa_tree_add_51_79_groupi_n_999);
  or csa_tree_add_51_79_groupi_g41657(csa_tree_add_51_79_groupi_n_4462 ,csa_tree_add_51_79_groupi_n_2214 ,csa_tree_add_51_79_groupi_n_909);
  or csa_tree_add_51_79_groupi_g41658(csa_tree_add_51_79_groupi_n_4461 ,csa_tree_add_51_79_groupi_n_2565 ,csa_tree_add_51_79_groupi_n_2965);
  or csa_tree_add_51_79_groupi_g41659(csa_tree_add_51_79_groupi_n_4460 ,csa_tree_add_51_79_groupi_n_2033 ,csa_tree_add_51_79_groupi_n_229);
  or csa_tree_add_51_79_groupi_g41660(csa_tree_add_51_79_groupi_n_4459 ,csa_tree_add_51_79_groupi_n_2673 ,csa_tree_add_51_79_groupi_n_406);
  or csa_tree_add_51_79_groupi_g41661(csa_tree_add_51_79_groupi_n_4458 ,csa_tree_add_51_79_groupi_n_2566 ,csa_tree_add_51_79_groupi_n_3389);
  or csa_tree_add_51_79_groupi_g41662(csa_tree_add_51_79_groupi_n_4457 ,csa_tree_add_51_79_groupi_n_2680 ,csa_tree_add_51_79_groupi_n_54);
  or csa_tree_add_51_79_groupi_g41663(csa_tree_add_51_79_groupi_n_4456 ,csa_tree_add_51_79_groupi_n_3219 ,csa_tree_add_51_79_groupi_n_3223);
  or csa_tree_add_51_79_groupi_g41664(csa_tree_add_51_79_groupi_n_4455 ,csa_tree_add_51_79_groupi_n_2792 ,csa_tree_add_51_79_groupi_n_446);
  or csa_tree_add_51_79_groupi_g41665(csa_tree_add_51_79_groupi_n_4454 ,csa_tree_add_51_79_groupi_n_2632 ,csa_tree_add_51_79_groupi_n_942);
  or csa_tree_add_51_79_groupi_g41666(csa_tree_add_51_79_groupi_n_4453 ,csa_tree_add_51_79_groupi_n_2225 ,csa_tree_add_51_79_groupi_n_402);
  or csa_tree_add_51_79_groupi_g41667(csa_tree_add_51_79_groupi_n_4452 ,csa_tree_add_51_79_groupi_n_2834 ,csa_tree_add_51_79_groupi_n_984);
  or csa_tree_add_51_79_groupi_g41668(csa_tree_add_51_79_groupi_n_4451 ,csa_tree_add_51_79_groupi_n_2627 ,csa_tree_add_51_79_groupi_n_924);
  or csa_tree_add_51_79_groupi_g41669(csa_tree_add_51_79_groupi_n_4450 ,csa_tree_add_51_79_groupi_n_2714 ,csa_tree_add_51_79_groupi_n_410);
  or csa_tree_add_51_79_groupi_g41670(csa_tree_add_51_79_groupi_n_4449 ,csa_tree_add_51_79_groupi_n_2352 ,csa_tree_add_51_79_groupi_n_1038);
  or csa_tree_add_51_79_groupi_g41671(csa_tree_add_51_79_groupi_n_4448 ,csa_tree_add_51_79_groupi_n_2191 ,csa_tree_add_51_79_groupi_n_1035);
  and csa_tree_add_51_79_groupi_g41672(csa_tree_add_51_79_groupi_n_4447 ,csa_tree_add_51_79_groupi_n_3790 ,csa_tree_add_51_79_groupi_n_3781);
  or csa_tree_add_51_79_groupi_g41673(csa_tree_add_51_79_groupi_n_4446 ,csa_tree_add_51_79_groupi_n_2262 ,csa_tree_add_51_79_groupi_n_1053);
  or csa_tree_add_51_79_groupi_g41674(csa_tree_add_51_79_groupi_n_4445 ,csa_tree_add_51_79_groupi_n_2126 ,csa_tree_add_51_79_groupi_n_918);
  or csa_tree_add_51_79_groupi_g41675(csa_tree_add_51_79_groupi_n_4444 ,csa_tree_add_51_79_groupi_n_2105 ,csa_tree_add_51_79_groupi_n_1050);
  or csa_tree_add_51_79_groupi_g41676(csa_tree_add_51_79_groupi_n_4443 ,csa_tree_add_51_79_groupi_n_2788 ,csa_tree_add_51_79_groupi_n_972);
  or csa_tree_add_51_79_groupi_g41677(csa_tree_add_51_79_groupi_n_4442 ,csa_tree_add_51_79_groupi_n_2029 ,csa_tree_add_51_79_groupi_n_933);
  or csa_tree_add_51_79_groupi_g41678(csa_tree_add_51_79_groupi_n_4441 ,csa_tree_add_51_79_groupi_n_2222 ,csa_tree_add_51_79_groupi_n_157);
  nor csa_tree_add_51_79_groupi_g41679(csa_tree_add_51_79_groupi_n_4440 ,csa_tree_add_51_79_groupi_n_2235 ,csa_tree_add_51_79_groupi_n_1029);
  or csa_tree_add_51_79_groupi_g41680(csa_tree_add_51_79_groupi_n_4439 ,csa_tree_add_51_79_groupi_n_2077 ,csa_tree_add_51_79_groupi_n_906);
  or csa_tree_add_51_79_groupi_g41681(csa_tree_add_51_79_groupi_n_4438 ,csa_tree_add_51_79_groupi_n_2805 ,csa_tree_add_51_79_groupi_n_349);
  or csa_tree_add_51_79_groupi_g41682(csa_tree_add_51_79_groupi_n_4437 ,csa_tree_add_51_79_groupi_n_2220 ,csa_tree_add_51_79_groupi_n_939);
  or csa_tree_add_51_79_groupi_g41683(csa_tree_add_51_79_groupi_n_4436 ,csa_tree_add_51_79_groupi_n_2243 ,csa_tree_add_51_79_groupi_n_1005);
  and csa_tree_add_51_79_groupi_g41684(csa_tree_add_51_79_groupi_n_4435 ,csa_tree_add_51_79_groupi_n_3267 ,csa_tree_add_51_79_groupi_n_3221);
  and csa_tree_add_51_79_groupi_g41685(csa_tree_add_51_79_groupi_n_4434 ,csa_tree_add_51_79_groupi_n_3262 ,csa_tree_add_51_79_groupi_n_3203);
  or csa_tree_add_51_79_groupi_g41686(csa_tree_add_51_79_groupi_n_4433 ,csa_tree_add_51_79_groupi_n_2732 ,csa_tree_add_51_79_groupi_n_1065);
  or csa_tree_add_51_79_groupi_g41687(csa_tree_add_51_79_groupi_n_4432 ,csa_tree_add_51_79_groupi_n_2096 ,csa_tree_add_51_79_groupi_n_434);
  or csa_tree_add_51_79_groupi_g41688(csa_tree_add_51_79_groupi_n_4431 ,csa_tree_add_51_79_groupi_n_2657 ,csa_tree_add_51_79_groupi_n_942);
  or csa_tree_add_51_79_groupi_g41689(csa_tree_add_51_79_groupi_n_4430 ,csa_tree_add_51_79_groupi_n_2642 ,csa_tree_add_51_79_groupi_n_1023);
  or csa_tree_add_51_79_groupi_g41690(csa_tree_add_51_79_groupi_n_4429 ,csa_tree_add_51_79_groupi_n_2676 ,csa_tree_add_51_79_groupi_n_945);
  or csa_tree_add_51_79_groupi_g41691(csa_tree_add_51_79_groupi_n_4428 ,csa_tree_add_51_79_groupi_n_2739 ,csa_tree_add_51_79_groupi_n_987);
  or csa_tree_add_51_79_groupi_g41692(csa_tree_add_51_79_groupi_n_4427 ,csa_tree_add_51_79_groupi_n_2633 ,csa_tree_add_51_79_groupi_n_960);
  or csa_tree_add_51_79_groupi_g41693(csa_tree_add_51_79_groupi_n_4426 ,csa_tree_add_51_79_groupi_n_2847 ,csa_tree_add_51_79_groupi_n_891);
  or csa_tree_add_51_79_groupi_g41694(csa_tree_add_51_79_groupi_n_4425 ,csa_tree_add_51_79_groupi_n_2208 ,csa_tree_add_51_79_groupi_n_1008);
  or csa_tree_add_51_79_groupi_g41695(csa_tree_add_51_79_groupi_n_4424 ,csa_tree_add_51_79_groupi_n_2670 ,csa_tree_add_51_79_groupi_n_460);
  or csa_tree_add_51_79_groupi_g41696(csa_tree_add_51_79_groupi_n_4423 ,csa_tree_add_51_79_groupi_n_2672 ,csa_tree_add_51_79_groupi_n_450);
  or csa_tree_add_51_79_groupi_g41697(csa_tree_add_51_79_groupi_n_4422 ,csa_tree_add_51_79_groupi_n_2803 ,csa_tree_add_51_79_groupi_n_496);
  or csa_tree_add_51_79_groupi_g41698(csa_tree_add_51_79_groupi_n_4421 ,csa_tree_add_51_79_groupi_n_2304 ,csa_tree_add_51_79_groupi_n_343);
  or csa_tree_add_51_79_groupi_g41699(csa_tree_add_51_79_groupi_n_4420 ,csa_tree_add_51_79_groupi_n_2674 ,csa_tree_add_51_79_groupi_n_49);
  or csa_tree_add_51_79_groupi_g41700(csa_tree_add_51_79_groupi_n_4419 ,csa_tree_add_51_79_groupi_n_2628 ,csa_tree_add_51_79_groupi_n_984);
  or csa_tree_add_51_79_groupi_g41701(csa_tree_add_51_79_groupi_n_4418 ,csa_tree_add_51_79_groupi_n_2830 ,csa_tree_add_51_79_groupi_n_490);
  or csa_tree_add_51_79_groupi_g41702(csa_tree_add_51_79_groupi_n_4417 ,csa_tree_add_51_79_groupi_n_2814 ,csa_tree_add_51_79_groupi_n_265);
  or csa_tree_add_51_79_groupi_g41703(csa_tree_add_51_79_groupi_n_4416 ,csa_tree_add_51_79_groupi_n_2285 ,csa_tree_add_51_79_groupi_n_498);
  or csa_tree_add_51_79_groupi_g41704(csa_tree_add_51_79_groupi_n_4415 ,csa_tree_add_51_79_groupi_n_2578 ,csa_tree_add_51_79_groupi_n_508);
  or csa_tree_add_51_79_groupi_g41705(csa_tree_add_51_79_groupi_n_4414 ,csa_tree_add_51_79_groupi_n_2305 ,csa_tree_add_51_79_groupi_n_1038);
  or csa_tree_add_51_79_groupi_g41706(csa_tree_add_51_79_groupi_n_4413 ,csa_tree_add_51_79_groupi_n_2131 ,csa_tree_add_51_79_groupi_n_442);
  or csa_tree_add_51_79_groupi_g41707(csa_tree_add_51_79_groupi_n_4412 ,csa_tree_add_51_79_groupi_n_2669 ,csa_tree_add_51_79_groupi_n_996);
  or csa_tree_add_51_79_groupi_g41708(csa_tree_add_51_79_groupi_n_4411 ,csa_tree_add_51_79_groupi_n_2581 ,csa_tree_add_51_79_groupi_n_430);
  or csa_tree_add_51_79_groupi_g41709(csa_tree_add_51_79_groupi_n_4410 ,csa_tree_add_51_79_groupi_n_2873 ,csa_tree_add_51_79_groupi_n_987);
  or csa_tree_add_51_79_groupi_g41710(csa_tree_add_51_79_groupi_n_4409 ,csa_tree_add_51_79_groupi_n_2668 ,csa_tree_add_51_79_groupi_n_963);
  or csa_tree_add_51_79_groupi_g41711(csa_tree_add_51_79_groupi_n_4408 ,csa_tree_add_51_79_groupi_n_2278 ,csa_tree_add_51_79_groupi_n_349);
  or csa_tree_add_51_79_groupi_g41712(csa_tree_add_51_79_groupi_n_4407 ,csa_tree_add_51_79_groupi_n_2667 ,csa_tree_add_51_79_groupi_n_514);
  or csa_tree_add_51_79_groupi_g41713(csa_tree_add_51_79_groupi_n_4406 ,csa_tree_add_51_79_groupi_n_2171 ,csa_tree_add_51_79_groupi_n_1068);
  or csa_tree_add_51_79_groupi_g41714(csa_tree_add_51_79_groupi_n_4405 ,csa_tree_add_51_79_groupi_n_2292 ,csa_tree_add_51_79_groupi_n_462);
  or csa_tree_add_51_79_groupi_g41715(csa_tree_add_51_79_groupi_n_4404 ,csa_tree_add_51_79_groupi_n_2777 ,csa_tree_add_51_79_groupi_n_438);
  or csa_tree_add_51_79_groupi_g41716(csa_tree_add_51_79_groupi_n_4403 ,csa_tree_add_51_79_groupi_n_2666 ,csa_tree_add_51_79_groupi_n_456);
  or csa_tree_add_51_79_groupi_g41717(csa_tree_add_51_79_groupi_n_4402 ,csa_tree_add_51_79_groupi_n_3275 ,csa_tree_add_51_79_groupi_n_3251);
  nor csa_tree_add_51_79_groupi_g41718(csa_tree_add_51_79_groupi_n_4401 ,csa_tree_add_51_79_groupi_n_3276 ,csa_tree_add_51_79_groupi_n_3252);
  or csa_tree_add_51_79_groupi_g41719(csa_tree_add_51_79_groupi_n_4400 ,csa_tree_add_51_79_groupi_n_2133 ,csa_tree_add_51_79_groupi_n_337);
  or csa_tree_add_51_79_groupi_g41720(csa_tree_add_51_79_groupi_n_4399 ,csa_tree_add_51_79_groupi_n_3288 ,csa_tree_add_51_79_groupi_n_3236);
  or csa_tree_add_51_79_groupi_g41721(csa_tree_add_51_79_groupi_n_4398 ,csa_tree_add_51_79_groupi_n_2186 ,csa_tree_add_51_79_groupi_n_1068);
  or csa_tree_add_51_79_groupi_g41722(csa_tree_add_51_79_groupi_n_4397 ,csa_tree_add_51_79_groupi_n_2318 ,csa_tree_add_51_79_groupi_n_385);
  or csa_tree_add_51_79_groupi_g41723(csa_tree_add_51_79_groupi_n_4396 ,csa_tree_add_51_79_groupi_n_3261 ,csa_tree_add_51_79_groupi_n_3195);
  or csa_tree_add_51_79_groupi_g41724(csa_tree_add_51_79_groupi_n_4395 ,csa_tree_add_51_79_groupi_n_2874 ,csa_tree_add_51_79_groupi_n_500);
  or csa_tree_add_51_79_groupi_g41725(csa_tree_add_51_79_groupi_n_4394 ,csa_tree_add_51_79_groupi_n_2858 ,csa_tree_add_51_79_groupi_n_909);
  nor csa_tree_add_51_79_groupi_g41726(csa_tree_add_51_79_groupi_n_4393 ,csa_tree_add_51_79_groupi_n_3279 ,csa_tree_add_51_79_groupi_n_3778);
  or csa_tree_add_51_79_groupi_g41727(csa_tree_add_51_79_groupi_n_4392 ,csa_tree_add_51_79_groupi_n_2021 ,csa_tree_add_51_79_groupi_n_957);
  or csa_tree_add_51_79_groupi_g41728(csa_tree_add_51_79_groupi_n_4391 ,csa_tree_add_51_79_groupi_n_2238 ,csa_tree_add_51_79_groupi_n_1008);
  or csa_tree_add_51_79_groupi_g41729(csa_tree_add_51_79_groupi_n_4390 ,csa_tree_add_51_79_groupi_n_3257 ,csa_tree_add_51_79_groupi_n_3294);
  or csa_tree_add_51_79_groupi_g41730(csa_tree_add_51_79_groupi_n_4389 ,csa_tree_add_51_79_groupi_n_2197 ,csa_tree_add_51_79_groupi_n_488);
  or csa_tree_add_51_79_groupi_g41731(csa_tree_add_51_79_groupi_n_4388 ,csa_tree_add_51_79_groupi_n_2682 ,csa_tree_add_51_79_groupi_n_930);
  or csa_tree_add_51_79_groupi_g41732(csa_tree_add_51_79_groupi_n_4387 ,csa_tree_add_51_79_groupi_n_2044 ,csa_tree_add_51_79_groupi_n_229);
  or csa_tree_add_51_79_groupi_g41733(csa_tree_add_51_79_groupi_n_4386 ,csa_tree_add_51_79_groupi_n_2230 ,csa_tree_add_51_79_groupi_n_418);
  or csa_tree_add_51_79_groupi_g41734(csa_tree_add_51_79_groupi_n_4385 ,csa_tree_add_51_79_groupi_n_2838 ,csa_tree_add_51_79_groupi_n_981);
  or csa_tree_add_51_79_groupi_g41735(csa_tree_add_51_79_groupi_n_4384 ,csa_tree_add_51_79_groupi_n_2849 ,csa_tree_add_51_79_groupi_n_482);
  or csa_tree_add_51_79_groupi_g41736(csa_tree_add_51_79_groupi_n_4383 ,csa_tree_add_51_79_groupi_n_2635 ,csa_tree_add_51_79_groupi_n_486);
  or csa_tree_add_51_79_groupi_g41737(csa_tree_add_51_79_groupi_n_4382 ,csa_tree_add_51_79_groupi_n_2241 ,csa_tree_add_51_79_groupi_n_897);
  or csa_tree_add_51_79_groupi_g41738(csa_tree_add_51_79_groupi_n_4381 ,csa_tree_add_51_79_groupi_n_2328 ,csa_tree_add_51_79_groupi_n_912);
  or csa_tree_add_51_79_groupi_g41739(csa_tree_add_51_79_groupi_n_4380 ,csa_tree_add_51_79_groupi_n_2309 ,csa_tree_add_51_79_groupi_n_355);
  or csa_tree_add_51_79_groupi_g41740(csa_tree_add_51_79_groupi_n_4379 ,csa_tree_add_51_79_groupi_n_2648 ,csa_tree_add_51_79_groupi_n_277);
  or csa_tree_add_51_79_groupi_g41741(csa_tree_add_51_79_groupi_n_4378 ,csa_tree_add_51_79_groupi_n_2072 ,csa_tree_add_51_79_groupi_n_918);
  or csa_tree_add_51_79_groupi_g41742(csa_tree_add_51_79_groupi_n_4377 ,csa_tree_add_51_79_groupi_n_2646 ,csa_tree_add_51_79_groupi_n_975);
  or csa_tree_add_51_79_groupi_g41743(csa_tree_add_51_79_groupi_n_4376 ,csa_tree_add_51_79_groupi_n_2211 ,csa_tree_add_51_79_groupi_n_1032);
  or csa_tree_add_51_79_groupi_g41744(csa_tree_add_51_79_groupi_n_4375 ,csa_tree_add_51_79_groupi_n_2645 ,csa_tree_add_51_79_groupi_n_1026);
  or csa_tree_add_51_79_groupi_g41745(csa_tree_add_51_79_groupi_n_4374 ,csa_tree_add_51_79_groupi_n_2831 ,csa_tree_add_51_79_groupi_n_492);
  or csa_tree_add_51_79_groupi_g41746(csa_tree_add_51_79_groupi_n_4373 ,csa_tree_add_51_79_groupi_n_2859 ,csa_tree_add_51_79_groupi_n_1029);
  or csa_tree_add_51_79_groupi_g41747(csa_tree_add_51_79_groupi_n_4372 ,csa_tree_add_51_79_groupi_n_2821 ,csa_tree_add_51_79_groupi_n_468);
  or csa_tree_add_51_79_groupi_g41748(csa_tree_add_51_79_groupi_n_4371 ,csa_tree_add_51_79_groupi_n_2659 ,csa_tree_add_51_79_groupi_n_163);
  or csa_tree_add_51_79_groupi_g41749(csa_tree_add_51_79_groupi_n_4370 ,csa_tree_add_51_79_groupi_n_2368 ,csa_tree_add_51_79_groupi_n_948);
  nor csa_tree_add_51_79_groupi_g41750(csa_tree_add_51_79_groupi_n_4369 ,csa_tree_add_51_79_groupi_n_2202 ,csa_tree_add_51_79_groupi_n_1035);
  or csa_tree_add_51_79_groupi_g41751(csa_tree_add_51_79_groupi_n_4368 ,csa_tree_add_51_79_groupi_n_2585 ,csa_tree_add_51_79_groupi_n_520);
  or csa_tree_add_51_79_groupi_g41752(csa_tree_add_51_79_groupi_n_4367 ,csa_tree_add_51_79_groupi_n_3293 ,csa_tree_add_51_79_groupi_n_3209);
  and csa_tree_add_51_79_groupi_g41753(csa_tree_add_51_79_groupi_n_4366 ,csa_tree_add_51_79_groupi_n_3293 ,csa_tree_add_51_79_groupi_n_3209);
  or csa_tree_add_51_79_groupi_g41754(csa_tree_add_51_79_groupi_n_4365 ,csa_tree_add_51_79_groupi_n_3198 ,csa_tree_add_51_79_groupi_n_3201);
  or csa_tree_add_51_79_groupi_g41755(csa_tree_add_51_79_groupi_n_4364 ,csa_tree_add_51_79_groupi_n_1958 ,csa_tree_add_51_79_groupi_n_474);
  or csa_tree_add_51_79_groupi_g41756(csa_tree_add_51_79_groupi_n_4363 ,csa_tree_add_51_79_groupi_n_2712 ,csa_tree_add_51_79_groupi_n_436);
  or csa_tree_add_51_79_groupi_g41757(csa_tree_add_51_79_groupi_n_4362 ,csa_tree_add_51_79_groupi_n_2622 ,csa_tree_add_51_79_groupi_n_476);
  nor csa_tree_add_51_79_groupi_g41758(csa_tree_add_51_79_groupi_n_4361 ,csa_tree_add_51_79_groupi_n_3255 ,csa_tree_add_51_79_groupi_n_3823);
  or csa_tree_add_51_79_groupi_g41759(csa_tree_add_51_79_groupi_n_4360 ,csa_tree_add_51_79_groupi_n_2114 ,csa_tree_add_51_79_groupi_n_1047);
  or csa_tree_add_51_79_groupi_g41760(csa_tree_add_51_79_groupi_n_4359 ,csa_tree_add_51_79_groupi_n_2818 ,csa_tree_add_51_79_groupi_n_518);
  or csa_tree_add_51_79_groupi_g41761(csa_tree_add_51_79_groupi_n_4358 ,csa_tree_add_51_79_groupi_n_3784 ,csa_tree_add_51_79_groupi_n_3826);
  or csa_tree_add_51_79_groupi_g41762(csa_tree_add_51_79_groupi_n_4357 ,csa_tree_add_51_79_groupi_n_2709 ,csa_tree_add_51_79_groupi_n_1062);
  or csa_tree_add_51_79_groupi_g41763(csa_tree_add_51_79_groupi_n_4356 ,csa_tree_add_51_79_groupi_n_2687 ,csa_tree_add_51_79_groupi_n_1056);
  or csa_tree_add_51_79_groupi_g41764(csa_tree_add_51_79_groupi_n_4355 ,csa_tree_add_51_79_groupi_n_2688 ,csa_tree_add_51_79_groupi_n_927);
  or csa_tree_add_51_79_groupi_g41765(csa_tree_add_51_79_groupi_n_4354 ,csa_tree_add_51_79_groupi_n_2639 ,csa_tree_add_51_79_groupi_n_470);
  or csa_tree_add_51_79_groupi_g41766(csa_tree_add_51_79_groupi_n_4353 ,csa_tree_add_51_79_groupi_n_2836 ,csa_tree_add_51_79_groupi_n_458);
  and csa_tree_add_51_79_groupi_g41767(csa_tree_add_51_79_groupi_n_4352 ,csa_tree_add_51_79_groupi_n_3804 ,csa_tree_add_51_79_groupi_n_3210);
  or csa_tree_add_51_79_groupi_g41768(csa_tree_add_51_79_groupi_n_4351 ,csa_tree_add_51_79_groupi_n_2119 ,csa_tree_add_51_79_groupi_n_915);
  or csa_tree_add_51_79_groupi_g41769(csa_tree_add_51_79_groupi_n_4350 ,csa_tree_add_51_79_groupi_n_2811 ,csa_tree_add_51_79_groupi_n_1023);
  or csa_tree_add_51_79_groupi_g41770(csa_tree_add_51_79_groupi_n_4349 ,csa_tree_add_51_79_groupi_n_2199 ,csa_tree_add_51_79_groupi_n_252);
  or csa_tree_add_51_79_groupi_g41771(csa_tree_add_51_79_groupi_n_4348 ,csa_tree_add_51_79_groupi_n_2815 ,csa_tree_add_51_79_groupi_n_954);
  or csa_tree_add_51_79_groupi_g41772(csa_tree_add_51_79_groupi_n_4347 ,csa_tree_add_51_79_groupi_n_2155 ,csa_tree_add_51_79_groupi_n_79);
  or csa_tree_add_51_79_groupi_g41773(csa_tree_add_51_79_groupi_n_4346 ,csa_tree_add_51_79_groupi_n_2213 ,csa_tree_add_51_79_groupi_n_1044);
  or csa_tree_add_51_79_groupi_g41774(csa_tree_add_51_79_groupi_n_4345 ,csa_tree_add_51_79_groupi_n_2577 ,csa_tree_add_51_79_groupi_n_506);
  and csa_tree_add_51_79_groupi_g41775(csa_tree_add_51_79_groupi_n_4344 ,csa_tree_add_51_79_groupi_n_2567 ,csa_tree_add_51_79_groupi_n_3536);
  or csa_tree_add_51_79_groupi_g41776(csa_tree_add_51_79_groupi_n_4343 ,csa_tree_add_51_79_groupi_n_2723 ,csa_tree_add_51_79_groupi_n_951);
  or csa_tree_add_51_79_groupi_g41777(csa_tree_add_51_79_groupi_n_4342 ,csa_tree_add_51_79_groupi_n_2781 ,csa_tree_add_51_79_groupi_n_1065);
  or csa_tree_add_51_79_groupi_g41778(csa_tree_add_51_79_groupi_n_4341 ,csa_tree_add_51_79_groupi_n_2621 ,csa_tree_add_51_79_groupi_n_966);
  or csa_tree_add_51_79_groupi_g41779(csa_tree_add_51_79_groupi_n_4340 ,csa_tree_add_51_79_groupi_n_2153 ,csa_tree_add_51_79_groupi_n_109);
  or csa_tree_add_51_79_groupi_g41780(csa_tree_add_51_79_groupi_n_4339 ,csa_tree_add_51_79_groupi_n_2613 ,csa_tree_add_51_79_groupi_n_199);
  or csa_tree_add_51_79_groupi_g41781(csa_tree_add_51_79_groupi_n_4338 ,csa_tree_add_51_79_groupi_n_2797 ,csa_tree_add_51_79_groupi_n_1017);
  or csa_tree_add_51_79_groupi_g41782(csa_tree_add_51_79_groupi_n_4337 ,csa_tree_add_51_79_groupi_n_2616 ,csa_tree_add_51_79_groupi_n_454);
  or csa_tree_add_51_79_groupi_g41783(csa_tree_add_51_79_groupi_n_4336 ,csa_tree_add_51_79_groupi_n_2865 ,csa_tree_add_51_79_groupi_n_969);
  or csa_tree_add_51_79_groupi_g41784(csa_tree_add_51_79_groupi_n_4335 ,csa_tree_add_51_79_groupi_n_2694 ,csa_tree_add_51_79_groupi_n_241);
  or csa_tree_add_51_79_groupi_g41785(csa_tree_add_51_79_groupi_n_4334 ,csa_tree_add_51_79_groupi_n_2692 ,csa_tree_add_51_79_groupi_n_151);
  or csa_tree_add_51_79_groupi_g41786(csa_tree_add_51_79_groupi_n_4333 ,csa_tree_add_51_79_groupi_n_2608 ,csa_tree_add_51_79_groupi_n_903);
  or csa_tree_add_51_79_groupi_g41787(csa_tree_add_51_79_groupi_n_4332 ,csa_tree_add_51_79_groupi_n_2636 ,csa_tree_add_51_79_groupi_n_924);
  or csa_tree_add_51_79_groupi_g41788(csa_tree_add_51_79_groupi_n_4331 ,csa_tree_add_51_79_groupi_n_2200 ,csa_tree_add_51_79_groupi_n_79);
  or csa_tree_add_51_79_groupi_g41789(csa_tree_add_51_79_groupi_n_4330 ,csa_tree_add_51_79_groupi_n_2884 ,csa_tree_add_51_79_groupi_n_452);
  or csa_tree_add_51_79_groupi_g41790(csa_tree_add_51_79_groupi_n_4329 ,csa_tree_add_51_79_groupi_n_2595 ,csa_tree_add_51_79_groupi_n_55);
  or csa_tree_add_51_79_groupi_g41791(csa_tree_add_51_79_groupi_n_4328 ,csa_tree_add_51_79_groupi_n_2205 ,csa_tree_add_51_79_groupi_n_939);
  or csa_tree_add_51_79_groupi_g41792(csa_tree_add_51_79_groupi_n_4327 ,csa_tree_add_51_79_groupi_n_2025 ,csa_tree_add_51_79_groupi_n_894);
  or csa_tree_add_51_79_groupi_g41793(csa_tree_add_51_79_groupi_n_4326 ,csa_tree_add_51_79_groupi_n_2603 ,csa_tree_add_51_79_groupi_n_900);
  or csa_tree_add_51_79_groupi_g41794(csa_tree_add_51_79_groupi_n_4325 ,csa_tree_add_51_79_groupi_n_2356 ,csa_tree_add_51_79_groupi_n_1020);
  or csa_tree_add_51_79_groupi_g41795(csa_tree_add_51_79_groupi_n_4324 ,csa_tree_add_51_79_groupi_n_2760 ,csa_tree_add_51_79_groupi_n_1065);
  or csa_tree_add_51_79_groupi_g41796(csa_tree_add_51_79_groupi_n_4323 ,csa_tree_add_51_79_groupi_n_1813 ,csa_tree_add_51_79_groupi_n_990);
  or csa_tree_add_51_79_groupi_g41797(csa_tree_add_51_79_groupi_n_4322 ,csa_tree_add_51_79_groupi_n_2178 ,csa_tree_add_51_79_groupi_n_247);
  or csa_tree_add_51_79_groupi_g41798(csa_tree_add_51_79_groupi_n_4321 ,csa_tree_add_51_79_groupi_n_2087 ,csa_tree_add_51_79_groupi_n_480);
  or csa_tree_add_51_79_groupi_g41799(csa_tree_add_51_79_groupi_n_4320 ,csa_tree_add_51_79_groupi_n_3265 ,csa_tree_add_51_79_groupi_n_3287);
  and csa_tree_add_51_79_groupi_g41800(csa_tree_add_51_79_groupi_n_4319 ,csa_tree_add_51_79_groupi_n_3265 ,csa_tree_add_51_79_groupi_n_3287);
  or csa_tree_add_51_79_groupi_g41801(csa_tree_add_51_79_groupi_n_4318 ,csa_tree_add_51_79_groupi_n_2109 ,csa_tree_add_51_79_groupi_n_960);
  and csa_tree_add_51_79_groupi_g41802(csa_tree_add_51_79_groupi_n_4317 ,csa_tree_add_51_79_groupi_n_3208 ,csa_tree_add_51_79_groupi_n_3200);
  or csa_tree_add_51_79_groupi_g41803(csa_tree_add_51_79_groupi_n_4316 ,csa_tree_add_51_79_groupi_n_3754 ,csa_tree_add_51_79_groupi_n_3248);
  or csa_tree_add_51_79_groupi_g41804(csa_tree_add_51_79_groupi_n_4315 ,csa_tree_add_51_79_groupi_n_2775 ,csa_tree_add_51_79_groupi_n_1002);
  or csa_tree_add_51_79_groupi_g41805(csa_tree_add_51_79_groupi_n_4314 ,csa_tree_add_51_79_groupi_n_2620 ,csa_tree_add_51_79_groupi_n_85);
  or csa_tree_add_51_79_groupi_g41806(csa_tree_add_51_79_groupi_n_4313 ,csa_tree_add_51_79_groupi_n_2826 ,csa_tree_add_51_79_groupi_n_984);
  or csa_tree_add_51_79_groupi_g41807(csa_tree_add_51_79_groupi_n_4312 ,csa_tree_add_51_79_groupi_n_2588 ,csa_tree_add_51_79_groupi_n_906);
  or csa_tree_add_51_79_groupi_g41808(csa_tree_add_51_79_groupi_n_4311 ,csa_tree_add_51_79_groupi_n_2223 ,csa_tree_add_51_79_groupi_n_1047);
  or csa_tree_add_51_79_groupi_g41809(csa_tree_add_51_79_groupi_n_4310 ,csa_tree_add_51_79_groupi_n_1940 ,csa_tree_add_51_79_groupi_n_67);
  or csa_tree_add_51_79_groupi_g41810(csa_tree_add_51_79_groupi_n_4309 ,csa_tree_add_51_79_groupi_n_2032 ,csa_tree_add_51_79_groupi_n_999);
  or csa_tree_add_51_79_groupi_g41811(csa_tree_add_51_79_groupi_n_4308 ,csa_tree_add_51_79_groupi_n_2340 ,csa_tree_add_51_79_groupi_n_987);
  or csa_tree_add_51_79_groupi_g41812(csa_tree_add_51_79_groupi_n_4307 ,csa_tree_add_51_79_groupi_n_2198 ,csa_tree_add_51_79_groupi_n_978);
  or csa_tree_add_51_79_groupi_g41813(csa_tree_add_51_79_groupi_n_4306 ,csa_tree_add_51_79_groupi_n_2728 ,csa_tree_add_51_79_groupi_n_912);
  or csa_tree_add_51_79_groupi_g41814(csa_tree_add_51_79_groupi_n_4713 ,csa_tree_add_51_79_groupi_n_3776 ,csa_tree_add_51_79_groupi_n_3744);
  and csa_tree_add_51_79_groupi_g41815(csa_tree_add_51_79_groupi_n_4712 ,csa_tree_add_51_79_groupi_n_3250 ,csa_tree_add_51_79_groupi_n_3786);
  or csa_tree_add_51_79_groupi_g41816(csa_tree_add_51_79_groupi_n_4711 ,csa_tree_add_51_79_groupi_n_3273 ,csa_tree_add_51_79_groupi_n_3736);
  not csa_tree_add_51_79_groupi_g41829(csa_tree_add_51_79_groupi_n_4282 ,csa_tree_add_51_79_groupi_n_4283);
  not csa_tree_add_51_79_groupi_g41830(csa_tree_add_51_79_groupi_n_4281 ,csa_tree_add_51_79_groupi_n_4280);
  not csa_tree_add_51_79_groupi_g41831(csa_tree_add_51_79_groupi_n_4278 ,csa_tree_add_51_79_groupi_n_4279);
  not csa_tree_add_51_79_groupi_g41832(csa_tree_add_51_79_groupi_n_4277 ,csa_tree_add_51_79_groupi_n_4276);
  not csa_tree_add_51_79_groupi_g41833(csa_tree_add_51_79_groupi_n_4274 ,csa_tree_add_51_79_groupi_n_4275);
  not csa_tree_add_51_79_groupi_g41834(csa_tree_add_51_79_groupi_n_4272 ,csa_tree_add_51_79_groupi_n_4273);
  not csa_tree_add_51_79_groupi_g41835(csa_tree_add_51_79_groupi_n_4270 ,csa_tree_add_51_79_groupi_n_4271);
  not csa_tree_add_51_79_groupi_g41836(csa_tree_add_51_79_groupi_n_4269 ,csa_tree_add_51_79_groupi_n_4268);
  not csa_tree_add_51_79_groupi_g41837(csa_tree_add_51_79_groupi_n_4266 ,csa_tree_add_51_79_groupi_n_4265);
  not csa_tree_add_51_79_groupi_g41838(csa_tree_add_51_79_groupi_n_4263 ,csa_tree_add_51_79_groupi_n_4264);
  not csa_tree_add_51_79_groupi_g41839(csa_tree_add_51_79_groupi_n_4261 ,csa_tree_add_51_79_groupi_n_4262);
  not csa_tree_add_51_79_groupi_g41840(csa_tree_add_51_79_groupi_n_4259 ,csa_tree_add_51_79_groupi_n_4258);
  not csa_tree_add_51_79_groupi_g41841(csa_tree_add_51_79_groupi_n_4256 ,csa_tree_add_51_79_groupi_n_4257);
  not csa_tree_add_51_79_groupi_g41842(csa_tree_add_51_79_groupi_n_4255 ,csa_tree_add_51_79_groupi_n_4254);
  not csa_tree_add_51_79_groupi_g41843(csa_tree_add_51_79_groupi_n_4252 ,csa_tree_add_51_79_groupi_n_4253);
  not csa_tree_add_51_79_groupi_g41844(csa_tree_add_51_79_groupi_n_4251 ,csa_tree_add_51_79_groupi_n_4250);
  not csa_tree_add_51_79_groupi_g41845(csa_tree_add_51_79_groupi_n_4248 ,csa_tree_add_51_79_groupi_n_4249);
  not csa_tree_add_51_79_groupi_g41846(csa_tree_add_51_79_groupi_n_4247 ,csa_tree_add_51_79_groupi_n_4246);
  not csa_tree_add_51_79_groupi_g41847(csa_tree_add_51_79_groupi_n_4245 ,csa_tree_add_51_79_groupi_n_4244);
  not csa_tree_add_51_79_groupi_g41848(csa_tree_add_51_79_groupi_n_4242 ,csa_tree_add_51_79_groupi_n_4241);
  not csa_tree_add_51_79_groupi_g41849(csa_tree_add_51_79_groupi_n_4239 ,csa_tree_add_51_79_groupi_n_4240);
  not csa_tree_add_51_79_groupi_g41850(csa_tree_add_51_79_groupi_n_4238 ,csa_tree_add_51_79_groupi_n_4237);
  not csa_tree_add_51_79_groupi_g41851(csa_tree_add_51_79_groupi_n_4232 ,csa_tree_add_51_79_groupi_n_4233);
  not csa_tree_add_51_79_groupi_g41852(csa_tree_add_51_79_groupi_n_4228 ,csa_tree_add_51_79_groupi_n_4227);
  or csa_tree_add_51_79_groupi_g41853(csa_tree_add_51_79_groupi_n_4224 ,csa_tree_add_51_79_groupi_n_2855 ,csa_tree_add_51_79_groupi_n_49);
  or csa_tree_add_51_79_groupi_g41854(csa_tree_add_51_79_groupi_n_4223 ,csa_tree_add_51_79_groupi_n_2416 ,csa_tree_add_51_79_groupi_n_127);
  or csa_tree_add_51_79_groupi_g41855(csa_tree_add_51_79_groupi_n_4222 ,csa_tree_add_51_79_groupi_n_2045 ,csa_tree_add_51_79_groupi_n_921);
  or csa_tree_add_51_79_groupi_g41856(csa_tree_add_51_79_groupi_n_4221 ,csa_tree_add_51_79_groupi_n_2366 ,csa_tree_add_51_79_groupi_n_1014);
  or csa_tree_add_51_79_groupi_g41857(csa_tree_add_51_79_groupi_n_4220 ,csa_tree_add_51_79_groupi_n_2327 ,csa_tree_add_51_79_groupi_n_343);
  or csa_tree_add_51_79_groupi_g41858(csa_tree_add_51_79_groupi_n_4219 ,csa_tree_add_51_79_groupi_n_2136 ,csa_tree_add_51_79_groupi_n_133);
  or csa_tree_add_51_79_groupi_g41859(csa_tree_add_51_79_groupi_n_4218 ,csa_tree_add_51_79_groupi_n_2793 ,csa_tree_add_51_79_groupi_n_163);
  or csa_tree_add_51_79_groupi_g41860(csa_tree_add_51_79_groupi_n_4217 ,csa_tree_add_51_79_groupi_n_2825 ,csa_tree_add_51_79_groupi_n_265);
  or csa_tree_add_51_79_groupi_g41861(csa_tree_add_51_79_groupi_n_4216 ,csa_tree_add_51_79_groupi_n_2042 ,csa_tree_add_51_79_groupi_n_223);
  or csa_tree_add_51_79_groupi_g41862(csa_tree_add_51_79_groupi_n_4215 ,csa_tree_add_51_79_groupi_n_2737 ,csa_tree_add_51_79_groupi_n_217);
  or csa_tree_add_51_79_groupi_g41863(csa_tree_add_51_79_groupi_n_4214 ,csa_tree_add_51_79_groupi_n_2756 ,csa_tree_add_51_79_groupi_n_1050);
  or csa_tree_add_51_79_groupi_g41864(csa_tree_add_51_79_groupi_n_4213 ,csa_tree_add_51_79_groupi_n_2151 ,csa_tree_add_51_79_groupi_n_367);
  or csa_tree_add_51_79_groupi_g41865(csa_tree_add_51_79_groupi_n_4212 ,csa_tree_add_51_79_groupi_n_2583 ,csa_tree_add_51_79_groupi_n_448);
  or csa_tree_add_51_79_groupi_g41866(csa_tree_add_51_79_groupi_n_4211 ,csa_tree_add_51_79_groupi_n_2115 ,csa_tree_add_51_79_groupi_n_145);
  or csa_tree_add_51_79_groupi_g41867(csa_tree_add_51_79_groupi_n_4210 ,csa_tree_add_51_79_groupi_n_2090 ,csa_tree_add_51_79_groupi_n_103);
  or csa_tree_add_51_79_groupi_g41868(csa_tree_add_51_79_groupi_n_4209 ,csa_tree_add_51_79_groupi_n_2291 ,csa_tree_add_51_79_groupi_n_211);
  or csa_tree_add_51_79_groupi_g41869(csa_tree_add_51_79_groupi_n_4208 ,csa_tree_add_51_79_groupi_n_2619 ,csa_tree_add_51_79_groupi_n_933);
  or csa_tree_add_51_79_groupi_g41870(csa_tree_add_51_79_groupi_n_4207 ,csa_tree_add_51_79_groupi_n_2068 ,csa_tree_add_51_79_groupi_n_993);
  or csa_tree_add_51_79_groupi_g41871(csa_tree_add_51_79_groupi_n_4206 ,csa_tree_add_51_79_groupi_n_2016 ,csa_tree_add_51_79_groupi_n_942);
  or csa_tree_add_51_79_groupi_g41872(csa_tree_add_51_79_groupi_n_4205 ,csa_tree_add_51_79_groupi_n_2572 ,csa_tree_add_51_79_groupi_n_133);
  or csa_tree_add_51_79_groupi_g41873(csa_tree_add_51_79_groupi_n_4204 ,csa_tree_add_51_79_groupi_n_2018 ,csa_tree_add_51_79_groupi_n_504);
  or csa_tree_add_51_79_groupi_g41874(csa_tree_add_51_79_groupi_n_4203 ,csa_tree_add_51_79_groupi_n_1800 ,csa_tree_add_51_79_groupi_n_169);
  or csa_tree_add_51_79_groupi_g41875(csa_tree_add_51_79_groupi_n_4202 ,csa_tree_add_51_79_groupi_n_2299 ,csa_tree_add_51_79_groupi_n_61);
  or csa_tree_add_51_79_groupi_g41876(csa_tree_add_51_79_groupi_n_4201 ,csa_tree_add_51_79_groupi_n_2226 ,csa_tree_add_51_79_groupi_n_1062);
  or csa_tree_add_51_79_groupi_g41877(csa_tree_add_51_79_groupi_n_4200 ,csa_tree_add_51_79_groupi_n_2203 ,csa_tree_add_51_79_groupi_n_45);
  or csa_tree_add_51_79_groupi_g41878(csa_tree_add_51_79_groupi_n_4199 ,csa_tree_add_51_79_groupi_n_2841 ,csa_tree_add_51_79_groupi_n_502);
  or csa_tree_add_51_79_groupi_g41879(csa_tree_add_51_79_groupi_n_4198 ,csa_tree_add_51_79_groupi_n_2810 ,csa_tree_add_51_79_groupi_n_355);
  or csa_tree_add_51_79_groupi_g41880(csa_tree_add_51_79_groupi_n_4197 ,csa_tree_add_51_79_groupi_n_2785 ,csa_tree_add_51_79_groupi_n_918);
  or csa_tree_add_51_79_groupi_g41881(csa_tree_add_51_79_groupi_n_4196 ,csa_tree_add_51_79_groupi_n_2584 ,csa_tree_add_51_79_groupi_n_307);
  or csa_tree_add_51_79_groupi_g41882(csa_tree_add_51_79_groupi_n_4195 ,csa_tree_add_51_79_groupi_n_2606 ,csa_tree_add_51_79_groupi_n_121);
  or csa_tree_add_51_79_groupi_g41883(csa_tree_add_51_79_groupi_n_4194 ,csa_tree_add_51_79_groupi_n_3199 ,csa_tree_add_51_79_groupi_n_3298);
  or csa_tree_add_51_79_groupi_g41884(csa_tree_add_51_79_groupi_n_4193 ,csa_tree_add_51_79_groupi_n_2157 ,csa_tree_add_51_79_groupi_n_444);
  or csa_tree_add_51_79_groupi_g41885(csa_tree_add_51_79_groupi_n_4192 ,csa_tree_add_51_79_groupi_n_3230 ,csa_tree_add_51_79_groupi_n_3270);
  and csa_tree_add_51_79_groupi_g41886(csa_tree_add_51_79_groupi_n_4191 ,csa_tree_add_51_79_groupi_n_3230 ,csa_tree_add_51_79_groupi_n_3270);
  or csa_tree_add_51_79_groupi_g41887(csa_tree_add_51_79_groupi_n_4190 ,csa_tree_add_51_79_groupi_n_2695 ,csa_tree_add_51_79_groupi_n_271);
  or csa_tree_add_51_79_groupi_g41888(csa_tree_add_51_79_groupi_n_4189 ,csa_tree_add_51_79_groupi_n_2653 ,csa_tree_add_51_79_groupi_n_936);
  or csa_tree_add_51_79_groupi_g41889(csa_tree_add_51_79_groupi_n_4188 ,csa_tree_add_51_79_groupi_n_2218 ,csa_tree_add_51_79_groupi_n_1068);
  or csa_tree_add_51_79_groupi_g41890(csa_tree_add_51_79_groupi_n_4187 ,csa_tree_add_51_79_groupi_n_2027 ,csa_tree_add_51_79_groupi_n_510);
  or csa_tree_add_51_79_groupi_g41891(csa_tree_add_51_79_groupi_n_4186 ,csa_tree_add_51_79_groupi_n_3737 ,csa_tree_add_51_79_groupi_n_3243);
  or csa_tree_add_51_79_groupi_g41892(csa_tree_add_51_79_groupi_n_4185 ,csa_tree_add_51_79_groupi_n_2283 ,csa_tree_add_51_79_groupi_n_283);
  or csa_tree_add_51_79_groupi_g41893(csa_tree_add_51_79_groupi_n_4184 ,csa_tree_add_51_79_groupi_n_2615 ,csa_tree_add_51_79_groupi_n_906);
  or csa_tree_add_51_79_groupi_g41894(csa_tree_add_51_79_groupi_n_4183 ,csa_tree_add_51_79_groupi_n_2123 ,csa_tree_add_51_79_groupi_n_440);
  or csa_tree_add_51_79_groupi_g41895(csa_tree_add_51_79_groupi_n_4182 ,csa_tree_add_51_79_groupi_n_2311 ,csa_tree_add_51_79_groupi_n_1020);
  or csa_tree_add_51_79_groupi_g41896(csa_tree_add_51_79_groupi_n_4181 ,csa_tree_add_51_79_groupi_n_2869 ,csa_tree_add_51_79_groupi_n_187);
  or csa_tree_add_51_79_groupi_g41897(csa_tree_add_51_79_groupi_n_4180 ,csa_tree_add_51_79_groupi_n_2183 ,csa_tree_add_51_79_groupi_n_1005);
  or csa_tree_add_51_79_groupi_g41898(csa_tree_add_51_79_groupi_n_4179 ,csa_tree_add_51_79_groupi_n_2034 ,csa_tree_add_51_79_groupi_n_211);
  or csa_tree_add_51_79_groupi_g41899(csa_tree_add_51_79_groupi_n_4178 ,csa_tree_add_51_79_groupi_n_2721 ,csa_tree_add_51_79_groupi_n_61);
  or csa_tree_add_51_79_groupi_g41900(csa_tree_add_51_79_groupi_n_4177 ,csa_tree_add_51_79_groupi_n_2089 ,csa_tree_add_51_79_groupi_n_951);
  or csa_tree_add_51_79_groupi_g41901(csa_tree_add_51_79_groupi_n_4176 ,csa_tree_add_51_79_groupi_n_2587 ,csa_tree_add_51_79_groupi_n_1029);
  or csa_tree_add_51_79_groupi_g41902(csa_tree_add_51_79_groupi_n_4175 ,csa_tree_add_51_79_groupi_n_2780 ,csa_tree_add_51_79_groupi_n_240);
  or csa_tree_add_51_79_groupi_g41903(csa_tree_add_51_79_groupi_n_4174 ,csa_tree_add_51_79_groupi_n_2091 ,csa_tree_add_51_79_groupi_n_121);
  or csa_tree_add_51_79_groupi_g41904(csa_tree_add_51_79_groupi_n_4173 ,csa_tree_add_51_79_groupi_n_2661 ,csa_tree_add_51_79_groupi_n_891);
  and csa_tree_add_51_79_groupi_g41905(csa_tree_add_51_79_groupi_n_4172 ,csa_tree_add_51_79_groupi_n_3207 ,csa_tree_add_51_79_groupi_n_3224);
  or csa_tree_add_51_79_groupi_g41906(csa_tree_add_51_79_groupi_n_4171 ,csa_tree_add_51_79_groupi_n_2195 ,csa_tree_add_51_79_groupi_n_91);
  or csa_tree_add_51_79_groupi_g41907(csa_tree_add_51_79_groupi_n_4170 ,csa_tree_add_51_79_groupi_n_2866 ,csa_tree_add_51_79_groupi_n_307);
  or csa_tree_add_51_79_groupi_g41908(csa_tree_add_51_79_groupi_n_4169 ,csa_tree_add_51_79_groupi_n_2579 ,csa_tree_add_51_79_groupi_n_228);
  or csa_tree_add_51_79_groupi_g41909(csa_tree_add_51_79_groupi_n_4168 ,csa_tree_add_51_79_groupi_n_2727 ,csa_tree_add_51_79_groupi_n_379);
  or csa_tree_add_51_79_groupi_g41910(csa_tree_add_51_79_groupi_n_4167 ,csa_tree_add_51_79_groupi_n_2852 ,csa_tree_add_51_79_groupi_n_373);
  or csa_tree_add_51_79_groupi_g41911(csa_tree_add_51_79_groupi_n_4166 ,csa_tree_add_51_79_groupi_n_2059 ,csa_tree_add_51_79_groupi_n_289);
  or csa_tree_add_51_79_groupi_g41912(csa_tree_add_51_79_groupi_n_4165 ,csa_tree_add_51_79_groupi_n_2663 ,csa_tree_add_51_79_groupi_n_397);
  or csa_tree_add_51_79_groupi_g41913(csa_tree_add_51_79_groupi_n_4164 ,csa_tree_add_51_79_groupi_n_2273 ,csa_tree_add_51_79_groupi_n_1053);
  or csa_tree_add_51_79_groupi_g41914(csa_tree_add_51_79_groupi_n_4163 ,csa_tree_add_51_79_groupi_n_2248 ,csa_tree_add_51_79_groupi_n_295);
  or csa_tree_add_51_79_groupi_g41915(csa_tree_add_51_79_groupi_n_4162 ,csa_tree_add_51_79_groupi_n_2689 ,csa_tree_add_51_79_groupi_n_325);
  or csa_tree_add_51_79_groupi_g41916(csa_tree_add_51_79_groupi_n_4161 ,csa_tree_add_51_79_groupi_n_2598 ,csa_tree_add_51_79_groupi_n_957);
  or csa_tree_add_51_79_groupi_g41917(csa_tree_add_51_79_groupi_n_4160 ,csa_tree_add_51_79_groupi_n_2681 ,csa_tree_add_51_79_groupi_n_993);
  or csa_tree_add_51_79_groupi_g41918(csa_tree_add_51_79_groupi_n_4159 ,csa_tree_add_51_79_groupi_n_2638 ,csa_tree_add_51_79_groupi_n_348);
  or csa_tree_add_51_79_groupi_g41919(csa_tree_add_51_79_groupi_n_4158 ,csa_tree_add_51_79_groupi_n_2125 ,csa_tree_add_51_79_groupi_n_1011);
  or csa_tree_add_51_79_groupi_g41920(csa_tree_add_51_79_groupi_n_4157 ,csa_tree_add_51_79_groupi_n_2827 ,csa_tree_add_51_79_groupi_n_1038);
  or csa_tree_add_51_79_groupi_g41921(csa_tree_add_51_79_groupi_n_4156 ,csa_tree_add_51_79_groupi_n_2624 ,csa_tree_add_51_79_groupi_n_1017);
  or csa_tree_add_51_79_groupi_g41922(csa_tree_add_51_79_groupi_n_4155 ,csa_tree_add_51_79_groupi_n_2745 ,csa_tree_add_51_79_groupi_n_271);
  or csa_tree_add_51_79_groupi_g41923(csa_tree_add_51_79_groupi_n_4154 ,csa_tree_add_51_79_groupi_n_2644 ,csa_tree_add_51_79_groupi_n_379);
  or csa_tree_add_51_79_groupi_g41924(csa_tree_add_51_79_groupi_n_4153 ,csa_tree_add_51_79_groupi_n_2187 ,csa_tree_add_51_79_groupi_n_412);
  or csa_tree_add_51_79_groupi_g41925(csa_tree_add_51_79_groupi_n_4152 ,csa_tree_add_51_79_groupi_n_2088 ,csa_tree_add_51_79_groupi_n_1065);
  and csa_tree_add_51_79_groupi_g41926(csa_tree_add_51_79_groupi_n_4151 ,csa_tree_add_51_79_groupi_n_3206 ,csa_tree_add_51_79_groupi_n_3194);
  or csa_tree_add_51_79_groupi_g41927(csa_tree_add_51_79_groupi_n_4150 ,csa_tree_add_51_79_groupi_n_2730 ,csa_tree_add_51_79_groupi_n_181);
  or csa_tree_add_51_79_groupi_g41928(csa_tree_add_51_79_groupi_n_4149 ,csa_tree_add_51_79_groupi_n_2049 ,csa_tree_add_51_79_groupi_n_397);
  or csa_tree_add_51_79_groupi_g41929(csa_tree_add_51_79_groupi_n_4148 ,csa_tree_add_51_79_groupi_n_2170 ,csa_tree_add_51_79_groupi_n_283);
  or csa_tree_add_51_79_groupi_g41930(csa_tree_add_51_79_groupi_n_4147 ,csa_tree_add_51_79_groupi_n_2355 ,csa_tree_add_51_79_groupi_n_1026);
  or csa_tree_add_51_79_groupi_g41931(csa_tree_add_51_79_groupi_n_4146 ,csa_tree_add_51_79_groupi_n_2110 ,csa_tree_add_51_79_groupi_n_909);
  or csa_tree_add_51_79_groupi_g41932(csa_tree_add_51_79_groupi_n_4145 ,csa_tree_add_51_79_groupi_n_2324 ,csa_tree_add_51_79_groupi_n_103);
  or csa_tree_add_51_79_groupi_g41933(csa_tree_add_51_79_groupi_n_4144 ,csa_tree_add_51_79_groupi_n_1794 ,csa_tree_add_51_79_groupi_n_85);
  or csa_tree_add_51_79_groupi_g41934(csa_tree_add_51_79_groupi_n_4143 ,csa_tree_add_51_79_groupi_n_1893 ,csa_tree_add_51_79_groupi_n_385);
  or csa_tree_add_51_79_groupi_g41935(csa_tree_add_51_79_groupi_n_4142 ,csa_tree_add_51_79_groupi_n_2050 ,csa_tree_add_51_79_groupi_n_139);
  or csa_tree_add_51_79_groupi_g41936(csa_tree_add_51_79_groupi_n_4141 ,csa_tree_add_51_79_groupi_n_1956 ,csa_tree_add_51_79_groupi_n_205);
  or csa_tree_add_51_79_groupi_g41937(csa_tree_add_51_79_groupi_n_4140 ,csa_tree_add_51_79_groupi_n_2270 ,csa_tree_add_51_79_groupi_n_1059);
  or csa_tree_add_51_79_groupi_g41938(csa_tree_add_51_79_groupi_n_4139 ,csa_tree_add_51_79_groupi_n_2671 ,csa_tree_add_51_79_groupi_n_313);
  or csa_tree_add_51_79_groupi_g41939(csa_tree_add_51_79_groupi_n_4138 ,csa_tree_add_51_79_groupi_n_1881 ,csa_tree_add_51_79_groupi_n_199);
  or csa_tree_add_51_79_groupi_g41940(csa_tree_add_51_79_groupi_n_4137 ,csa_tree_add_51_79_groupi_n_2053 ,csa_tree_add_51_79_groupi_n_894);
  or csa_tree_add_51_79_groupi_g41941(csa_tree_add_51_79_groupi_n_4136 ,csa_tree_add_51_79_groupi_n_3262 ,csa_tree_add_51_79_groupi_n_3203);
  or csa_tree_add_51_79_groupi_g41942(csa_tree_add_51_79_groupi_n_4135 ,csa_tree_add_51_79_groupi_n_2074 ,csa_tree_add_51_79_groupi_n_1050);
  or csa_tree_add_51_79_groupi_g41943(csa_tree_add_51_79_groupi_n_4134 ,csa_tree_add_51_79_groupi_n_2614 ,csa_tree_add_51_79_groupi_n_361);
  or csa_tree_add_51_79_groupi_g41944(csa_tree_add_51_79_groupi_n_4133 ,csa_tree_add_51_79_groupi_n_2599 ,csa_tree_add_51_79_groupi_n_319);
  or csa_tree_add_51_79_groupi_g41945(csa_tree_add_51_79_groupi_n_4132 ,csa_tree_add_51_79_groupi_n_2308 ,csa_tree_add_51_79_groupi_n_945);
  or csa_tree_add_51_79_groupi_g41946(csa_tree_add_51_79_groupi_n_4131 ,csa_tree_add_51_79_groupi_n_3254 ,csa_tree_add_51_79_groupi_n_3822);
  or csa_tree_add_51_79_groupi_g41947(csa_tree_add_51_79_groupi_n_4130 ,csa_tree_add_51_79_groupi_n_1965 ,csa_tree_add_51_79_groupi_n_175);
  or csa_tree_add_51_79_groupi_g41948(csa_tree_add_51_79_groupi_n_4129 ,csa_tree_add_51_79_groupi_n_2835 ,csa_tree_add_51_79_groupi_n_187);
  or csa_tree_add_51_79_groupi_g41949(csa_tree_add_51_79_groupi_n_4128 ,csa_tree_add_51_79_groupi_n_2210 ,csa_tree_add_51_79_groupi_n_337);
  or csa_tree_add_51_79_groupi_g41950(csa_tree_add_51_79_groupi_n_4127 ,csa_tree_add_51_79_groupi_n_2686 ,csa_tree_add_51_79_groupi_n_289);
  or csa_tree_add_51_79_groupi_g41951(csa_tree_add_51_79_groupi_n_4126 ,csa_tree_add_51_79_groupi_n_2656 ,csa_tree_add_51_79_groupi_n_373);
  or csa_tree_add_51_79_groupi_g41952(csa_tree_add_51_79_groupi_n_4125 ,csa_tree_add_51_79_groupi_n_2319 ,csa_tree_add_51_79_groupi_n_319);
  or csa_tree_add_51_79_groupi_g41953(csa_tree_add_51_79_groupi_n_4124 ,csa_tree_add_51_79_groupi_n_2696 ,csa_tree_add_51_79_groupi_n_313);
  or csa_tree_add_51_79_groupi_g41954(csa_tree_add_51_79_groupi_n_4123 ,csa_tree_add_51_79_groupi_n_2594 ,csa_tree_add_51_79_groupi_n_915);
  or csa_tree_add_51_79_groupi_g41955(csa_tree_add_51_79_groupi_n_4122 ,csa_tree_add_51_79_groupi_n_2776 ,csa_tree_add_51_79_groupi_n_361);
  or csa_tree_add_51_79_groupi_g41956(csa_tree_add_51_79_groupi_n_4121 ,csa_tree_add_51_79_groupi_n_1896 ,csa_tree_add_51_79_groupi_n_984);
  or csa_tree_add_51_79_groupi_g41957(csa_tree_add_51_79_groupi_n_4120 ,csa_tree_add_51_79_groupi_n_2189 ,csa_tree_add_51_79_groupi_n_73);
  or csa_tree_add_51_79_groupi_g41958(csa_tree_add_51_79_groupi_n_4119 ,csa_tree_add_51_79_groupi_n_2596 ,csa_tree_add_51_79_groupi_n_169);
  or csa_tree_add_51_79_groupi_g41959(csa_tree_add_51_79_groupi_n_4118 ,csa_tree_add_51_79_groupi_n_1876 ,csa_tree_add_51_79_groupi_n_301);
  or csa_tree_add_51_79_groupi_g41960(csa_tree_add_51_79_groupi_n_4117 ,csa_tree_add_51_79_groupi_n_3208 ,csa_tree_add_51_79_groupi_n_3200);
  or csa_tree_add_51_79_groupi_g41961(csa_tree_add_51_79_groupi_n_4116 ,csa_tree_add_51_79_groupi_n_2017 ,csa_tree_add_51_79_groupi_n_193);
  or csa_tree_add_51_79_groupi_g41962(csa_tree_add_51_79_groupi_n_4115 ,csa_tree_add_51_79_groupi_n_2799 ,csa_tree_add_51_79_groupi_n_942);
  or csa_tree_add_51_79_groupi_g41963(csa_tree_add_51_79_groupi_n_4114 ,csa_tree_add_51_79_groupi_n_2067 ,csa_tree_add_51_79_groupi_n_127);
  or csa_tree_add_51_79_groupi_g41964(csa_tree_add_51_79_groupi_n_4113 ,csa_tree_add_51_79_groupi_n_2224 ,csa_tree_add_51_79_groupi_n_1035);
  or csa_tree_add_51_79_groupi_g41965(csa_tree_add_51_79_groupi_n_4112 ,csa_tree_add_51_79_groupi_n_2152 ,csa_tree_add_51_79_groupi_n_109);
  or csa_tree_add_51_79_groupi_g41966(csa_tree_add_51_79_groupi_n_4111 ,csa_tree_add_51_79_groupi_n_2677 ,csa_tree_add_51_79_groupi_n_331);
  or csa_tree_add_51_79_groupi_g41967(csa_tree_add_51_79_groupi_n_4110 ,csa_tree_add_51_79_groupi_n_2798 ,csa_tree_add_51_79_groupi_n_139);
  or csa_tree_add_51_79_groupi_g41968(csa_tree_add_51_79_groupi_n_4109 ,csa_tree_add_51_79_groupi_n_2763 ,csa_tree_add_51_79_groupi_n_175);
  or csa_tree_add_51_79_groupi_g41969(csa_tree_add_51_79_groupi_n_4108 ,csa_tree_add_51_79_groupi_n_2037 ,csa_tree_add_51_79_groupi_n_331);
  or csa_tree_add_51_79_groupi_g41970(csa_tree_add_51_79_groupi_n_4107 ,csa_tree_add_51_79_groupi_n_2065 ,csa_tree_add_51_79_groupi_n_145);
  or csa_tree_add_51_79_groupi_g41971(csa_tree_add_51_79_groupi_n_4106 ,csa_tree_add_51_79_groupi_n_2219 ,csa_tree_add_51_79_groupi_n_295);
  or csa_tree_add_51_79_groupi_g41972(csa_tree_add_51_79_groupi_n_4105 ,csa_tree_add_51_79_groupi_n_2300 ,csa_tree_add_51_79_groupi_n_936);
  or csa_tree_add_51_79_groupi_g41973(csa_tree_add_51_79_groupi_n_4104 ,csa_tree_add_51_79_groupi_n_2172 ,csa_tree_add_51_79_groupi_n_259);
  or csa_tree_add_51_79_groupi_g41974(csa_tree_add_51_79_groupi_n_4103 ,csa_tree_add_51_79_groupi_n_2028 ,csa_tree_add_51_79_groupi_n_900);
  or csa_tree_add_51_79_groupi_g41975(csa_tree_add_51_79_groupi_n_4102 ,csa_tree_add_51_79_groupi_n_2631 ,csa_tree_add_51_79_groupi_n_927);
  or csa_tree_add_51_79_groupi_g41976(csa_tree_add_51_79_groupi_n_4101 ,csa_tree_add_51_79_groupi_n_2882 ,csa_tree_add_51_79_groupi_n_217);
  or csa_tree_add_51_79_groupi_g41977(csa_tree_add_51_79_groupi_n_4100 ,csa_tree_add_51_79_groupi_n_2580 ,csa_tree_add_51_79_groupi_n_924);
  or csa_tree_add_51_79_groupi_g41978(csa_tree_add_51_79_groupi_n_4099 ,csa_tree_add_51_79_groupi_n_2700 ,csa_tree_add_51_79_groupi_n_325);
  or csa_tree_add_51_79_groupi_g41979(csa_tree_add_51_79_groupi_n_4098 ,csa_tree_add_51_79_groupi_n_2685 ,csa_tree_add_51_79_groupi_n_906);
  or csa_tree_add_51_79_groupi_g41980(csa_tree_add_51_79_groupi_n_4097 ,csa_tree_add_51_79_groupi_n_2697 ,csa_tree_add_51_79_groupi_n_1056);
  or csa_tree_add_51_79_groupi_g41981(csa_tree_add_51_79_groupi_n_4096 ,csa_tree_add_51_79_groupi_n_2085 ,csa_tree_add_51_79_groupi_n_391);
  or csa_tree_add_51_79_groupi_g41982(csa_tree_add_51_79_groupi_n_4095 ,csa_tree_add_51_79_groupi_n_2881 ,csa_tree_add_51_79_groupi_n_193);
  or csa_tree_add_51_79_groupi_g41983(csa_tree_add_51_79_groupi_n_4094 ,csa_tree_add_51_79_groupi_n_2698 ,csa_tree_add_51_79_groupi_n_132);
  or csa_tree_add_51_79_groupi_g41984(csa_tree_add_51_79_groupi_n_4093 ,csa_tree_add_51_79_groupi_n_2843 ,csa_tree_add_51_79_groupi_n_223);
  or csa_tree_add_51_79_groupi_g41985(csa_tree_add_51_79_groupi_n_4092 ,csa_tree_add_51_79_groupi_n_2562 ,csa_tree_add_51_79_groupi_n_3007);
  or csa_tree_add_51_79_groupi_g41986(csa_tree_add_51_79_groupi_n_4091 ,csa_tree_add_51_79_groupi_n_2604 ,csa_tree_add_51_79_groupi_n_963);
  nor csa_tree_add_51_79_groupi_g41987(csa_tree_add_51_79_groupi_n_4090 ,csa_tree_add_51_79_groupi_n_3785 ,csa_tree_add_51_79_groupi_n_3827);
  or csa_tree_add_51_79_groupi_g41988(csa_tree_add_51_79_groupi_n_4089 ,csa_tree_add_51_79_groupi_n_2611 ,csa_tree_add_51_79_groupi_n_915);
  or csa_tree_add_51_79_groupi_g41989(csa_tree_add_51_79_groupi_n_4088 ,csa_tree_add_51_79_groupi_n_2650 ,csa_tree_add_51_79_groupi_n_67);
  or csa_tree_add_51_79_groupi_g41990(csa_tree_add_51_79_groupi_n_4087 ,csa_tree_add_51_79_groupi_n_2783 ,csa_tree_add_51_79_groupi_n_97);
  or csa_tree_add_51_79_groupi_g41991(csa_tree_add_51_79_groupi_n_4086 ,csa_tree_add_51_79_groupi_n_2740 ,csa_tree_add_51_79_groupi_n_55);
  or csa_tree_add_51_79_groupi_g41992(csa_tree_add_51_79_groupi_n_4085 ,csa_tree_add_51_79_groupi_n_2809 ,csa_tree_add_51_79_groupi_n_996);
  or csa_tree_add_51_79_groupi_g41993(csa_tree_add_51_79_groupi_n_4084 ,csa_tree_add_51_79_groupi_n_2600 ,csa_tree_add_51_79_groupi_n_999);
  or csa_tree_add_51_79_groupi_g41994(csa_tree_add_51_79_groupi_n_4083 ,csa_tree_add_51_79_groupi_n_2062 ,csa_tree_add_51_79_groupi_n_372);
  or csa_tree_add_51_79_groupi_g41995(csa_tree_add_51_79_groupi_n_4082 ,csa_tree_add_51_79_groupi_n_2612 ,csa_tree_add_51_79_groupi_n_1038);
  or csa_tree_add_51_79_groupi_g41996(csa_tree_add_51_79_groupi_n_4081 ,csa_tree_add_51_79_groupi_n_2747 ,csa_tree_add_51_79_groupi_n_972);
  or csa_tree_add_51_79_groupi_g41997(csa_tree_add_51_79_groupi_n_4080 ,csa_tree_add_51_79_groupi_n_3283 ,csa_tree_add_51_79_groupi_n_3299);
  or csa_tree_add_51_79_groupi_g41998(csa_tree_add_51_79_groupi_n_4079 ,csa_tree_add_51_79_groupi_n_2879 ,csa_tree_add_51_79_groupi_n_1062);
  or csa_tree_add_51_79_groupi_g41999(csa_tree_add_51_79_groupi_n_4078 ,csa_tree_add_51_79_groupi_n_2192 ,csa_tree_add_51_79_groupi_n_277);
  or csa_tree_add_51_79_groupi_g42000(csa_tree_add_51_79_groupi_n_4077 ,csa_tree_add_51_79_groupi_n_2738 ,csa_tree_add_51_79_groupi_n_930);
  and csa_tree_add_51_79_groupi_g42001(csa_tree_add_51_79_groupi_n_4076 ,csa_tree_add_51_79_groupi_n_3288 ,csa_tree_add_51_79_groupi_n_3236);
  or csa_tree_add_51_79_groupi_g42002(csa_tree_add_51_79_groupi_n_4075 ,csa_tree_add_51_79_groupi_n_2320 ,csa_tree_add_51_79_groupi_n_264);
  or csa_tree_add_51_79_groupi_g42003(csa_tree_add_51_79_groupi_n_4074 ,csa_tree_add_51_79_groupi_n_2817 ,csa_tree_add_51_79_groupi_n_990);
  or csa_tree_add_51_79_groupi_g42004(csa_tree_add_51_79_groupi_n_4073 ,csa_tree_add_51_79_groupi_n_2371 ,csa_tree_add_51_79_groupi_n_270);
  or csa_tree_add_51_79_groupi_g42005(csa_tree_add_51_79_groupi_n_4072 ,csa_tree_add_51_79_groupi_n_1905 ,csa_tree_add_51_79_groupi_n_282);
  or csa_tree_add_51_79_groupi_g42006(csa_tree_add_51_79_groupi_n_4071 ,csa_tree_add_51_79_groupi_n_2179 ,csa_tree_add_51_79_groupi_n_1008);
  or csa_tree_add_51_79_groupi_g42007(csa_tree_add_51_79_groupi_n_4070 ,csa_tree_add_51_79_groupi_n_1793 ,csa_tree_add_51_79_groupi_n_330);
  or csa_tree_add_51_79_groupi_g42008(csa_tree_add_51_79_groupi_n_4069 ,csa_tree_add_51_79_groupi_n_2336 ,csa_tree_add_51_79_groupi_n_312);
  or csa_tree_add_51_79_groupi_g42009(csa_tree_add_51_79_groupi_n_4068 ,csa_tree_add_51_79_groupi_n_2138 ,csa_tree_add_51_79_groupi_n_91);
  or csa_tree_add_51_79_groupi_g42010(csa_tree_add_51_79_groupi_n_4067 ,csa_tree_add_51_79_groupi_n_2334 ,csa_tree_add_51_79_groupi_n_360);
  or csa_tree_add_51_79_groupi_g42011(csa_tree_add_51_79_groupi_n_4066 ,csa_tree_add_51_79_groupi_n_2084 ,csa_tree_add_51_79_groupi_n_205);
  or csa_tree_add_51_79_groupi_g42012(csa_tree_add_51_79_groupi_n_4065 ,csa_tree_add_51_79_groupi_n_2717 ,csa_tree_add_51_79_groupi_n_987);
  or csa_tree_add_51_79_groupi_g42013(csa_tree_add_51_79_groupi_n_4064 ,csa_tree_add_51_79_groupi_n_2726 ,csa_tree_add_51_79_groupi_n_1020);
  or csa_tree_add_51_79_groupi_g42014(csa_tree_add_51_79_groupi_n_4063 ,csa_tree_add_51_79_groupi_n_2221 ,csa_tree_add_51_79_groupi_n_1044);
  nor csa_tree_add_51_79_groupi_g42015(csa_tree_add_51_79_groupi_n_4062 ,csa_tree_add_51_79_groupi_n_2560 ,csa_tree_add_51_79_groupi_n_3003);
  or csa_tree_add_51_79_groupi_g42016(csa_tree_add_51_79_groupi_n_4061 ,csa_tree_add_51_79_groupi_n_2162 ,csa_tree_add_51_79_groupi_n_73);
  or csa_tree_add_51_79_groupi_g42017(csa_tree_add_51_79_groupi_n_4060 ,csa_tree_add_51_79_groupi_n_3278 ,csa_tree_add_51_79_groupi_n_3777);
  or csa_tree_add_51_79_groupi_g42018(csa_tree_add_51_79_groupi_n_4059 ,csa_tree_add_51_79_groupi_n_2163 ,csa_tree_add_51_79_groupi_n_1035);
  and csa_tree_add_51_79_groupi_g42019(csa_tree_add_51_79_groupi_n_4058 ,csa_tree_add_51_79_groupi_n_3796 ,csa_tree_add_51_79_groupi_n_3244);
  nor csa_tree_add_51_79_groupi_g42020(csa_tree_add_51_79_groupi_n_4057 ,csa_tree_add_51_79_groupi_n_2147 ,csa_tree_add_51_79_groupi_n_1032);
  or csa_tree_add_51_79_groupi_g42021(csa_tree_add_51_79_groupi_n_4056 ,csa_tree_add_51_79_groupi_n_2215 ,csa_tree_add_51_79_groupi_n_1059);
  or csa_tree_add_51_79_groupi_g42022(csa_tree_add_51_79_groupi_n_4055 ,csa_tree_add_51_79_groupi_n_2148 ,csa_tree_add_51_79_groupi_n_367);
  or csa_tree_add_51_79_groupi_g42023(csa_tree_add_51_79_groupi_n_4054 ,csa_tree_add_51_79_groupi_n_2684 ,csa_tree_add_51_79_groupi_n_1047);
  or csa_tree_add_51_79_groupi_g42024(csa_tree_add_51_79_groupi_n_4053 ,csa_tree_add_51_79_groupi_n_1925 ,csa_tree_add_51_79_groupi_n_391);
  or csa_tree_add_51_79_groupi_g42025(csa_tree_add_51_79_groupi_n_4052 ,csa_tree_add_51_79_groupi_n_2209 ,csa_tree_add_51_79_groupi_n_1005);
  or csa_tree_add_51_79_groupi_g42026(csa_tree_add_51_79_groupi_n_4051 ,csa_tree_add_51_79_groupi_n_2634 ,csa_tree_add_51_79_groupi_n_276);
  or csa_tree_add_51_79_groupi_g42027(csa_tree_add_51_79_groupi_n_4050 ,csa_tree_add_51_79_groupi_n_2081 ,csa_tree_add_51_79_groupi_n_210);
  or csa_tree_add_51_79_groupi_g42028(csa_tree_add_51_79_groupi_n_4049 ,csa_tree_add_51_79_groupi_n_2791 ,csa_tree_add_51_79_groupi_n_1014);
  or csa_tree_add_51_79_groupi_g42029(csa_tree_add_51_79_groupi_n_4048 ,csa_tree_add_51_79_groupi_n_2344 ,csa_tree_add_51_79_groupi_n_306);
  and csa_tree_add_51_79_groupi_g42030(csa_tree_add_51_79_groupi_n_4047 ,csa_tree_add_51_79_groupi_n_3257 ,csa_tree_add_51_79_groupi_n_3294);
  or csa_tree_add_51_79_groupi_g42031(csa_tree_add_51_79_groupi_n_4046 ,csa_tree_add_51_79_groupi_n_2609 ,csa_tree_add_51_79_groupi_n_97);
  or csa_tree_add_51_79_groupi_g42032(csa_tree_add_51_79_groupi_n_4045 ,csa_tree_add_51_79_groupi_n_3206 ,csa_tree_add_51_79_groupi_n_3194);
  or csa_tree_add_51_79_groupi_g42033(csa_tree_add_51_79_groupi_n_4044 ,csa_tree_add_51_79_groupi_n_2086 ,csa_tree_add_51_79_groupi_n_1002);
  or csa_tree_add_51_79_groupi_g42034(csa_tree_add_51_79_groupi_n_4043 ,csa_tree_add_51_79_groupi_n_2173 ,csa_tree_add_51_79_groupi_n_90);
  nor csa_tree_add_51_79_groupi_g42035(csa_tree_add_51_79_groupi_n_4042 ,csa_tree_add_51_79_groupi_n_3284 ,csa_tree_add_51_79_groupi_n_3300);
  or csa_tree_add_51_79_groupi_g42036(csa_tree_add_51_79_groupi_n_4041 ,csa_tree_add_51_79_groupi_n_2030 ,csa_tree_add_51_79_groupi_n_151);
  or csa_tree_add_51_79_groupi_g42037(csa_tree_add_51_79_groupi_n_4040 ,csa_tree_add_51_79_groupi_n_2743 ,csa_tree_add_51_79_groupi_n_948);
  or csa_tree_add_51_79_groupi_g42038(csa_tree_add_51_79_groupi_n_4039 ,csa_tree_add_51_79_groupi_n_2180 ,csa_tree_add_51_79_groupi_n_46);
  or csa_tree_add_51_79_groupi_g42039(csa_tree_add_51_79_groupi_n_4038 ,csa_tree_add_51_79_groupi_n_2058 ,csa_tree_add_51_79_groupi_n_918);
  or csa_tree_add_51_79_groupi_g42040(csa_tree_add_51_79_groupi_n_4037 ,csa_tree_add_51_79_groupi_n_2052 ,csa_tree_add_51_79_groupi_n_957);
  or csa_tree_add_51_79_groupi_g42041(csa_tree_add_51_79_groupi_n_4036 ,csa_tree_add_51_79_groupi_n_2076 ,csa_tree_add_51_79_groupi_n_378);
  or csa_tree_add_51_79_groupi_g42042(csa_tree_add_51_79_groupi_n_4035 ,csa_tree_add_51_79_groupi_n_2177 ,csa_tree_add_51_79_groupi_n_897);
  or csa_tree_add_51_79_groupi_g42043(csa_tree_add_51_79_groupi_n_4034 ,csa_tree_add_51_79_groupi_n_2111 ,csa_tree_add_51_79_groupi_n_324);
  or csa_tree_add_51_79_groupi_g42044(csa_tree_add_51_79_groupi_n_4033 ,csa_tree_add_51_79_groupi_n_2367 ,csa_tree_add_51_79_groupi_n_1056);
  or csa_tree_add_51_79_groupi_g42045(csa_tree_add_51_79_groupi_n_4032 ,csa_tree_add_51_79_groupi_n_2043 ,csa_tree_add_51_79_groupi_n_1023);
  or csa_tree_add_51_79_groupi_g42046(csa_tree_add_51_79_groupi_n_4031 ,csa_tree_add_51_79_groupi_n_2071 ,csa_tree_add_51_79_groupi_n_120);
  or csa_tree_add_51_79_groupi_g42047(csa_tree_add_51_79_groupi_n_4030 ,csa_tree_add_51_79_groupi_n_2193 ,csa_tree_add_51_79_groupi_n_259);
  nor csa_tree_add_51_79_groupi_g42048(csa_tree_add_51_79_groupi_n_4029 ,csa_tree_add_51_79_groupi_n_3755 ,csa_tree_add_51_79_groupi_n_3249);
  or csa_tree_add_51_79_groupi_g42049(csa_tree_add_51_79_groupi_n_4028 ,csa_tree_add_51_79_groupi_n_2326 ,csa_tree_add_51_79_groupi_n_354);
  or csa_tree_add_51_79_groupi_g42050(csa_tree_add_51_79_groupi_n_4027 ,csa_tree_add_51_79_groupi_n_2618 ,csa_tree_add_51_79_groupi_n_186);
  or csa_tree_add_51_79_groupi_g42051(csa_tree_add_51_79_groupi_n_4026 ,csa_tree_add_51_79_groupi_n_2258 ,csa_tree_add_51_79_groupi_n_366);
  or csa_tree_add_51_79_groupi_g42052(csa_tree_add_51_79_groupi_n_4025 ,csa_tree_add_51_79_groupi_n_2699 ,csa_tree_add_51_79_groupi_n_115);
  or csa_tree_add_51_79_groupi_g42053(csa_tree_add_51_79_groupi_n_4024 ,csa_tree_add_51_79_groupi_n_2864 ,csa_tree_add_51_79_groupi_n_978);
  or csa_tree_add_51_79_groupi_g42054(csa_tree_add_51_79_groupi_n_4023 ,csa_tree_add_51_79_groupi_n_2075 ,csa_tree_add_51_79_groupi_n_204);
  or csa_tree_add_51_79_groupi_g42055(csa_tree_add_51_79_groupi_n_4022 ,csa_tree_add_51_79_groupi_n_2678 ,csa_tree_add_51_79_groupi_n_960);
  or csa_tree_add_51_79_groupi_g42056(csa_tree_add_51_79_groupi_n_4021 ,csa_tree_add_51_79_groupi_n_2751 ,csa_tree_add_51_79_groupi_n_181);
  or csa_tree_add_51_79_groupi_g42057(csa_tree_add_51_79_groupi_n_4020 ,csa_tree_add_51_79_groupi_n_2041 ,csa_tree_add_51_79_groupi_n_912);
  or csa_tree_add_51_79_groupi_g42058(csa_tree_add_51_79_groupi_n_4019 ,csa_tree_add_51_79_groupi_n_2064 ,csa_tree_add_51_79_groupi_n_174);
  or csa_tree_add_51_79_groupi_g42059(csa_tree_add_51_79_groupi_n_4018 ,csa_tree_add_51_79_groupi_n_2787 ,csa_tree_add_51_79_groupi_n_1026);
  and csa_tree_add_51_79_groupi_g42060(csa_tree_add_51_79_groupi_n_4017 ,csa_tree_add_51_79_groupi_n_3205 ,csa_tree_add_51_79_groupi_n_3277);
  or csa_tree_add_51_79_groupi_g42061(csa_tree_add_51_79_groupi_n_4016 ,csa_tree_add_51_79_groupi_n_3790 ,csa_tree_add_51_79_groupi_n_3781);
  and csa_tree_add_51_79_groupi_g42062(csa_tree_add_51_79_groupi_n_4015 ,csa_tree_add_51_79_groupi_n_3737 ,csa_tree_add_51_79_groupi_n_3243);
  or csa_tree_add_51_79_groupi_g42063(csa_tree_add_51_79_groupi_n_4014 ,csa_tree_add_51_79_groupi_n_2778 ,csa_tree_add_51_79_groupi_n_241);
  or csa_tree_add_51_79_groupi_g42064(csa_tree_add_51_79_groupi_n_4013 ,csa_tree_add_51_79_groupi_n_2592 ,csa_tree_add_51_79_groupi_n_301);
  or csa_tree_add_51_79_groupi_g42065(csa_tree_add_51_79_groupi_n_4012 ,csa_tree_add_51_79_groupi_n_1852 ,csa_tree_add_51_79_groupi_n_933);
  or csa_tree_add_51_79_groupi_g42066(csa_tree_add_51_79_groupi_n_4011 ,csa_tree_add_51_79_groupi_n_2307 ,csa_tree_add_51_79_groupi_n_216);
  or csa_tree_add_51_79_groupi_g42067(csa_tree_add_51_79_groupi_n_4010 ,csa_tree_add_51_79_groupi_n_2691 ,csa_tree_add_51_79_groupi_n_235);
  or csa_tree_add_51_79_groupi_g42068(csa_tree_add_51_79_groupi_n_4009 ,csa_tree_add_51_79_groupi_n_2095 ,csa_tree_add_51_79_groupi_n_924);
  or csa_tree_add_51_79_groupi_g42069(csa_tree_add_51_79_groupi_n_4008 ,csa_tree_add_51_79_groupi_n_2629 ,csa_tree_add_51_79_groupi_n_126);
  or csa_tree_add_51_79_groupi_g42070(csa_tree_add_51_79_groupi_n_4007 ,csa_tree_add_51_79_groupi_n_2247 ,csa_tree_add_51_79_groupi_n_1011);
  or csa_tree_add_51_79_groupi_g42071(csa_tree_add_51_79_groupi_n_4006 ,csa_tree_add_51_79_groupi_n_2804 ,csa_tree_add_51_79_groupi_n_1038);
  or csa_tree_add_51_79_groupi_g42072(csa_tree_add_51_79_groupi_n_4005 ,csa_tree_add_51_79_groupi_n_2736 ,csa_tree_add_51_79_groupi_n_969);
  or csa_tree_add_51_79_groupi_g42073(csa_tree_add_51_79_groupi_n_4004 ,csa_tree_add_51_79_groupi_n_2098 ,csa_tree_add_51_79_groupi_n_894);
  nor csa_tree_add_51_79_groupi_g42074(csa_tree_add_51_79_groupi_n_4003 ,csa_tree_add_51_79_groupi_n_2255 ,csa_tree_add_51_79_groupi_n_1044);
  or csa_tree_add_51_79_groupi_g42075(csa_tree_add_51_79_groupi_n_4002 ,csa_tree_add_51_79_groupi_n_2779 ,csa_tree_add_51_79_groupi_n_978);
  or csa_tree_add_51_79_groupi_g42076(csa_tree_add_51_79_groupi_n_4001 ,csa_tree_add_51_79_groupi_n_2602 ,csa_tree_add_51_79_groupi_n_396);
  or csa_tree_add_51_79_groupi_g42077(csa_tree_add_51_79_groupi_n_4000 ,csa_tree_add_51_79_groupi_n_2099 ,csa_tree_add_51_79_groupi_n_927);
  or csa_tree_add_51_79_groupi_g42078(csa_tree_add_51_79_groupi_n_3999 ,csa_tree_add_51_79_groupi_n_1814 ,csa_tree_add_51_79_groupi_n_939);
  or csa_tree_add_51_79_groupi_g42079(csa_tree_add_51_79_groupi_n_3998 ,csa_tree_add_51_79_groupi_n_2097 ,csa_tree_add_51_79_groupi_n_966);
  or csa_tree_add_51_79_groupi_g42080(csa_tree_add_51_79_groupi_n_3997 ,csa_tree_add_51_79_groupi_n_2102 ,csa_tree_add_51_79_groupi_n_1050);
  or csa_tree_add_51_79_groupi_g42081(csa_tree_add_51_79_groupi_n_3996 ,csa_tree_add_51_79_groupi_n_1823 ,csa_tree_add_51_79_groupi_n_1053);
  nor csa_tree_add_51_79_groupi_g42082(csa_tree_add_51_79_groupi_n_3995 ,csa_tree_add_51_79_groupi_n_2101 ,csa_tree_add_51_79_groupi_n_1065);
  or csa_tree_add_51_79_groupi_g42083(csa_tree_add_51_79_groupi_n_3994 ,csa_tree_add_51_79_groupi_n_2104 ,csa_tree_add_51_79_groupi_n_945);
  or csa_tree_add_51_79_groupi_g42084(csa_tree_add_51_79_groupi_n_3993 ,csa_tree_add_51_79_groupi_n_1818 ,csa_tree_add_51_79_groupi_n_294);
  or csa_tree_add_51_79_groupi_g42085(csa_tree_add_51_79_groupi_n_3992 ,csa_tree_add_51_79_groupi_n_1816 ,csa_tree_add_51_79_groupi_n_336);
  or csa_tree_add_51_79_groupi_g42086(csa_tree_add_51_79_groupi_n_3991 ,csa_tree_add_51_79_groupi_n_2675 ,csa_tree_add_51_79_groupi_n_84);
  or csa_tree_add_51_79_groupi_g42087(csa_tree_add_51_79_groupi_n_3990 ,csa_tree_add_51_79_groupi_n_2116 ,csa_tree_add_51_79_groupi_n_1017);
  or csa_tree_add_51_79_groupi_g42088(csa_tree_add_51_79_groupi_n_3989 ,csa_tree_add_51_79_groupi_n_2665 ,csa_tree_add_51_79_groupi_n_318);
  or csa_tree_add_51_79_groupi_g42089(csa_tree_add_51_79_groupi_n_3988 ,csa_tree_add_51_79_groupi_n_2806 ,csa_tree_add_51_79_groupi_n_416);
  nor csa_tree_add_51_79_groupi_g42090(csa_tree_add_51_79_groupi_n_3987 ,csa_tree_add_51_79_groupi_n_2107 ,csa_tree_add_51_79_groupi_n_1056);
  or csa_tree_add_51_79_groupi_g42091(csa_tree_add_51_79_groupi_n_3986 ,csa_tree_add_51_79_groupi_n_2832 ,csa_tree_add_51_79_groupi_n_891);
  and csa_tree_add_51_79_groupi_g42092(csa_tree_add_51_79_groupi_n_3985 ,csa_tree_add_51_79_groupi_n_3199 ,csa_tree_add_51_79_groupi_n_3298);
  or csa_tree_add_51_79_groupi_g42093(csa_tree_add_51_79_groupi_n_3984 ,csa_tree_add_51_79_groupi_n_2707 ,csa_tree_add_51_79_groupi_n_180);
  nor csa_tree_add_51_79_groupi_g42094(csa_tree_add_51_79_groupi_n_3983 ,csa_tree_add_51_79_groupi_n_2590 ,csa_tree_add_51_79_groupi_n_1062);
  or csa_tree_add_51_79_groupi_g42095(csa_tree_add_51_79_groupi_n_3982 ,csa_tree_add_51_79_groupi_n_2130 ,csa_tree_add_51_79_groupi_n_157);
  or csa_tree_add_51_79_groupi_g42096(csa_tree_add_51_79_groupi_n_3981 ,csa_tree_add_51_79_groupi_n_2144 ,csa_tree_add_51_79_groupi_n_402);
  or csa_tree_add_51_79_groupi_g42097(csa_tree_add_51_79_groupi_n_3980 ,csa_tree_add_51_79_groupi_n_2132 ,csa_tree_add_51_79_groupi_n_72);
  or csa_tree_add_51_79_groupi_g42098(csa_tree_add_51_79_groupi_n_3979 ,csa_tree_add_51_79_groupi_n_2261 ,csa_tree_add_51_79_groupi_n_78);
  or csa_tree_add_51_79_groupi_g42099(csa_tree_add_51_79_groupi_n_3978 ,csa_tree_add_51_79_groupi_n_2862 ,csa_tree_add_51_79_groupi_n_222);
  or csa_tree_add_51_79_groupi_g42100(csa_tree_add_51_79_groupi_n_3977 ,csa_tree_add_51_79_groupi_n_2749 ,csa_tree_add_51_79_groupi_n_144);
  or csa_tree_add_51_79_groupi_g42101(csa_tree_add_51_79_groupi_n_3976 ,csa_tree_add_51_79_groupi_n_2610 ,csa_tree_add_51_79_groupi_n_288);
  or csa_tree_add_51_79_groupi_g42102(csa_tree_add_51_79_groupi_n_3975 ,csa_tree_add_51_79_groupi_n_2143 ,csa_tree_add_51_79_groupi_n_1044);
  or csa_tree_add_51_79_groupi_g42103(csa_tree_add_51_79_groupi_n_3974 ,csa_tree_add_51_79_groupi_n_2640 ,csa_tree_add_51_79_groupi_n_903);
  and csa_tree_add_51_79_groupi_g42104(csa_tree_add_51_79_groupi_n_3973 ,csa_tree_add_51_79_groupi_n_3266 ,csa_tree_add_51_79_groupi_n_3263);
  or csa_tree_add_51_79_groupi_g42105(csa_tree_add_51_79_groupi_n_3972 ,csa_tree_add_51_79_groupi_n_2078 ,csa_tree_add_51_79_groupi_n_912);
  or csa_tree_add_51_79_groupi_g42106(csa_tree_add_51_79_groupi_n_3971 ,csa_tree_add_51_79_groupi_n_2127 ,csa_tree_add_51_79_groupi_n_963);
  or csa_tree_add_51_79_groupi_g42107(csa_tree_add_51_79_groupi_n_3970 ,csa_tree_add_51_79_groupi_n_1815 ,csa_tree_add_51_79_groupi_n_46);
  nor csa_tree_add_51_79_groupi_g42108(csa_tree_add_51_79_groupi_n_3969 ,csa_tree_add_51_79_groupi_n_2121 ,csa_tree_add_51_79_groupi_n_1026);
  or csa_tree_add_51_79_groupi_g42109(csa_tree_add_51_79_groupi_n_3968 ,csa_tree_add_51_79_groupi_n_2129 ,csa_tree_add_51_79_groupi_n_921);
  or csa_tree_add_51_79_groupi_g42110(csa_tree_add_51_79_groupi_n_3967 ,csa_tree_add_51_79_groupi_n_2204 ,csa_tree_add_51_79_groupi_n_1041);
  or csa_tree_add_51_79_groupi_g42111(csa_tree_add_51_79_groupi_n_3966 ,csa_tree_add_51_79_groupi_n_2702 ,csa_tree_add_51_79_groupi_n_1026);
  or csa_tree_add_51_79_groupi_g42112(csa_tree_add_51_79_groupi_n_3965 ,csa_tree_add_51_79_groupi_n_2716 ,csa_tree_add_51_79_groupi_n_948);
  or csa_tree_add_51_79_groupi_g42113(csa_tree_add_51_79_groupi_n_3964 ,csa_tree_add_51_79_groupi_n_2784 ,csa_tree_add_51_79_groupi_n_900);
  and csa_tree_add_51_79_groupi_g42114(csa_tree_add_51_79_groupi_n_3963 ,csa_tree_add_51_79_groupi_n_3245 ,csa_tree_add_51_79_groupi_n_3763);
  or csa_tree_add_51_79_groupi_g42115(csa_tree_add_51_79_groupi_n_3962 ,csa_tree_add_51_79_groupi_n_2733 ,csa_tree_add_51_79_groupi_n_930);
  or csa_tree_add_51_79_groupi_g42116(csa_tree_add_51_79_groupi_n_3961 ,csa_tree_add_51_79_groupi_n_2744 ,csa_tree_add_51_79_groupi_n_987);
  or csa_tree_add_51_79_groupi_g42117(csa_tree_add_51_79_groupi_n_3960 ,csa_tree_add_51_79_groupi_n_2139 ,csa_tree_add_51_79_groupi_n_1023);
  or csa_tree_add_51_79_groupi_g42118(csa_tree_add_51_79_groupi_n_3959 ,csa_tree_add_51_79_groupi_n_2140 ,csa_tree_add_51_79_groupi_n_996);
  or csa_tree_add_51_79_groupi_g42119(csa_tree_add_51_79_groupi_n_3958 ,csa_tree_add_51_79_groupi_n_1799 ,csa_tree_add_51_79_groupi_n_247);
  or csa_tree_add_51_79_groupi_g42120(csa_tree_add_51_79_groupi_n_3957 ,csa_tree_add_51_79_groupi_n_2782 ,csa_tree_add_51_79_groupi_n_1020);
  or csa_tree_add_51_79_groupi_g42121(csa_tree_add_51_79_groupi_n_3956 ,csa_tree_add_51_79_groupi_n_1797 ,csa_tree_add_51_79_groupi_n_897);
  or csa_tree_add_51_79_groupi_g42122(csa_tree_add_51_79_groupi_n_3955 ,csa_tree_add_51_79_groupi_n_2369 ,csa_tree_add_51_79_groupi_n_975);
  or csa_tree_add_51_79_groupi_g42123(csa_tree_add_51_79_groupi_n_3954 ,csa_tree_add_51_79_groupi_n_2274 ,csa_tree_add_51_79_groupi_n_972);
  or csa_tree_add_51_79_groupi_g42124(csa_tree_add_51_79_groupi_n_3953 ,csa_tree_add_51_79_groupi_n_2141 ,csa_tree_add_51_79_groupi_n_300);
  or csa_tree_add_51_79_groupi_g42125(csa_tree_add_51_79_groupi_n_3952 ,csa_tree_add_51_79_groupi_n_2853 ,csa_tree_add_51_79_groupi_n_162);
  or csa_tree_add_51_79_groupi_g42126(csa_tree_add_51_79_groupi_n_3951 ,csa_tree_add_51_79_groupi_n_2883 ,csa_tree_add_51_79_groupi_n_936);
  or csa_tree_add_51_79_groupi_g42127(csa_tree_add_51_79_groupi_n_3950 ,csa_tree_add_51_79_groupi_n_2265 ,csa_tree_add_51_79_groupi_n_258);
  or csa_tree_add_51_79_groupi_g42128(csa_tree_add_51_79_groupi_n_3949 ,csa_tree_add_51_79_groupi_n_3307 ,csa_tree_add_51_79_groupi_n_3274);
  and csa_tree_add_51_79_groupi_g42129(csa_tree_add_51_79_groupi_n_3948 ,csa_tree_add_51_79_groupi_n_3307 ,csa_tree_add_51_79_groupi_n_3274);
  or csa_tree_add_51_79_groupi_g42130(csa_tree_add_51_79_groupi_n_3947 ,csa_tree_add_51_79_groupi_n_3289 ,csa_tree_add_51_79_groupi_n_3202);
  or csa_tree_add_51_79_groupi_g42131(csa_tree_add_51_79_groupi_n_3946 ,csa_tree_add_51_79_groupi_n_2142 ,csa_tree_add_51_79_groupi_n_975);
  and csa_tree_add_51_79_groupi_g42132(csa_tree_add_51_79_groupi_n_3945 ,csa_tree_add_51_79_groupi_n_3289 ,csa_tree_add_51_79_groupi_n_3202);
  and csa_tree_add_51_79_groupi_g42133(csa_tree_add_51_79_groupi_n_3944 ,csa_tree_add_51_79_groupi_n_3225 ,csa_tree_add_51_79_groupi_n_3253);
  or csa_tree_add_51_79_groupi_g42134(csa_tree_add_51_79_groupi_n_3943 ,csa_tree_add_51_79_groupi_n_2185 ,csa_tree_add_51_79_groupi_n_115);
  or csa_tree_add_51_79_groupi_g42135(csa_tree_add_51_79_groupi_n_3942 ,csa_tree_add_51_79_groupi_n_3212 ,csa_tree_add_51_79_groupi_n_3749);
  or csa_tree_add_51_79_groupi_g42136(csa_tree_add_51_79_groupi_n_3941 ,csa_tree_add_51_79_groupi_n_2718 ,csa_tree_add_51_79_groupi_n_342);
  or csa_tree_add_51_79_groupi_g42137(csa_tree_add_51_79_groupi_n_3940 ,csa_tree_add_51_79_groupi_n_2154 ,csa_tree_add_51_79_groupi_n_1053);
  or csa_tree_add_51_79_groupi_g42138(csa_tree_add_51_79_groupi_n_3939 ,csa_tree_add_51_79_groupi_n_1803 ,csa_tree_add_51_79_groupi_n_253);
  or csa_tree_add_51_79_groupi_g42139(csa_tree_add_51_79_groupi_n_3938 ,csa_tree_add_51_79_groupi_n_2240 ,csa_tree_add_51_79_groupi_n_96);
  or csa_tree_add_51_79_groupi_g42140(csa_tree_add_51_79_groupi_n_3937 ,csa_tree_add_51_79_groupi_n_2706 ,csa_tree_add_51_79_groupi_n_235);
  or csa_tree_add_51_79_groupi_g42141(csa_tree_add_51_79_groupi_n_3936 ,csa_tree_add_51_79_groupi_n_2040 ,csa_tree_add_51_79_groupi_n_993);
  and csa_tree_add_51_79_groupi_g42142(csa_tree_add_51_79_groupi_n_3935 ,csa_tree_add_51_79_groupi_n_3753 ,csa_tree_add_51_79_groupi_n_3297);
  or csa_tree_add_51_79_groupi_g42143(csa_tree_add_51_79_groupi_n_3934 ,csa_tree_add_51_79_groupi_n_1821 ,csa_tree_add_51_79_groupi_n_1059);
  or csa_tree_add_51_79_groupi_g42144(csa_tree_add_51_79_groupi_n_3933 ,csa_tree_add_51_79_groupi_n_2250 ,csa_tree_add_51_79_groupi_n_1065);
  or csa_tree_add_51_79_groupi_g42145(csa_tree_add_51_79_groupi_n_3932 ,csa_tree_add_51_79_groupi_n_2252 ,csa_tree_add_51_79_groupi_n_1014);
  nor csa_tree_add_51_79_groupi_g42146(csa_tree_add_51_79_groupi_n_3931 ,csa_tree_add_51_79_groupi_n_2257 ,csa_tree_add_51_79_groupi_n_1059);
  nor csa_tree_add_51_79_groupi_g42147(csa_tree_add_51_79_groupi_n_3930 ,csa_tree_add_51_79_groupi_n_3213 ,csa_tree_add_51_79_groupi_n_3750);
  or csa_tree_add_51_79_groupi_g42148(csa_tree_add_51_79_groupi_n_3929 ,csa_tree_add_51_79_groupi_n_2293 ,csa_tree_add_51_79_groupi_n_918);
  or csa_tree_add_51_79_groupi_g42149(csa_tree_add_51_79_groupi_n_3928 ,csa_tree_add_51_79_groupi_n_3753 ,csa_tree_add_51_79_groupi_n_3297);
  or csa_tree_add_51_79_groupi_g42150(csa_tree_add_51_79_groupi_n_3927 ,csa_tree_add_51_79_groupi_n_2295 ,csa_tree_add_51_79_groupi_n_192);
  or csa_tree_add_51_79_groupi_g42151(csa_tree_add_51_79_groupi_n_3926 ,csa_tree_add_51_79_groupi_n_2275 ,csa_tree_add_51_79_groupi_n_1056);
  or csa_tree_add_51_79_groupi_g42152(csa_tree_add_51_79_groupi_n_3925 ,csa_tree_add_51_79_groupi_n_2135 ,csa_tree_add_51_79_groupi_n_1041);
  or csa_tree_add_51_79_groupi_g42153(csa_tree_add_51_79_groupi_n_3924 ,csa_tree_add_51_79_groupi_n_2315 ,csa_tree_add_51_79_groupi_n_942);
  or csa_tree_add_51_79_groupi_g42154(csa_tree_add_51_79_groupi_n_3923 ,csa_tree_add_51_79_groupi_n_2063 ,csa_tree_add_51_79_groupi_n_1029);
  nor csa_tree_add_51_79_groupi_g42155(csa_tree_add_51_79_groupi_n_3922 ,csa_tree_add_51_79_groupi_n_2264 ,csa_tree_add_51_79_groupi_n_1017);
  or csa_tree_add_51_79_groupi_g42156(csa_tree_add_51_79_groupi_n_3921 ,csa_tree_add_51_79_groupi_n_2316 ,csa_tree_add_51_79_groupi_n_915);
  nor csa_tree_add_51_79_groupi_g42157(csa_tree_add_51_79_groupi_n_3920 ,csa_tree_add_51_79_groupi_n_2282 ,csa_tree_add_51_79_groupi_n_1023);
  or csa_tree_add_51_79_groupi_g42158(csa_tree_add_51_79_groupi_n_3919 ,csa_tree_add_51_79_groupi_n_2303 ,csa_tree_add_51_79_groupi_n_957);
  or csa_tree_add_51_79_groupi_g42159(csa_tree_add_51_79_groupi_n_3918 ,csa_tree_add_51_79_groupi_n_2249 ,csa_tree_add_51_79_groupi_n_966);
  or csa_tree_add_51_79_groupi_g42160(csa_tree_add_51_79_groupi_n_3917 ,csa_tree_add_51_79_groupi_n_2317 ,csa_tree_add_51_79_groupi_n_981);
  or csa_tree_add_51_79_groupi_g42161(csa_tree_add_51_79_groupi_n_3916 ,csa_tree_add_51_79_groupi_n_2314 ,csa_tree_add_51_79_groupi_n_906);
  or csa_tree_add_51_79_groupi_g42162(csa_tree_add_51_79_groupi_n_3915 ,csa_tree_add_51_79_groupi_n_2313 ,csa_tree_add_51_79_groupi_n_1047);
  or csa_tree_add_51_79_groupi_g42163(csa_tree_add_51_79_groupi_n_3914 ,csa_tree_add_51_79_groupi_n_2701 ,csa_tree_add_51_79_groupi_n_168);
  or csa_tree_add_51_79_groupi_g42164(csa_tree_add_51_79_groupi_n_3913 ,csa_tree_add_51_79_groupi_n_2093 ,csa_tree_add_51_79_groupi_n_1017);
  or csa_tree_add_51_79_groupi_g42165(csa_tree_add_51_79_groupi_n_3912 ,csa_tree_add_51_79_groupi_n_2134 ,csa_tree_add_51_79_groupi_n_1035);
  or csa_tree_add_51_79_groupi_g42166(csa_tree_add_51_79_groupi_n_3911 ,csa_tree_add_51_79_groupi_n_2217 ,csa_tree_add_51_79_groupi_n_1032);
  or csa_tree_add_51_79_groupi_g42167(csa_tree_add_51_79_groupi_n_3910 ,csa_tree_add_51_79_groupi_n_3796 ,csa_tree_add_51_79_groupi_n_3244);
  or csa_tree_add_51_79_groupi_g42168(csa_tree_add_51_79_groupi_n_3909 ,csa_tree_add_51_79_groupi_n_2276 ,csa_tree_add_51_79_groupi_n_951);
  or csa_tree_add_51_79_groupi_g42169(csa_tree_add_51_79_groupi_n_3908 ,csa_tree_add_51_79_groupi_n_2296 ,csa_tree_add_51_79_groupi_n_921);
  and csa_tree_add_51_79_groupi_g42170(csa_tree_add_51_79_groupi_n_3907 ,csa_tree_add_51_79_groupi_n_3198 ,csa_tree_add_51_79_groupi_n_3201);
  or csa_tree_add_51_79_groupi_g42171(csa_tree_add_51_79_groupi_n_3906 ,csa_tree_add_51_79_groupi_n_2031 ,csa_tree_add_51_79_groupi_n_138);
  or csa_tree_add_51_79_groupi_g42172(csa_tree_add_51_79_groupi_n_3905 ,csa_tree_add_51_79_groupi_n_1863 ,csa_tree_add_51_79_groupi_n_234);
  or csa_tree_add_51_79_groupi_g42173(csa_tree_add_51_79_groupi_n_3904 ,csa_tree_add_51_79_groupi_n_2703 ,csa_tree_add_51_79_groupi_n_981);
  or csa_tree_add_51_79_groupi_g42174(csa_tree_add_51_79_groupi_n_3903 ,csa_tree_add_51_79_groupi_n_2774 ,csa_tree_add_51_79_groupi_n_1002);
  or csa_tree_add_51_79_groupi_g42175(csa_tree_add_51_79_groupi_n_3902 ,csa_tree_add_51_79_groupi_n_1822 ,csa_tree_add_51_79_groupi_n_1005);
  or csa_tree_add_51_79_groupi_g42176(csa_tree_add_51_79_groupi_n_3901 ,csa_tree_add_51_79_groupi_n_2306 ,csa_tree_add_51_79_groupi_n_954);
  or csa_tree_add_51_79_groupi_g42177(csa_tree_add_51_79_groupi_n_3900 ,csa_tree_add_51_79_groupi_n_2649 ,csa_tree_add_51_79_groupi_n_969);
  or csa_tree_add_51_79_groupi_g42178(csa_tree_add_51_79_groupi_n_3899 ,csa_tree_add_51_79_groupi_n_2272 ,csa_tree_add_51_79_groupi_n_939);
  or csa_tree_add_51_79_groupi_g42179(csa_tree_add_51_79_groupi_n_3898 ,csa_tree_add_51_79_groupi_n_1817 ,csa_tree_add_51_79_groupi_n_1008);
  or csa_tree_add_51_79_groupi_g42180(csa_tree_add_51_79_groupi_n_3897 ,csa_tree_add_51_79_groupi_n_2302 ,csa_tree_add_51_79_groupi_n_999);
  or csa_tree_add_51_79_groupi_g42181(csa_tree_add_51_79_groupi_n_3896 ,csa_tree_add_51_79_groupi_n_2301 ,csa_tree_add_51_79_groupi_n_1062);
  or csa_tree_add_51_79_groupi_g42182(csa_tree_add_51_79_groupi_n_3895 ,csa_tree_add_51_79_groupi_n_2015 ,csa_tree_add_51_79_groupi_n_960);
  or csa_tree_add_51_79_groupi_g42183(csa_tree_add_51_79_groupi_n_3894 ,csa_tree_add_51_79_groupi_n_2112 ,csa_tree_add_51_79_groupi_n_984);
  nor csa_tree_add_51_79_groupi_g42184(csa_tree_add_51_79_groupi_n_3893 ,csa_tree_add_51_79_groupi_n_2024 ,csa_tree_add_51_79_groupi_n_1020);
  or csa_tree_add_51_79_groupi_g42185(csa_tree_add_51_79_groupi_n_3892 ,csa_tree_add_51_79_groupi_n_2605 ,csa_tree_add_51_79_groupi_n_390);
  or csa_tree_add_51_79_groupi_g42186(csa_tree_add_51_79_groupi_n_3891 ,csa_tree_add_51_79_groupi_n_2294 ,csa_tree_add_51_79_groupi_n_114);
  or csa_tree_add_51_79_groupi_g42187(csa_tree_add_51_79_groupi_n_3890 ,csa_tree_add_51_79_groupi_n_1071 ,csa_tree_add_51_79_groupi_n_3282);
  or csa_tree_add_51_79_groupi_g42188(csa_tree_add_51_79_groupi_n_3889 ,csa_tree_add_51_79_groupi_n_2297 ,csa_tree_add_51_79_groupi_n_933);
  or csa_tree_add_51_79_groupi_g42189(csa_tree_add_51_79_groupi_n_3888 ,csa_tree_add_51_79_groupi_n_2807 ,csa_tree_add_51_79_groupi_n_909);
  or csa_tree_add_51_79_groupi_g42190(csa_tree_add_51_79_groupi_n_3887 ,csa_tree_add_51_79_groupi_n_2289 ,csa_tree_add_51_79_groupi_n_951);
  or csa_tree_add_51_79_groupi_g42191(csa_tree_add_51_79_groupi_n_3886 ,csa_tree_add_51_79_groupi_n_2287 ,csa_tree_add_51_79_groupi_n_999);
  or csa_tree_add_51_79_groupi_g42192(csa_tree_add_51_79_groupi_n_3885 ,csa_tree_add_51_79_groupi_n_1806 ,csa_tree_add_51_79_groupi_n_1011);
  or csa_tree_add_51_79_groupi_g42193(csa_tree_add_51_79_groupi_n_3884 ,csa_tree_add_51_79_groupi_n_2060 ,csa_tree_add_51_79_groupi_n_891);
  or csa_tree_add_51_79_groupi_g42194(csa_tree_add_51_79_groupi_n_3883 ,csa_tree_add_51_79_groupi_n_2206 ,csa_tree_add_51_79_groupi_n_1044);
  or csa_tree_add_51_79_groupi_g42195(csa_tree_add_51_79_groupi_n_3882 ,csa_tree_add_51_79_groupi_n_3245 ,csa_tree_add_51_79_groupi_n_3763);
  or csa_tree_add_51_79_groupi_g42196(csa_tree_add_51_79_groupi_n_3881 ,csa_tree_add_51_79_groupi_n_2288 ,csa_tree_add_51_79_groupi_n_990);
  and csa_tree_add_51_79_groupi_g42197(csa_tree_add_51_79_groupi_n_4305 ,csa_tree_add_51_79_groupi_n_3776 ,csa_tree_add_51_79_groupi_n_3744);
  and csa_tree_add_51_79_groupi_g42198(csa_tree_add_51_79_groupi_n_4304 ,csa_tree_add_51_79_groupi_n_3247 ,csa_tree_add_51_79_groupi_n_3743);
  or csa_tree_add_51_79_groupi_g42199(csa_tree_add_51_79_groupi_n_4303 ,csa_tree_add_51_79_groupi_n_3247 ,csa_tree_add_51_79_groupi_n_3743);
  xnor csa_tree_add_51_79_groupi_g42200(csa_tree_add_51_79_groupi_n_3880 ,csa_tree_add_51_79_groupi_n_2558 ,csa_tree_add_51_79_groupi_n_2552);
  xnor csa_tree_add_51_79_groupi_g42201(csa_tree_add_51_79_groupi_n_3879 ,csa_tree_add_51_79_groupi_n_2553 ,csa_tree_add_51_79_groupi_n_2554);
  xnor csa_tree_add_51_79_groupi_g42202(csa_tree_add_51_79_groupi_n_3878 ,csa_tree_add_51_79_groupi_n_2557 ,csa_tree_add_51_79_groupi_n_2556);
  or csa_tree_add_51_79_groupi_g42203(csa_tree_add_51_79_groupi_n_4302 ,csa_tree_add_51_79_groupi_n_3250 ,csa_tree_add_51_79_groupi_n_3786);
  xnor csa_tree_add_51_79_groupi_g42204(csa_tree_add_51_79_groupi_n_3877 ,csa_tree_add_51_79_groupi_n_2546 ,csa_tree_add_51_79_groupi_n_2566);
  xnor csa_tree_add_51_79_groupi_g42205(csa_tree_add_51_79_groupi_n_3876 ,csa_tree_add_51_79_groupi_n_2541 ,csa_tree_add_51_79_groupi_n_2550);
  xnor csa_tree_add_51_79_groupi_g42206(csa_tree_add_51_79_groupi_n_3875 ,csa_tree_add_51_79_groupi_n_2547 ,csa_tree_add_51_79_groupi_n_2559);
  xnor csa_tree_add_51_79_groupi_g42207(csa_tree_add_51_79_groupi_n_3874 ,csa_tree_add_51_79_groupi_n_2551 ,csa_tree_add_51_79_groupi_n_2565);
  xor csa_tree_add_51_79_groupi_g42208(csa_tree_add_51_79_groupi_n_3873 ,csa_tree_add_51_79_groupi_n_2555 ,csa_tree_add_51_79_groupi_n_2570);
  or csa_tree_add_51_79_groupi_g42209(csa_tree_add_51_79_groupi_n_4301 ,csa_tree_add_51_79_groupi_n_1532 ,csa_tree_add_51_79_groupi_n_3069);
  or csa_tree_add_51_79_groupi_g42210(csa_tree_add_51_79_groupi_n_4300 ,csa_tree_add_51_79_groupi_n_1555 ,csa_tree_add_51_79_groupi_n_2896);
  or csa_tree_add_51_79_groupi_g42211(csa_tree_add_51_79_groupi_n_4299 ,csa_tree_add_51_79_groupi_n_1544 ,csa_tree_add_51_79_groupi_n_3475);
  or csa_tree_add_51_79_groupi_g42212(csa_tree_add_51_79_groupi_n_4298 ,csa_tree_add_51_79_groupi_n_1613 ,csa_tree_add_51_79_groupi_n_3469);
  or csa_tree_add_51_79_groupi_g42213(csa_tree_add_51_79_groupi_n_4297 ,csa_tree_add_51_79_groupi_n_1546 ,csa_tree_add_51_79_groupi_n_3466);
  or csa_tree_add_51_79_groupi_g42214(csa_tree_add_51_79_groupi_n_4296 ,csa_tree_add_51_79_groupi_n_1609 ,csa_tree_add_51_79_groupi_n_3566);
  or csa_tree_add_51_79_groupi_g42215(csa_tree_add_51_79_groupi_n_4295 ,csa_tree_add_51_79_groupi_n_1535 ,csa_tree_add_51_79_groupi_n_3548);
  or csa_tree_add_51_79_groupi_g42216(csa_tree_add_51_79_groupi_n_4294 ,csa_tree_add_51_79_groupi_n_1616 ,csa_tree_add_51_79_groupi_n_3157);
  or csa_tree_add_51_79_groupi_g42217(csa_tree_add_51_79_groupi_n_4293 ,csa_tree_add_51_79_groupi_n_1534 ,csa_tree_add_51_79_groupi_n_3053);
  or csa_tree_add_51_79_groupi_g42218(csa_tree_add_51_79_groupi_n_4292 ,csa_tree_add_51_79_groupi_n_1621 ,csa_tree_add_51_79_groupi_n_3042);
  or csa_tree_add_51_79_groupi_g42219(csa_tree_add_51_79_groupi_n_4291 ,csa_tree_add_51_79_groupi_n_1549 ,csa_tree_add_51_79_groupi_n_3406);
  or csa_tree_add_51_79_groupi_g42220(csa_tree_add_51_79_groupi_n_4290 ,csa_tree_add_51_79_groupi_n_1618 ,csa_tree_add_51_79_groupi_n_3036);
  or csa_tree_add_51_79_groupi_g42221(csa_tree_add_51_79_groupi_n_4289 ,csa_tree_add_51_79_groupi_n_1551 ,csa_tree_add_51_79_groupi_n_3393);
  or csa_tree_add_51_79_groupi_g42222(csa_tree_add_51_79_groupi_n_4288 ,csa_tree_add_51_79_groupi_n_1615 ,csa_tree_add_51_79_groupi_n_3070);
  or csa_tree_add_51_79_groupi_g42223(csa_tree_add_51_79_groupi_n_4287 ,csa_tree_add_51_79_groupi_n_1624 ,csa_tree_add_51_79_groupi_n_3575);
  or csa_tree_add_51_79_groupi_g42224(csa_tree_add_51_79_groupi_n_4286 ,csa_tree_add_51_79_groupi_n_1623 ,csa_tree_add_51_79_groupi_n_3407);
  and csa_tree_add_51_79_groupi_g42225(csa_tree_add_51_79_groupi_n_4285 ,csa_tree_add_51_79_groupi_n_2393 ,csa_tree_add_51_79_groupi_n_3424);
  and csa_tree_add_51_79_groupi_g42226(csa_tree_add_51_79_groupi_n_4284 ,csa_tree_add_51_79_groupi_n_3273 ,csa_tree_add_51_79_groupi_n_3736);
  or csa_tree_add_51_79_groupi_g42227(csa_tree_add_51_79_groupi_n_4283 ,csa_tree_add_51_79_groupi_n_1620 ,csa_tree_add_51_79_groupi_n_3688);
  or csa_tree_add_51_79_groupi_g42228(csa_tree_add_51_79_groupi_n_4280 ,csa_tree_add_51_79_groupi_n_1619 ,csa_tree_add_51_79_groupi_n_3381);
  or csa_tree_add_51_79_groupi_g42229(csa_tree_add_51_79_groupi_n_4279 ,csa_tree_add_51_79_groupi_n_1598 ,csa_tree_add_51_79_groupi_n_3382);
  or csa_tree_add_51_79_groupi_g42230(csa_tree_add_51_79_groupi_n_4276 ,csa_tree_add_51_79_groupi_n_1552 ,csa_tree_add_51_79_groupi_n_3067);
  or csa_tree_add_51_79_groupi_g42231(csa_tree_add_51_79_groupi_n_4275 ,csa_tree_add_51_79_groupi_n_1531 ,csa_tree_add_51_79_groupi_n_3481);
  or csa_tree_add_51_79_groupi_g42232(csa_tree_add_51_79_groupi_n_4273 ,csa_tree_add_51_79_groupi_n_1533 ,csa_tree_add_51_79_groupi_n_3130);
  or csa_tree_add_51_79_groupi_g42233(csa_tree_add_51_79_groupi_n_4271 ,csa_tree_add_51_79_groupi_n_1605 ,csa_tree_add_51_79_groupi_n_3511);
  or csa_tree_add_51_79_groupi_g42234(csa_tree_add_51_79_groupi_n_4268 ,csa_tree_add_51_79_groupi_n_1538 ,csa_tree_add_51_79_groupi_n_3493);
  or csa_tree_add_51_79_groupi_g42235(csa_tree_add_51_79_groupi_n_4267 ,csa_tree_add_51_79_groupi_n_1626 ,csa_tree_add_51_79_groupi_n_3463);
  or csa_tree_add_51_79_groupi_g42236(csa_tree_add_51_79_groupi_n_4265 ,csa_tree_add_51_79_groupi_n_1548 ,csa_tree_add_51_79_groupi_n_3477);
  or csa_tree_add_51_79_groupi_g42237(csa_tree_add_51_79_groupi_n_4264 ,csa_tree_add_51_79_groupi_n_1596 ,csa_tree_add_51_79_groupi_n_3476);
  or csa_tree_add_51_79_groupi_g42238(csa_tree_add_51_79_groupi_n_4262 ,csa_tree_add_51_79_groupi_n_1611 ,csa_tree_add_51_79_groupi_n_3088);
  or csa_tree_add_51_79_groupi_g42239(csa_tree_add_51_79_groupi_n_4260 ,csa_tree_add_51_79_groupi_n_1627 ,csa_tree_add_51_79_groupi_n_3046);
  or csa_tree_add_51_79_groupi_g42240(csa_tree_add_51_79_groupi_n_4258 ,csa_tree_add_51_79_groupi_n_1541 ,csa_tree_add_51_79_groupi_n_3074);
  or csa_tree_add_51_79_groupi_g42241(csa_tree_add_51_79_groupi_n_4257 ,csa_tree_add_51_79_groupi_n_1603 ,csa_tree_add_51_79_groupi_n_3142);
  or csa_tree_add_51_79_groupi_g42242(csa_tree_add_51_79_groupi_n_4254 ,csa_tree_add_51_79_groupi_n_1608 ,csa_tree_add_51_79_groupi_n_3572);
  or csa_tree_add_51_79_groupi_g42243(csa_tree_add_51_79_groupi_n_4253 ,csa_tree_add_51_79_groupi_n_1600 ,csa_tree_add_51_79_groupi_n_3049);
  or csa_tree_add_51_79_groupi_g42244(csa_tree_add_51_79_groupi_n_4250 ,csa_tree_add_51_79_groupi_n_1604 ,csa_tree_add_51_79_groupi_n_3472);
  or csa_tree_add_51_79_groupi_g42245(csa_tree_add_51_79_groupi_n_4249 ,csa_tree_add_51_79_groupi_n_1543 ,csa_tree_add_51_79_groupi_n_3471);
  or csa_tree_add_51_79_groupi_g42246(csa_tree_add_51_79_groupi_n_4246 ,csa_tree_add_51_79_groupi_n_1545 ,csa_tree_add_51_79_groupi_n_3408);
  or csa_tree_add_51_79_groupi_g42247(csa_tree_add_51_79_groupi_n_4244 ,csa_tree_add_51_79_groupi_n_1597 ,csa_tree_add_51_79_groupi_n_3066);
  or csa_tree_add_51_79_groupi_g42248(csa_tree_add_51_79_groupi_n_4243 ,csa_tree_add_51_79_groupi_n_1556 ,csa_tree_add_51_79_groupi_n_2898);
  or csa_tree_add_51_79_groupi_g42249(csa_tree_add_51_79_groupi_n_4241 ,csa_tree_add_51_79_groupi_n_1602 ,csa_tree_add_51_79_groupi_n_3031);
  or csa_tree_add_51_79_groupi_g42250(csa_tree_add_51_79_groupi_n_4240 ,csa_tree_add_51_79_groupi_n_1614 ,csa_tree_add_51_79_groupi_n_2980);
  or csa_tree_add_51_79_groupi_g42251(csa_tree_add_51_79_groupi_n_4237 ,csa_tree_add_51_79_groupi_n_1536 ,csa_tree_add_51_79_groupi_n_3571);
  or csa_tree_add_51_79_groupi_g42252(csa_tree_add_51_79_groupi_n_4236 ,csa_tree_add_51_79_groupi_n_1625 ,csa_tree_add_51_79_groupi_n_3062);
  or csa_tree_add_51_79_groupi_g42253(csa_tree_add_51_79_groupi_n_4235 ,csa_tree_add_51_79_groupi_n_1554 ,csa_tree_add_51_79_groupi_n_3039);
  or csa_tree_add_51_79_groupi_g42254(csa_tree_add_51_79_groupi_n_4234 ,csa_tree_add_51_79_groupi_n_1553 ,csa_tree_add_51_79_groupi_n_3045);
  or csa_tree_add_51_79_groupi_g42255(csa_tree_add_51_79_groupi_n_4233 ,csa_tree_add_51_79_groupi_n_1595 ,csa_tree_add_51_79_groupi_n_3057);
  or csa_tree_add_51_79_groupi_g42256(csa_tree_add_51_79_groupi_n_4231 ,csa_tree_add_51_79_groupi_n_1622 ,csa_tree_add_51_79_groupi_n_3110);
  or csa_tree_add_51_79_groupi_g42257(csa_tree_add_51_79_groupi_n_4230 ,csa_tree_add_51_79_groupi_n_1557 ,csa_tree_add_51_79_groupi_n_2897);
  xnor csa_tree_add_51_79_groupi_g42258(csa_tree_add_51_79_groupi_n_4229 ,csa_tree_add_51_79_groupi_n_2568 ,csa_tree_add_51_79_groupi_n_2563);
  or csa_tree_add_51_79_groupi_g42259(csa_tree_add_51_79_groupi_n_4227 ,csa_tree_add_51_79_groupi_n_1547 ,csa_tree_add_51_79_groupi_n_3693);
  and csa_tree_add_51_79_groupi_g42260(csa_tree_add_51_79_groupi_n_4226 ,csa_tree_add_51_79_groupi_n_2389 ,csa_tree_add_51_79_groupi_n_3559);
  and csa_tree_add_51_79_groupi_g42261(csa_tree_add_51_79_groupi_n_4225 ,csa_tree_add_51_79_groupi_n_2417 ,csa_tree_add_51_79_groupi_n_3704);
  not csa_tree_add_51_79_groupi_g42262(csa_tree_add_51_79_groupi_n_3871 ,csa_tree_add_51_79_groupi_n_3870);
  not csa_tree_add_51_79_groupi_g42263(csa_tree_add_51_79_groupi_n_3867 ,csa_tree_add_51_79_groupi_n_3866);
  not csa_tree_add_51_79_groupi_g42264(csa_tree_add_51_79_groupi_n_3858 ,csa_tree_add_51_79_groupi_n_3857);
  not csa_tree_add_51_79_groupi_g42265(csa_tree_add_51_79_groupi_n_3855 ,csa_tree_add_51_79_groupi_n_3854);
  not csa_tree_add_51_79_groupi_g42266(csa_tree_add_51_79_groupi_n_3850 ,csa_tree_add_51_79_groupi_n_3849);
  not csa_tree_add_51_79_groupi_g42267(csa_tree_add_51_79_groupi_n_3847 ,csa_tree_add_51_79_groupi_n_3846);
  not csa_tree_add_51_79_groupi_g42268(csa_tree_add_51_79_groupi_n_3829 ,csa_tree_add_51_79_groupi_n_3828);
  not csa_tree_add_51_79_groupi_g42269(csa_tree_add_51_79_groupi_n_3826 ,csa_tree_add_51_79_groupi_n_3827);
  not csa_tree_add_51_79_groupi_g42270(csa_tree_add_51_79_groupi_n_3824 ,csa_tree_add_51_79_groupi_n_3825);
  not csa_tree_add_51_79_groupi_g42271(csa_tree_add_51_79_groupi_n_3822 ,csa_tree_add_51_79_groupi_n_3823);
  not csa_tree_add_51_79_groupi_g42272(csa_tree_add_51_79_groupi_n_3820 ,csa_tree_add_51_79_groupi_n_3821);
  not csa_tree_add_51_79_groupi_g42273(csa_tree_add_51_79_groupi_n_3818 ,csa_tree_add_51_79_groupi_n_3819);
  not csa_tree_add_51_79_groupi_g42274(csa_tree_add_51_79_groupi_n_3816 ,csa_tree_add_51_79_groupi_n_3817);
  not csa_tree_add_51_79_groupi_g42275(csa_tree_add_51_79_groupi_n_3814 ,csa_tree_add_51_79_groupi_n_3813);
  not csa_tree_add_51_79_groupi_g42276(csa_tree_add_51_79_groupi_n_3811 ,csa_tree_add_51_79_groupi_n_3812);
  not csa_tree_add_51_79_groupi_g42277(csa_tree_add_51_79_groupi_n_3809 ,csa_tree_add_51_79_groupi_n_3810);
  not csa_tree_add_51_79_groupi_g42278(csa_tree_add_51_79_groupi_n_3807 ,csa_tree_add_51_79_groupi_n_3808);
  not csa_tree_add_51_79_groupi_g42279(csa_tree_add_51_79_groupi_n_3805 ,csa_tree_add_51_79_groupi_n_3806);
  not csa_tree_add_51_79_groupi_g42280(csa_tree_add_51_79_groupi_n_3802 ,csa_tree_add_51_79_groupi_n_3803);
  not csa_tree_add_51_79_groupi_g42281(csa_tree_add_51_79_groupi_n_3798 ,csa_tree_add_51_79_groupi_n_3799);
  not csa_tree_add_51_79_groupi_g42282(csa_tree_add_51_79_groupi_n_3793 ,csa_tree_add_51_79_groupi_n_3794);
  not csa_tree_add_51_79_groupi_g42283(csa_tree_add_51_79_groupi_n_3791 ,csa_tree_add_51_79_groupi_n_3792);
  not csa_tree_add_51_79_groupi_g42284(csa_tree_add_51_79_groupi_n_3788 ,csa_tree_add_51_79_groupi_n_3789);
  not csa_tree_add_51_79_groupi_g42285(csa_tree_add_51_79_groupi_n_3784 ,csa_tree_add_51_79_groupi_n_3785);
  not csa_tree_add_51_79_groupi_g42286(csa_tree_add_51_79_groupi_n_3782 ,csa_tree_add_51_79_groupi_n_3783);
  not csa_tree_add_51_79_groupi_g42287(csa_tree_add_51_79_groupi_n_3779 ,csa_tree_add_51_79_groupi_n_3780);
  not csa_tree_add_51_79_groupi_g42288(csa_tree_add_51_79_groupi_n_3777 ,csa_tree_add_51_79_groupi_n_3778);
  not csa_tree_add_51_79_groupi_g42289(csa_tree_add_51_79_groupi_n_3774 ,csa_tree_add_51_79_groupi_n_3775);
  not csa_tree_add_51_79_groupi_g42290(csa_tree_add_51_79_groupi_n_3772 ,csa_tree_add_51_79_groupi_n_3773);
  not csa_tree_add_51_79_groupi_g42291(csa_tree_add_51_79_groupi_n_3770 ,csa_tree_add_51_79_groupi_n_3771);
  not csa_tree_add_51_79_groupi_g42292(csa_tree_add_51_79_groupi_n_3768 ,csa_tree_add_51_79_groupi_n_3769);
  not csa_tree_add_51_79_groupi_g42293(csa_tree_add_51_79_groupi_n_3766 ,csa_tree_add_51_79_groupi_n_3767);
  not csa_tree_add_51_79_groupi_g42294(csa_tree_add_51_79_groupi_n_3764 ,csa_tree_add_51_79_groupi_n_3765);
  not csa_tree_add_51_79_groupi_g42295(csa_tree_add_51_79_groupi_n_3761 ,csa_tree_add_51_79_groupi_n_3762);
  not csa_tree_add_51_79_groupi_g42296(csa_tree_add_51_79_groupi_n_3759 ,csa_tree_add_51_79_groupi_n_3760);
  not csa_tree_add_51_79_groupi_g42297(csa_tree_add_51_79_groupi_n_3756 ,csa_tree_add_51_79_groupi_n_3757);
  not csa_tree_add_51_79_groupi_g42298(csa_tree_add_51_79_groupi_n_3754 ,csa_tree_add_51_79_groupi_n_3755);
  not csa_tree_add_51_79_groupi_g42299(csa_tree_add_51_79_groupi_n_3751 ,csa_tree_add_51_79_groupi_n_3752);
  not csa_tree_add_51_79_groupi_g42300(csa_tree_add_51_79_groupi_n_3749 ,csa_tree_add_51_79_groupi_n_3750);
  not csa_tree_add_51_79_groupi_g42301(csa_tree_add_51_79_groupi_n_3747 ,csa_tree_add_51_79_groupi_n_3748);
  not csa_tree_add_51_79_groupi_g42302(csa_tree_add_51_79_groupi_n_3745 ,csa_tree_add_51_79_groupi_n_3746);
  not csa_tree_add_51_79_groupi_g42303(csa_tree_add_51_79_groupi_n_3741 ,csa_tree_add_51_79_groupi_n_3740);
  not csa_tree_add_51_79_groupi_g42304(csa_tree_add_51_79_groupi_n_3736 ,csa_tree_add_51_79_groupi_n_3735);
  not csa_tree_add_51_79_groupi_g42305(csa_tree_add_51_79_groupi_n_3733 ,csa_tree_add_51_79_groupi_n_3734);
  or csa_tree_add_51_79_groupi_g42306(csa_tree_add_51_79_groupi_n_3704 ,csa_tree_add_51_79_groupi_n_1781 ,csa_tree_add_51_79_groupi_n_2429);
  or csa_tree_add_51_79_groupi_g42307(csa_tree_add_51_79_groupi_n_3703 ,csa_tree_add_51_79_groupi_n_601 ,csa_tree_add_51_79_groupi_n_2631);
  or csa_tree_add_51_79_groupi_g42308(csa_tree_add_51_79_groupi_n_3702 ,csa_tree_add_51_79_groupi_n_595 ,csa_tree_add_51_79_groupi_n_2083);
  or csa_tree_add_51_79_groupi_g42309(csa_tree_add_51_79_groupi_n_3701 ,csa_tree_add_51_79_groupi_n_593 ,csa_tree_add_51_79_groupi_n_2297);
  or csa_tree_add_51_79_groupi_g42310(csa_tree_add_51_79_groupi_n_3700 ,csa_tree_add_51_79_groupi_n_531 ,csa_tree_add_51_79_groupi_n_2095);
  or csa_tree_add_51_79_groupi_g42311(csa_tree_add_51_79_groupi_n_3699 ,csa_tree_add_51_79_groupi_n_557 ,csa_tree_add_51_79_groupi_n_2656);
  or csa_tree_add_51_79_groupi_g42312(csa_tree_add_51_79_groupi_n_3698 ,csa_tree_add_51_79_groupi_n_588 ,csa_tree_add_51_79_groupi_n_2676);
  or csa_tree_add_51_79_groupi_g42313(csa_tree_add_51_79_groupi_n_3697 ,csa_tree_add_51_79_groupi_n_590 ,csa_tree_add_51_79_groupi_n_2298);
  or csa_tree_add_51_79_groupi_g42314(csa_tree_add_51_79_groupi_n_3696 ,csa_tree_add_51_79_groupi_n_552 ,csa_tree_add_51_79_groupi_n_2810);
  or csa_tree_add_51_79_groupi_g42315(csa_tree_add_51_79_groupi_n_3695 ,csa_tree_add_51_79_groupi_n_544 ,csa_tree_add_51_79_groupi_n_2841);
  or csa_tree_add_51_79_groupi_g42316(csa_tree_add_51_79_groupi_n_3694 ,csa_tree_add_51_79_groupi_n_526 ,csa_tree_add_51_79_groupi_n_2830);
  nor csa_tree_add_51_79_groupi_g42317(csa_tree_add_51_79_groupi_n_3693 ,csa_tree_add_51_79_groupi_n_1704 ,csa_tree_add_51_79_groupi_n_2421);
  or csa_tree_add_51_79_groupi_g42318(csa_tree_add_51_79_groupi_n_3692 ,csa_tree_add_51_79_groupi_n_536 ,csa_tree_add_51_79_groupi_n_2098);
  or csa_tree_add_51_79_groupi_g42319(csa_tree_add_51_79_groupi_n_3691 ,csa_tree_add_51_79_groupi_n_533 ,csa_tree_add_51_79_groupi_n_2285);
  or csa_tree_add_51_79_groupi_g42320(csa_tree_add_51_79_groupi_n_3690 ,csa_tree_add_51_79_groupi_n_554 ,csa_tree_add_51_79_groupi_n_2578);
  or csa_tree_add_51_79_groupi_g42321(csa_tree_add_51_79_groupi_n_3689 ,csa_tree_add_51_79_groupi_n_881 ,csa_tree_add_51_79_groupi_n_2870);
  nor csa_tree_add_51_79_groupi_g42322(csa_tree_add_51_79_groupi_n_3688 ,csa_tree_add_51_79_groupi_n_1680 ,csa_tree_add_51_79_groupi_n_2430);
  or csa_tree_add_51_79_groupi_g42323(csa_tree_add_51_79_groupi_n_3687 ,csa_tree_add_51_79_groupi_n_546 ,csa_tree_add_51_79_groupi_n_2293);
  or csa_tree_add_51_79_groupi_g42324(csa_tree_add_51_79_groupi_n_3686 ,csa_tree_add_51_79_groupi_n_598 ,csa_tree_add_51_79_groupi_n_2314);
  or csa_tree_add_51_79_groupi_g42325(csa_tree_add_51_79_groupi_n_3685 ,csa_tree_add_51_79_groupi_n_538 ,csa_tree_add_51_79_groupi_n_2818);
  or csa_tree_add_51_79_groupi_g42326(csa_tree_add_51_79_groupi_n_3684 ,csa_tree_add_51_79_groupi_n_528 ,csa_tree_add_51_79_groupi_n_2883);
  or csa_tree_add_51_79_groupi_g42327(csa_tree_add_51_79_groupi_n_3683 ,csa_tree_add_51_79_groupi_n_603 ,csa_tree_add_51_79_groupi_n_2099);
  or csa_tree_add_51_79_groupi_g42328(csa_tree_add_51_79_groupi_n_3682 ,csa_tree_add_51_79_groupi_n_605 ,csa_tree_add_51_79_groupi_n_2685);
  or csa_tree_add_51_79_groupi_g42329(csa_tree_add_51_79_groupi_n_3681 ,csa_tree_add_51_79_groupi_n_886 ,csa_tree_add_51_79_groupi_n_2300);
  or csa_tree_add_51_79_groupi_g42330(csa_tree_add_51_79_groupi_n_3680 ,csa_tree_add_51_79_groupi_n_523 ,csa_tree_add_51_79_groupi_n_2037);
  or csa_tree_add_51_79_groupi_g42331(csa_tree_add_51_79_groupi_n_3679 ,csa_tree_add_51_79_groupi_n_821 ,csa_tree_add_51_79_groupi_n_2584);
  or csa_tree_add_51_79_groupi_g42332(csa_tree_add_51_79_groupi_n_3678 ,csa_tree_add_51_79_groupi_n_541 ,csa_tree_add_51_79_groupi_n_2315);
  or csa_tree_add_51_79_groupi_g42333(csa_tree_add_51_79_groupi_n_3677 ,csa_tree_add_51_79_groupi_n_888 ,csa_tree_add_51_79_groupi_n_2651);
  or csa_tree_add_51_79_groupi_g42334(csa_tree_add_51_79_groupi_n_3676 ,csa_tree_add_51_79_groupi_n_549 ,csa_tree_add_51_79_groupi_n_2308);
  or csa_tree_add_51_79_groupi_g42335(csa_tree_add_51_79_groupi_n_3675 ,csa_tree_add_51_79_groupi_n_862 ,csa_tree_add_51_79_groupi_n_2309);
  or csa_tree_add_51_79_groupi_g42336(csa_tree_add_51_79_groupi_n_3674 ,csa_tree_add_51_79_groupi_n_559 ,csa_tree_add_51_79_groupi_n_2667);
  or csa_tree_add_51_79_groupi_g42337(csa_tree_add_51_79_groupi_n_3673 ,csa_tree_add_51_79_groupi_n_876 ,csa_tree_add_51_79_groupi_n_2877);
  or csa_tree_add_51_79_groupi_g42338(csa_tree_add_51_79_groupi_n_3672 ,csa_tree_add_51_79_groupi_n_862 ,csa_tree_add_51_79_groupi_n_2824);
  or csa_tree_add_51_79_groupi_g42339(csa_tree_add_51_79_groupi_n_3671 ,csa_tree_add_51_79_groupi_n_864 ,csa_tree_add_51_79_groupi_n_2038);
  or csa_tree_add_51_79_groupi_g42340(csa_tree_add_51_79_groupi_n_3670 ,csa_tree_add_51_79_groupi_n_886 ,csa_tree_add_51_79_groupi_n_2283);
  or csa_tree_add_51_79_groupi_g42341(csa_tree_add_51_79_groupi_n_3669 ,csa_tree_add_51_79_groupi_n_857 ,csa_tree_add_51_79_groupi_n_2022);
  or csa_tree_add_51_79_groupi_g42342(csa_tree_add_51_79_groupi_n_3668 ,csa_tree_add_51_79_groupi_n_857 ,csa_tree_add_51_79_groupi_n_2035);
  or csa_tree_add_51_79_groupi_g42343(csa_tree_add_51_79_groupi_n_3667 ,csa_tree_add_51_79_groupi_n_823 ,csa_tree_add_51_79_groupi_n_2614);
  or csa_tree_add_51_79_groupi_g42344(csa_tree_add_51_79_groupi_n_3666 ,csa_tree_add_51_79_groupi_n_871 ,csa_tree_add_51_79_groupi_n_2016);
  or csa_tree_add_51_79_groupi_g42345(csa_tree_add_51_79_groupi_n_3665 ,csa_tree_add_51_79_groupi_n_528 ,csa_tree_add_51_79_groupi_n_2574);
  or csa_tree_add_51_79_groupi_g42346(csa_tree_add_51_79_groupi_n_3664 ,csa_tree_add_51_79_groupi_n_526 ,csa_tree_add_51_79_groupi_n_2625);
  or csa_tree_add_51_79_groupi_g42347(csa_tree_add_51_79_groupi_n_3663 ,csa_tree_add_51_79_groupi_n_821 ,csa_tree_add_51_79_groupi_n_2803);
  or csa_tree_add_51_79_groupi_g42348(csa_tree_add_51_79_groupi_n_3662 ,csa_tree_add_51_79_groupi_n_888 ,csa_tree_add_51_79_groupi_n_2316);
  or csa_tree_add_51_79_groupi_g42349(csa_tree_add_51_79_groupi_n_3661 ,csa_tree_add_51_79_groupi_n_871 ,csa_tree_add_51_79_groupi_n_2799);
  or csa_tree_add_51_79_groupi_g42350(csa_tree_add_51_79_groupi_n_3660 ,csa_tree_add_51_79_groupi_n_603 ,csa_tree_add_51_79_groupi_n_2688);
  or csa_tree_add_51_79_groupi_g42351(csa_tree_add_51_79_groupi_n_3659 ,csa_tree_add_51_79_groupi_n_2169 ,csa_tree_add_51_79_groupi_n_1369);
  or csa_tree_add_51_79_groupi_g42352(csa_tree_add_51_79_groupi_n_3658 ,csa_tree_add_51_79_groupi_n_886 ,csa_tree_add_51_79_groupi_n_2170);
  or csa_tree_add_51_79_groupi_g42353(csa_tree_add_51_79_groupi_n_3657 ,csa_tree_add_51_79_groupi_n_2679 ,csa_tree_add_51_79_groupi_n_1384);
  or csa_tree_add_51_79_groupi_g42354(csa_tree_add_51_79_groupi_n_3656 ,csa_tree_add_51_79_groupi_n_881 ,csa_tree_add_51_79_groupi_n_2627);
  or csa_tree_add_51_79_groupi_g42355(csa_tree_add_51_79_groupi_n_3655 ,csa_tree_add_51_79_groupi_n_607 ,csa_tree_add_51_79_groupi_n_2767);
  or csa_tree_add_51_79_groupi_g42356(csa_tree_add_51_79_groupi_n_3654 ,csa_tree_add_51_79_groupi_n_2139 ,csa_tree_add_51_79_groupi_n_706);
  or csa_tree_add_51_79_groupi_g42357(csa_tree_add_51_79_groupi_n_3653 ,csa_tree_add_51_79_groupi_n_828 ,csa_tree_add_51_79_groupi_n_2619);
  or csa_tree_add_51_79_groupi_g42358(csa_tree_add_51_79_groupi_n_3652 ,csa_tree_add_51_79_groupi_n_523 ,csa_tree_add_51_79_groupi_n_2108);
  or csa_tree_add_51_79_groupi_g42359(csa_tree_add_51_79_groupi_n_3651 ,csa_tree_add_51_79_groupi_n_864 ,csa_tree_add_51_79_groupi_n_2735);
  or csa_tree_add_51_79_groupi_g42360(csa_tree_add_51_79_groupi_n_3650 ,csa_tree_add_51_79_groupi_n_823 ,csa_tree_add_51_79_groupi_n_2615);
  or csa_tree_add_51_79_groupi_g42361(csa_tree_add_51_79_groupi_n_3649 ,csa_tree_add_51_79_groupi_n_2876 ,csa_tree_add_51_79_groupi_n_1336);
  or csa_tree_add_51_79_groupi_g42362(csa_tree_add_51_79_groupi_n_3648 ,csa_tree_add_51_79_groupi_n_828 ,csa_tree_add_51_79_groupi_n_2047);
  or csa_tree_add_51_79_groupi_g42363(csa_tree_add_51_79_groupi_n_3647 ,csa_tree_add_51_79_groupi_n_2195 ,csa_tree_add_51_79_groupi_n_1417);
  or csa_tree_add_51_79_groupi_g42364(csa_tree_add_51_79_groupi_n_3646 ,csa_tree_add_51_79_groupi_n_607 ,csa_tree_add_51_79_groupi_n_2812);
  or csa_tree_add_51_79_groupi_g42365(csa_tree_add_51_79_groupi_n_3645 ,csa_tree_add_51_79_groupi_n_605 ,csa_tree_add_51_79_groupi_n_2588);
  or csa_tree_add_51_79_groupi_g42366(csa_tree_add_51_79_groupi_n_3644 ,csa_tree_add_51_79_groupi_n_2729 ,csa_tree_add_51_79_groupi_n_682);
  or csa_tree_add_51_79_groupi_g42367(csa_tree_add_51_79_groupi_n_3643 ,csa_tree_add_51_79_groupi_n_598 ,csa_tree_add_51_79_groupi_n_2312);
  or csa_tree_add_51_79_groupi_g42368(csa_tree_add_51_79_groupi_n_3642 ,csa_tree_add_51_79_groupi_n_2305 ,csa_tree_add_51_79_groupi_n_736);
  or csa_tree_add_51_79_groupi_g42369(csa_tree_add_51_79_groupi_n_3641 ,csa_tree_add_51_79_groupi_n_869 ,csa_tree_add_51_79_groupi_n_2126);
  or csa_tree_add_51_79_groupi_g42370(csa_tree_add_51_79_groupi_n_3640 ,csa_tree_add_51_79_groupi_n_869 ,csa_tree_add_51_79_groupi_n_2848);
  or csa_tree_add_51_79_groupi_g42371(csa_tree_add_51_79_groupi_n_3639 ,csa_tree_add_51_79_groupi_n_554 ,csa_tree_add_51_79_groupi_n_2807);
  or csa_tree_add_51_79_groupi_g42372(csa_tree_add_51_79_groupi_n_3638 ,csa_tree_add_51_79_groupi_n_541 ,csa_tree_add_51_79_groupi_n_2745);
  or csa_tree_add_51_79_groupi_g42373(csa_tree_add_51_79_groupi_n_3637 ,csa_tree_add_51_79_groupi_n_590 ,csa_tree_add_51_79_groupi_n_2695);
  or csa_tree_add_51_79_groupi_g42374(csa_tree_add_51_79_groupi_n_3636 ,csa_tree_add_51_79_groupi_n_886 ,csa_tree_add_51_79_groupi_n_2683);
  or csa_tree_add_51_79_groupi_g42375(csa_tree_add_51_79_groupi_n_3635 ,csa_tree_add_51_79_groupi_n_601 ,csa_tree_add_51_79_groupi_n_2073);
  or csa_tree_add_51_79_groupi_g42376(csa_tree_add_51_79_groupi_n_3634 ,csa_tree_add_51_79_groupi_n_533 ,csa_tree_add_51_79_groupi_n_2580);
  or csa_tree_add_51_79_groupi_g42377(csa_tree_add_51_79_groupi_n_3633 ,csa_tree_add_51_79_groupi_n_552 ,csa_tree_add_51_79_groupi_n_2110);
  or csa_tree_add_51_79_groupi_g42378(csa_tree_add_51_79_groupi_n_3632 ,csa_tree_add_51_79_groupi_n_531 ,csa_tree_add_51_79_groupi_n_2636);
  or csa_tree_add_51_79_groupi_g42379(csa_tree_add_51_79_groupi_n_3631 ,csa_tree_add_51_79_groupi_n_546 ,csa_tree_add_51_79_groupi_n_2785);
  or csa_tree_add_51_79_groupi_g42380(csa_tree_add_51_79_groupi_n_3630 ,csa_tree_add_51_79_groupi_n_823 ,csa_tree_add_51_79_groupi_n_2776);
  or csa_tree_add_51_79_groupi_g42381(csa_tree_add_51_79_groupi_n_3629 ,csa_tree_add_51_79_groupi_n_876 ,csa_tree_add_51_79_groupi_n_2748);
  or csa_tree_add_51_79_groupi_g42382(csa_tree_add_51_79_groupi_n_3628 ,csa_tree_add_51_79_groupi_n_2253 ,csa_tree_add_51_79_groupi_n_697);
  or csa_tree_add_51_79_groupi_g42383(csa_tree_add_51_79_groupi_n_3627 ,csa_tree_add_51_79_groupi_n_549 ,csa_tree_add_51_79_groupi_n_2825);
  or csa_tree_add_51_79_groupi_g42384(csa_tree_add_51_79_groupi_n_3626 ,csa_tree_add_51_79_groupi_n_595 ,csa_tree_add_51_79_groupi_n_2677);
  or csa_tree_add_51_79_groupi_g42385(csa_tree_add_51_79_groupi_n_3625 ,csa_tree_add_51_79_groupi_n_588 ,csa_tree_add_51_79_groupi_n_2104);
  or csa_tree_add_51_79_groupi_g42386(csa_tree_add_51_79_groupi_n_3624 ,csa_tree_add_51_79_groupi_n_544 ,csa_tree_add_51_79_groupi_n_2072);
  or csa_tree_add_51_79_groupi_g42387(csa_tree_add_51_79_groupi_n_3623 ,csa_tree_add_51_79_groupi_n_871 ,csa_tree_add_51_79_groupi_n_2632);
  or csa_tree_add_51_79_groupi_g42388(csa_tree_add_51_79_groupi_n_3622 ,csa_tree_add_51_79_groupi_n_871 ,csa_tree_add_51_79_groupi_n_2657);
  or csa_tree_add_51_79_groupi_g42389(csa_tree_add_51_79_groupi_n_3621 ,csa_tree_add_51_79_groupi_n_559 ,csa_tree_add_51_79_groupi_n_2062);
  or csa_tree_add_51_79_groupi_g42390(csa_tree_add_51_79_groupi_n_3620 ,csa_tree_add_51_79_groupi_n_823 ,csa_tree_add_51_79_groupi_n_2630);
  or csa_tree_add_51_79_groupi_g42391(csa_tree_add_51_79_groupi_n_3619 ,csa_tree_add_51_79_groupi_n_538 ,csa_tree_add_51_79_groupi_n_2727);
  or csa_tree_add_51_79_groupi_g42392(csa_tree_add_51_79_groupi_n_3618 ,csa_tree_add_51_79_groupi_n_821 ,csa_tree_add_51_79_groupi_n_2048);
  or csa_tree_add_51_79_groupi_g42393(csa_tree_add_51_79_groupi_n_3617 ,csa_tree_add_51_79_groupi_n_862 ,csa_tree_add_51_79_groupi_n_2734);
  or csa_tree_add_51_79_groupi_g42394(csa_tree_add_51_79_groupi_n_3616 ,csa_tree_add_51_79_groupi_n_593 ,csa_tree_add_51_79_groupi_n_2610);
  or csa_tree_add_51_79_groupi_g42395(csa_tree_add_51_79_groupi_n_3615 ,csa_tree_add_51_79_groupi_n_869 ,csa_tree_add_51_79_groupi_n_2689);
  or csa_tree_add_51_79_groupi_g42396(csa_tree_add_51_79_groupi_n_3614 ,csa_tree_add_51_79_groupi_n_869 ,csa_tree_add_51_79_groupi_n_2700);
  or csa_tree_add_51_79_groupi_g42397(csa_tree_add_51_79_groupi_n_3613 ,csa_tree_add_51_79_groupi_n_862 ,csa_tree_add_51_79_groupi_n_2214);
  or csa_tree_add_51_79_groupi_g42398(csa_tree_add_51_79_groupi_n_3612 ,csa_tree_add_51_79_groupi_n_536 ,csa_tree_add_51_79_groupi_n_2076);
  or csa_tree_add_51_79_groupi_g42399(csa_tree_add_51_79_groupi_n_3611 ,csa_tree_add_51_79_groupi_n_821 ,csa_tree_add_51_79_groupi_n_2758);
  or csa_tree_add_51_79_groupi_g42400(csa_tree_add_51_79_groupi_n_3610 ,csa_tree_add_51_79_groupi_n_2211 ,csa_tree_add_51_79_groupi_n_1258);
  or csa_tree_add_51_79_groupi_g42401(csa_tree_add_51_79_groupi_n_3609 ,csa_tree_add_51_79_groupi_n_881 ,csa_tree_add_51_79_groupi_n_2696);
  or csa_tree_add_51_79_groupi_g42402(csa_tree_add_51_79_groupi_n_3608 ,csa_tree_add_51_79_groupi_n_888 ,csa_tree_add_51_79_groupi_n_2018);
  or csa_tree_add_51_79_groupi_g42403(csa_tree_add_51_79_groupi_n_3607 ,csa_tree_add_51_79_groupi_n_864 ,csa_tree_add_51_79_groupi_n_2851);
  or csa_tree_add_51_79_groupi_g42404(csa_tree_add_51_79_groupi_n_3606 ,csa_tree_add_51_79_groupi_n_557 ,csa_tree_add_51_79_groupi_n_2784);
  or csa_tree_add_51_79_groupi_g42405(csa_tree_add_51_79_groupi_n_3605 ,csa_tree_add_51_79_groupi_n_857 ,csa_tree_add_51_79_groupi_n_2875);
  or csa_tree_add_51_79_groupi_g42406(csa_tree_add_51_79_groupi_n_3604 ,csa_tree_add_51_79_groupi_n_864 ,csa_tree_add_51_79_groupi_n_2576);
  or csa_tree_add_51_79_groupi_g42407(csa_tree_add_51_79_groupi_n_3603 ,csa_tree_add_51_79_groupi_n_876 ,csa_tree_add_51_79_groupi_n_2644);
  or csa_tree_add_51_79_groupi_g42408(csa_tree_add_51_79_groupi_n_3602 ,csa_tree_add_51_79_groupi_n_876 ,csa_tree_add_51_79_groupi_n_2025);
  or csa_tree_add_51_79_groupi_g42409(csa_tree_add_51_79_groupi_n_3601 ,csa_tree_add_51_79_groupi_n_828 ,csa_tree_add_51_79_groupi_n_2831);
  or csa_tree_add_51_79_groupi_g42410(csa_tree_add_51_79_groupi_n_3600 ,csa_tree_add_51_79_groupi_n_828 ,csa_tree_add_51_79_groupi_n_2686);
  or csa_tree_add_51_79_groupi_g42411(csa_tree_add_51_79_groupi_n_3599 ,csa_tree_add_51_79_groupi_n_821 ,csa_tree_add_51_79_groupi_n_2866);
  or csa_tree_add_51_79_groupi_g42412(csa_tree_add_51_79_groupi_n_3598 ,csa_tree_add_51_79_groupi_n_823 ,csa_tree_add_51_79_groupi_n_2077);
  or csa_tree_add_51_79_groupi_g42413(csa_tree_add_51_79_groupi_n_3597 ,csa_tree_add_51_79_groupi_n_862 ,csa_tree_add_51_79_groupi_n_2113);
  or csa_tree_add_51_79_groupi_g42414(csa_tree_add_51_79_groupi_n_3596 ,csa_tree_add_51_79_groupi_n_828 ,csa_tree_add_51_79_groupi_n_2029);
  or csa_tree_add_51_79_groupi_g42415(csa_tree_add_51_79_groupi_n_3595 ,csa_tree_add_51_79_groupi_n_886 ,csa_tree_add_51_79_groupi_n_2061);
  or csa_tree_add_51_79_groupi_g42416(csa_tree_add_51_79_groupi_n_3594 ,csa_tree_add_51_79_groupi_n_876 ,csa_tree_add_51_79_groupi_n_2053);
  or csa_tree_add_51_79_groupi_g42417(csa_tree_add_51_79_groupi_n_3593 ,csa_tree_add_51_79_groupi_n_869 ,csa_tree_add_51_79_groupi_n_2058);
  or csa_tree_add_51_79_groupi_g42418(csa_tree_add_51_79_groupi_n_3592 ,csa_tree_add_51_79_groupi_n_540 ,csa_tree_add_51_79_groupi_n_2713);
  or csa_tree_add_51_79_groupi_g42419(csa_tree_add_51_79_groupi_n_3591 ,csa_tree_add_51_79_groupi_n_548 ,csa_tree_add_51_79_groupi_n_2814);
  or csa_tree_add_51_79_groupi_g42420(csa_tree_add_51_79_groupi_n_3590 ,csa_tree_add_51_79_groupi_n_888 ,csa_tree_add_51_79_groupi_n_2119);
  or csa_tree_add_51_79_groupi_g42421(csa_tree_add_51_79_groupi_n_3589 ,csa_tree_add_51_79_groupi_n_857 ,csa_tree_add_51_79_groupi_n_2028);
  or csa_tree_add_51_79_groupi_g42422(csa_tree_add_51_79_groupi_n_3588 ,csa_tree_add_51_79_groupi_n_857 ,csa_tree_add_51_79_groupi_n_2852);
  or csa_tree_add_51_79_groupi_g42423(csa_tree_add_51_79_groupi_n_3587 ,csa_tree_add_51_79_groupi_n_881 ,csa_tree_add_51_79_groupi_n_2880);
  or csa_tree_add_51_79_groupi_g42424(csa_tree_add_51_79_groupi_n_3586 ,csa_tree_add_51_79_groupi_n_522 ,csa_tree_add_51_79_groupi_n_2594);
  or csa_tree_add_51_79_groupi_g42425(csa_tree_add_51_79_groupi_n_3585 ,csa_tree_add_51_79_groupi_n_881 ,csa_tree_add_51_79_groupi_n_2771);
  or csa_tree_add_51_79_groupi_g42426(csa_tree_add_51_79_groupi_n_3584 ,csa_tree_add_51_79_groupi_n_2820 ,csa_tree_add_51_79_groupi_n_1339);
  or csa_tree_add_51_79_groupi_g42427(csa_tree_add_51_79_groupi_n_3583 ,csa_tree_add_51_79_groupi_n_2661 ,csa_tree_add_51_79_groupi_n_1402);
  or csa_tree_add_51_79_groupi_g42428(csa_tree_add_51_79_groupi_n_3582 ,csa_tree_add_51_79_groupi_n_2879 ,csa_tree_add_51_79_groupi_n_748);
  or csa_tree_add_51_79_groupi_g42429(csa_tree_add_51_79_groupi_n_3581 ,csa_tree_add_51_79_groupi_n_2774 ,csa_tree_add_51_79_groupi_n_1354);
  or csa_tree_add_51_79_groupi_g42430(csa_tree_add_51_79_groupi_n_3580 ,csa_tree_add_51_79_groupi_n_2248 ,csa_tree_add_51_79_groupi_n_673);
  or csa_tree_add_51_79_groupi_g42431(csa_tree_add_51_79_groupi_n_3579 ,csa_tree_add_51_79_groupi_n_2857 ,csa_tree_add_51_79_groupi_n_1264);
  or csa_tree_add_51_79_groupi_g42432(csa_tree_add_51_79_groupi_n_3578 ,csa_tree_add_51_79_groupi_n_2218 ,csa_tree_add_51_79_groupi_n_709);
  or csa_tree_add_51_79_groupi_g42433(csa_tree_add_51_79_groupi_n_3577 ,csa_tree_add_51_79_groupi_n_2760 ,csa_tree_add_51_79_groupi_n_712);
  or csa_tree_add_51_79_groupi_g42434(csa_tree_add_51_79_groupi_n_3576 ,csa_tree_add_51_79_groupi_n_2741 ,csa_tree_add_51_79_groupi_n_751);
  nor csa_tree_add_51_79_groupi_g42435(csa_tree_add_51_79_groupi_n_3575 ,csa_tree_add_51_79_groupi_n_1766 ,csa_tree_add_51_79_groupi_n_2401);
  or csa_tree_add_51_79_groupi_g42436(csa_tree_add_51_79_groupi_n_3574 ,csa_tree_add_51_79_groupi_n_2873 ,csa_tree_add_51_79_groupi_n_1294);
  or csa_tree_add_51_79_groupi_g42437(csa_tree_add_51_79_groupi_n_3573 ,csa_tree_add_51_79_groupi_n_2220 ,csa_tree_add_51_79_groupi_n_1318);
  nor csa_tree_add_51_79_groupi_g42438(csa_tree_add_51_79_groupi_n_3572 ,csa_tree_add_51_79_groupi_n_1714 ,csa_tree_add_51_79_groupi_n_2384);
  nor csa_tree_add_51_79_groupi_g42439(csa_tree_add_51_79_groupi_n_3571 ,csa_tree_add_51_79_groupi_n_1677 ,csa_tree_add_51_79_groupi_n_2431);
  or csa_tree_add_51_79_groupi_g42440(csa_tree_add_51_79_groupi_n_3570 ,csa_tree_add_51_79_groupi_n_2209 ,csa_tree_add_51_79_groupi_n_1426);
  or csa_tree_add_51_79_groupi_g42441(csa_tree_add_51_79_groupi_n_3569 ,csa_tree_add_51_79_groupi_n_2051 ,csa_tree_add_51_79_groupi_n_730);
  or csa_tree_add_51_79_groupi_g42442(csa_tree_add_51_79_groupi_n_3568 ,csa_tree_add_51_79_groupi_n_2177 ,csa_tree_add_51_79_groupi_n_1372);
  or csa_tree_add_51_79_groupi_g42443(csa_tree_add_51_79_groupi_n_3567 ,csa_tree_add_51_79_groupi_n_2609 ,csa_tree_add_51_79_groupi_n_1357);
  nor csa_tree_add_51_79_groupi_g42444(csa_tree_add_51_79_groupi_n_3566 ,csa_tree_add_51_79_groupi_n_1768 ,csa_tree_add_51_79_groupi_n_2392);
  or csa_tree_add_51_79_groupi_g42445(csa_tree_add_51_79_groupi_n_3565 ,csa_tree_add_51_79_groupi_n_2716 ,csa_tree_add_51_79_groupi_n_1336);
  and csa_tree_add_51_79_groupi_g42446(csa_tree_add_51_79_groupi_n_3564 ,csa_tree_add_51_79_groupi_n_2550 ,csa_tree_add_51_79_groupi_n_2541);
  or csa_tree_add_51_79_groupi_g42447(csa_tree_add_51_79_groupi_n_3563 ,csa_tree_add_51_79_groupi_n_2821 ,csa_tree_add_51_79_groupi_n_1420);
  or csa_tree_add_51_79_groupi_g42448(csa_tree_add_51_79_groupi_n_3562 ,csa_tree_add_51_79_groupi_n_2164 ,csa_tree_add_51_79_groupi_n_700);
  or csa_tree_add_51_79_groupi_g42449(csa_tree_add_51_79_groupi_n_3561 ,csa_tree_add_51_79_groupi_n_2744 ,csa_tree_add_51_79_groupi_n_1297);
  or csa_tree_add_51_79_groupi_g42450(csa_tree_add_51_79_groupi_n_3560 ,csa_tree_add_51_79_groupi_n_2681 ,csa_tree_add_51_79_groupi_n_1390);
  or csa_tree_add_51_79_groupi_g42451(csa_tree_add_51_79_groupi_n_3559 ,csa_tree_add_51_79_groupi_n_1787 ,csa_tree_add_51_79_groupi_n_2394);
  or csa_tree_add_51_79_groupi_g42452(csa_tree_add_51_79_groupi_n_3558 ,csa_tree_add_51_79_groupi_n_2755 ,csa_tree_add_51_79_groupi_n_1252);
  or csa_tree_add_51_79_groupi_g42453(csa_tree_add_51_79_groupi_n_3557 ,csa_tree_add_51_79_groupi_n_2751 ,csa_tree_add_51_79_groupi_n_1444);
  or csa_tree_add_51_79_groupi_g42454(csa_tree_add_51_79_groupi_n_3556 ,csa_tree_add_51_79_groupi_n_2813 ,csa_tree_add_51_79_groupi_n_1339);
  or csa_tree_add_51_79_groupi_g42455(csa_tree_add_51_79_groupi_n_3555 ,csa_tree_add_51_79_groupi_n_2290 ,csa_tree_add_51_79_groupi_n_1411);
  or csa_tree_add_51_79_groupi_g42456(csa_tree_add_51_79_groupi_n_3554 ,csa_tree_add_51_79_groupi_n_2266 ,csa_tree_add_51_79_groupi_n_1219);
  or csa_tree_add_51_79_groupi_g42457(csa_tree_add_51_79_groupi_n_3553 ,csa_tree_add_51_79_groupi_n_2237 ,csa_tree_add_51_79_groupi_n_694);
  or csa_tree_add_51_79_groupi_g42458(csa_tree_add_51_79_groupi_n_3552 ,csa_tree_add_51_79_groupi_n_2711 ,csa_tree_add_51_79_groupi_n_1324);
  or csa_tree_add_51_79_groupi_g42459(csa_tree_add_51_79_groupi_n_3551 ,csa_tree_add_51_79_groupi_n_2138 ,csa_tree_add_51_79_groupi_n_1417);
  or csa_tree_add_51_79_groupi_g42460(csa_tree_add_51_79_groupi_n_3550 ,csa_tree_add_51_79_groupi_n_2815 ,csa_tree_add_51_79_groupi_n_1342);
  or csa_tree_add_51_79_groupi_g42461(csa_tree_add_51_79_groupi_n_3549 ,csa_tree_add_51_79_groupi_n_2213 ,csa_tree_add_51_79_groupi_n_676);
  nor csa_tree_add_51_79_groupi_g42462(csa_tree_add_51_79_groupi_n_3548 ,csa_tree_add_51_79_groupi_n_1692 ,csa_tree_add_51_79_groupi_n_2413);
  or csa_tree_add_51_79_groupi_g42463(csa_tree_add_51_79_groupi_n_3547 ,csa_tree_add_51_79_groupi_n_2227 ,csa_tree_add_51_79_groupi_n_697);
  or csa_tree_add_51_79_groupi_g42464(csa_tree_add_51_79_groupi_n_3546 ,csa_tree_add_51_79_groupi_n_2224 ,csa_tree_add_51_79_groupi_n_673);
  or csa_tree_add_51_79_groupi_g42465(csa_tree_add_51_79_groupi_n_3545 ,csa_tree_add_51_79_groupi_n_2558 ,csa_tree_add_51_79_groupi_n_2552);
  or csa_tree_add_51_79_groupi_g42466(csa_tree_add_51_79_groupi_n_3544 ,csa_tree_add_51_79_groupi_n_2753 ,csa_tree_add_51_79_groupi_n_748);
  or csa_tree_add_51_79_groupi_g42467(csa_tree_add_51_79_groupi_n_3543 ,csa_tree_add_51_79_groupi_n_2737 ,csa_tree_add_51_79_groupi_n_1348);
  or csa_tree_add_51_79_groupi_g42468(csa_tree_add_51_79_groupi_n_3542 ,csa_tree_add_51_79_groupi_n_2137 ,csa_tree_add_51_79_groupi_n_673);
  or csa_tree_add_51_79_groupi_g42469(csa_tree_add_51_79_groupi_n_3541 ,csa_tree_add_51_79_groupi_n_2231 ,csa_tree_add_51_79_groupi_n_1261);
  or csa_tree_add_51_79_groupi_g42470(csa_tree_add_51_79_groupi_n_3540 ,csa_tree_add_51_79_groupi_n_2071 ,csa_tree_add_51_79_groupi_n_1270);
  or csa_tree_add_51_79_groupi_g42471(csa_tree_add_51_79_groupi_n_3539 ,csa_tree_add_51_79_groupi_n_2629 ,csa_tree_add_51_79_groupi_n_1393);
  or csa_tree_add_51_79_groupi_g42472(csa_tree_add_51_79_groupi_n_3538 ,csa_tree_add_51_79_groupi_n_2032 ,csa_tree_add_51_79_groupi_n_1312);
  or csa_tree_add_51_79_groupi_g42473(csa_tree_add_51_79_groupi_n_3537 ,csa_tree_add_51_79_groupi_n_2721 ,csa_tree_add_51_79_groupi_n_1237);
  or csa_tree_add_51_79_groupi_g42474(csa_tree_add_51_79_groupi_n_3536 ,csa_tree_add_51_79_groupi_n_2550 ,csa_tree_add_51_79_groupi_n_2541);
  or csa_tree_add_51_79_groupi_g42475(csa_tree_add_51_79_groupi_n_3535 ,csa_tree_add_51_79_groupi_n_2691 ,csa_tree_add_51_79_groupi_n_1330);
  or csa_tree_add_51_79_groupi_g42476(csa_tree_add_51_79_groupi_n_3534 ,csa_tree_add_51_79_groupi_n_2641 ,csa_tree_add_51_79_groupi_n_1351);
  or csa_tree_add_51_79_groupi_g42477(csa_tree_add_51_79_groupi_n_3533 ,csa_tree_add_51_79_groupi_n_2181 ,csa_tree_add_51_79_groupi_n_1243);
  or csa_tree_add_51_79_groupi_g42478(csa_tree_add_51_79_groupi_n_3532 ,csa_tree_add_51_79_groupi_n_2319 ,csa_tree_add_51_79_groupi_n_1276);
  or csa_tree_add_51_79_groupi_g42479(csa_tree_add_51_79_groupi_n_3531 ,csa_tree_add_51_79_groupi_n_2604 ,csa_tree_add_51_79_groupi_n_1360);
  or csa_tree_add_51_79_groupi_g42480(csa_tree_add_51_79_groupi_n_3530 ,csa_tree_add_51_79_groupi_n_2140 ,csa_tree_add_51_79_groupi_n_1441);
  or csa_tree_add_51_79_groupi_g42481(csa_tree_add_51_79_groupi_n_3529 ,csa_tree_add_51_79_groupi_n_2781 ,csa_tree_add_51_79_groupi_n_1225);
  or csa_tree_add_51_79_groupi_g42482(csa_tree_add_51_79_groupi_n_3528 ,csa_tree_add_51_79_groupi_n_2823 ,csa_tree_add_51_79_groupi_n_1327);
  or csa_tree_add_51_79_groupi_g42483(csa_tree_add_51_79_groupi_n_3527 ,csa_tree_add_51_79_groupi_n_2640 ,csa_tree_add_51_79_groupi_n_1387);
  or csa_tree_add_51_79_groupi_g42484(csa_tree_add_51_79_groupi_n_3526 ,csa_tree_add_51_79_groupi_n_2608 ,csa_tree_add_51_79_groupi_n_1384);
  or csa_tree_add_51_79_groupi_g42485(csa_tree_add_51_79_groupi_n_3525 ,csa_tree_add_51_79_groupi_n_2026 ,csa_tree_add_51_79_groupi_n_1429);
  or csa_tree_add_51_79_groupi_g42486(csa_tree_add_51_79_groupi_n_3524 ,csa_tree_add_51_79_groupi_n_2212 ,csa_tree_add_51_79_groupi_n_676);
  or csa_tree_add_51_79_groupi_g42487(csa_tree_add_51_79_groupi_n_3523 ,csa_tree_add_51_79_groupi_n_2114 ,csa_tree_add_51_79_groupi_n_739);
  or csa_tree_add_51_79_groupi_g42488(csa_tree_add_51_79_groupi_n_3522 ,csa_tree_add_51_79_groupi_n_2675 ,csa_tree_add_51_79_groupi_n_712);
  or csa_tree_add_51_79_groupi_g42489(csa_tree_add_51_79_groupi_n_3521 ,csa_tree_add_51_79_groupi_n_2153 ,csa_tree_add_51_79_groupi_n_658);
  or csa_tree_add_51_79_groupi_g42490(csa_tree_add_51_79_groupi_n_3520 ,csa_tree_add_51_79_groupi_n_2278 ,csa_tree_add_51_79_groupi_n_1387);
  or csa_tree_add_51_79_groupi_g42491(csa_tree_add_51_79_groupi_n_3519 ,csa_tree_add_51_79_groupi_n_2585 ,csa_tree_add_51_79_groupi_n_1414);
  or csa_tree_add_51_79_groupi_g42492(csa_tree_add_51_79_groupi_n_3518 ,csa_tree_add_51_79_groupi_n_2643 ,csa_tree_add_51_79_groupi_n_1240);
  or csa_tree_add_51_79_groupi_g42493(csa_tree_add_51_79_groupi_n_3517 ,csa_tree_add_51_79_groupi_n_2591 ,csa_tree_add_51_79_groupi_n_1228);
  or csa_tree_add_51_79_groupi_g42494(csa_tree_add_51_79_groupi_n_3516 ,csa_tree_add_51_79_groupi_n_2151 ,csa_tree_add_51_79_groupi_n_1369);
  or csa_tree_add_51_79_groupi_g42495(csa_tree_add_51_79_groupi_n_3515 ,csa_tree_add_51_79_groupi_n_2659 ,csa_tree_add_51_79_groupi_n_1324);
  or csa_tree_add_51_79_groupi_g42496(csa_tree_add_51_79_groupi_n_3514 ,csa_tree_add_51_79_groupi_n_2240 ,csa_tree_add_51_79_groupi_n_1354);
  or csa_tree_add_51_79_groupi_g42497(csa_tree_add_51_79_groupi_n_3513 ,csa_tree_add_51_79_groupi_n_2313 ,csa_tree_add_51_79_groupi_n_739);
  or csa_tree_add_51_79_groupi_g42498(csa_tree_add_51_79_groupi_n_3512 ,csa_tree_add_51_79_groupi_n_2178 ,csa_tree_add_51_79_groupi_n_676);
  nor csa_tree_add_51_79_groupi_g42499(csa_tree_add_51_79_groupi_n_3511 ,csa_tree_add_51_79_groupi_n_1742 ,csa_tree_add_51_79_groupi_n_2381);
  or csa_tree_add_51_79_groupi_g42500(csa_tree_add_51_79_groupi_n_3510 ,csa_tree_add_51_79_groupi_n_2063 ,csa_tree_add_51_79_groupi_n_730);
  or csa_tree_add_51_79_groupi_g42501(csa_tree_add_51_79_groupi_n_3509 ,csa_tree_add_51_79_groupi_n_2134 ,csa_tree_add_51_79_groupi_n_1219);
  or csa_tree_add_51_79_groupi_g42502(csa_tree_add_51_79_groupi_n_3508 ,csa_tree_add_51_79_groupi_n_2194 ,csa_tree_add_51_79_groupi_n_1231);
  or csa_tree_add_51_79_groupi_g42503(csa_tree_add_51_79_groupi_n_3507 ,csa_tree_add_51_79_groupi_n_2112 ,csa_tree_add_51_79_groupi_n_1438);
  or csa_tree_add_51_79_groupi_g42504(csa_tree_add_51_79_groupi_n_3506 ,csa_tree_add_51_79_groupi_n_2251 ,csa_tree_add_51_79_groupi_n_1321);
  or csa_tree_add_51_79_groupi_g42505(csa_tree_add_51_79_groupi_n_3505 ,csa_tree_add_51_79_groupi_n_2572 ,csa_tree_add_51_79_groupi_n_1381);
  or csa_tree_add_51_79_groupi_g42506(csa_tree_add_51_79_groupi_n_3504 ,csa_tree_add_51_79_groupi_n_2216 ,csa_tree_add_51_79_groupi_n_1300);
  or csa_tree_add_51_79_groupi_g42507(csa_tree_add_51_79_groupi_n_3503 ,csa_tree_add_51_79_groupi_n_2792 ,csa_tree_add_51_79_groupi_n_1357);
  or csa_tree_add_51_79_groupi_g42508(csa_tree_add_51_79_groupi_n_3502 ,csa_tree_add_51_79_groupi_n_2782 ,csa_tree_add_51_79_groupi_n_682);
  or csa_tree_add_51_79_groupi_g42509(csa_tree_add_51_79_groupi_n_3501 ,csa_tree_add_51_79_groupi_n_2173 ,csa_tree_add_51_79_groupi_n_1426);
  or csa_tree_add_51_79_groupi_g42510(csa_tree_add_51_79_groupi_n_3500 ,csa_tree_add_51_79_groupi_n_2793 ,csa_tree_add_51_79_groupi_n_1327);
  or csa_tree_add_51_79_groupi_g42511(csa_tree_add_51_79_groupi_n_3499 ,csa_tree_add_51_79_groupi_n_2184 ,csa_tree_add_51_79_groupi_n_1282);
  or csa_tree_add_51_79_groupi_g42512(csa_tree_add_51_79_groupi_n_3498 ,csa_tree_add_51_79_groupi_n_2310 ,csa_tree_add_51_79_groupi_n_1279);
  or csa_tree_add_51_79_groupi_g42513(csa_tree_add_51_79_groupi_n_3497 ,csa_tree_add_51_79_groupi_n_2612 ,csa_tree_add_51_79_groupi_n_1216);
  or csa_tree_add_51_79_groupi_g42514(csa_tree_add_51_79_groupi_n_3496 ,csa_tree_add_51_79_groupi_n_2822 ,csa_tree_add_51_79_groupi_n_1405);
  or csa_tree_add_51_79_groupi_g42515(csa_tree_add_51_79_groupi_n_3495 ,csa_tree_add_51_79_groupi_n_2041 ,csa_tree_add_51_79_groupi_n_1276);
  or csa_tree_add_51_79_groupi_g42516(csa_tree_add_51_79_groupi_n_3494 ,csa_tree_add_51_79_groupi_n_2019 ,csa_tree_add_51_79_groupi_n_1279);
  nor csa_tree_add_51_79_groupi_g42517(csa_tree_add_51_79_groupi_n_3493 ,csa_tree_add_51_79_groupi_n_1724 ,csa_tree_add_51_79_groupi_n_2383);
  or csa_tree_add_51_79_groupi_g42518(csa_tree_add_51_79_groupi_n_3492 ,csa_tree_add_51_79_groupi_n_2094 ,csa_tree_add_51_79_groupi_n_1390);
  or csa_tree_add_51_79_groupi_g42519(csa_tree_add_51_79_groupi_n_3491 ,csa_tree_add_51_79_groupi_n_2031 ,csa_tree_add_51_79_groupi_n_1306);
  or csa_tree_add_51_79_groupi_g42520(csa_tree_add_51_79_groupi_n_3490 ,csa_tree_add_51_79_groupi_n_2245 ,csa_tree_add_51_79_groupi_n_1285);
  or csa_tree_add_51_79_groupi_g42521(csa_tree_add_51_79_groupi_n_3489 ,csa_tree_add_51_79_groupi_n_2778 ,csa_tree_add_51_79_groupi_n_724);
  or csa_tree_add_51_79_groupi_g42522(csa_tree_add_51_79_groupi_n_3488 ,csa_tree_add_51_79_groupi_n_2874 ,csa_tree_add_51_79_groupi_n_1408);
  or csa_tree_add_51_79_groupi_g42523(csa_tree_add_51_79_groupi_n_3487 ,csa_tree_add_51_79_groupi_n_2844 ,csa_tree_add_51_79_groupi_n_1423);
  or csa_tree_add_51_79_groupi_g42524(csa_tree_add_51_79_groupi_n_3486 ,csa_tree_add_51_79_groupi_n_2853 ,csa_tree_add_51_79_groupi_n_1324);
  or csa_tree_add_51_79_groupi_g42525(csa_tree_add_51_79_groupi_n_3485 ,csa_tree_add_51_79_groupi_n_2743 ,csa_tree_add_51_79_groupi_n_1336);
  or csa_tree_add_51_79_groupi_g42526(csa_tree_add_51_79_groupi_n_3484 ,csa_tree_add_51_79_groupi_n_2033 ,csa_tree_add_51_79_groupi_n_1345);
  or csa_tree_add_51_79_groupi_g42527(csa_tree_add_51_79_groupi_n_3483 ,csa_tree_add_51_79_groupi_n_2271 ,csa_tree_add_51_79_groupi_n_1234);
  or csa_tree_add_51_79_groupi_g42528(csa_tree_add_51_79_groupi_n_3482 ,csa_tree_add_51_79_groupi_n_2750 ,csa_tree_add_51_79_groupi_n_1396);
  nor csa_tree_add_51_79_groupi_g42529(csa_tree_add_51_79_groupi_n_3481 ,csa_tree_add_51_79_groupi_n_1758 ,csa_tree_add_51_79_groupi_n_2380);
  or csa_tree_add_51_79_groupi_g42530(csa_tree_add_51_79_groupi_n_3480 ,csa_tree_add_51_79_groupi_n_2034 ,csa_tree_add_51_79_groupi_n_1363);
  or csa_tree_add_51_79_groupi_g42531(csa_tree_add_51_79_groupi_n_3479 ,csa_tree_add_51_79_groupi_n_2838 ,csa_tree_add_51_79_groupi_n_1411);
  or csa_tree_add_51_79_groupi_g42532(csa_tree_add_51_79_groupi_n_3478 ,csa_tree_add_51_79_groupi_n_2725 ,csa_tree_add_51_79_groupi_n_736);
  nor csa_tree_add_51_79_groupi_g42533(csa_tree_add_51_79_groupi_n_3477 ,csa_tree_add_51_79_groupi_n_1678 ,csa_tree_add_51_79_groupi_n_2426);
  nor csa_tree_add_51_79_groupi_g42534(csa_tree_add_51_79_groupi_n_3476 ,csa_tree_add_51_79_groupi_n_1681 ,csa_tree_add_51_79_groupi_n_2425);
  nor csa_tree_add_51_79_groupi_g42535(csa_tree_add_51_79_groupi_n_3475 ,csa_tree_add_51_79_groupi_n_1723 ,csa_tree_add_51_79_groupi_n_2400);
  or csa_tree_add_51_79_groupi_g42536(csa_tree_add_51_79_groupi_n_3474 ,csa_tree_add_51_79_groupi_n_2798 ,csa_tree_add_51_79_groupi_n_1309);
  or csa_tree_add_51_79_groupi_g42537(csa_tree_add_51_79_groupi_n_3473 ,csa_tree_add_51_79_groupi_n_2307 ,csa_tree_add_51_79_groupi_n_1348);
  nor csa_tree_add_51_79_groupi_g42538(csa_tree_add_51_79_groupi_n_3472 ,csa_tree_add_51_79_groupi_n_1700 ,csa_tree_add_51_79_groupi_n_2428);
  nor csa_tree_add_51_79_groupi_g42539(csa_tree_add_51_79_groupi_n_3471 ,csa_tree_add_51_79_groupi_n_1697 ,csa_tree_add_51_79_groupi_n_2424);
  or csa_tree_add_51_79_groupi_g42540(csa_tree_add_51_79_groupi_n_3470 ,csa_tree_add_51_79_groupi_n_2553 ,csa_tree_add_51_79_groupi_n_2554);
  nor csa_tree_add_51_79_groupi_g42541(csa_tree_add_51_79_groupi_n_3469 ,csa_tree_add_51_79_groupi_n_1754 ,csa_tree_add_51_79_groupi_n_2404);
  or csa_tree_add_51_79_groupi_g42542(csa_tree_add_51_79_groupi_n_3468 ,csa_tree_add_51_79_groupi_n_2682 ,csa_tree_add_51_79_groupi_n_1273);
  or csa_tree_add_51_79_groupi_g42543(csa_tree_add_51_79_groupi_n_3467 ,csa_tree_add_51_79_groupi_n_2259 ,csa_tree_add_51_79_groupi_n_658);
  nor csa_tree_add_51_79_groupi_g42544(csa_tree_add_51_79_groupi_n_3466 ,csa_tree_add_51_79_groupi_n_1729 ,csa_tree_add_51_79_groupi_n_2405);
  or csa_tree_add_51_79_groupi_g42545(csa_tree_add_51_79_groupi_n_3465 ,csa_tree_add_51_79_groupi_n_2102 ,csa_tree_add_51_79_groupi_n_1222);
  or csa_tree_add_51_79_groupi_g42546(csa_tree_add_51_79_groupi_n_3464 ,csa_tree_add_51_79_groupi_n_2183 ,csa_tree_add_51_79_groupi_n_1417);
  nor csa_tree_add_51_79_groupi_g42547(csa_tree_add_51_79_groupi_n_3463 ,csa_tree_add_51_79_groupi_n_1737 ,csa_tree_add_51_79_groupi_n_2420);
  or csa_tree_add_51_79_groupi_g42548(csa_tree_add_51_79_groupi_n_3462 ,csa_tree_add_51_79_groupi_n_2277 ,csa_tree_add_51_79_groupi_n_1432);
  or csa_tree_add_51_79_groupi_g42549(csa_tree_add_51_79_groupi_n_3461 ,csa_tree_add_51_79_groupi_n_2808 ,csa_tree_add_51_79_groupi_n_1351);
  or csa_tree_add_51_79_groupi_g42550(csa_tree_add_51_79_groupi_n_3460 ,csa_tree_add_51_79_groupi_n_2130 ,csa_tree_add_51_79_groupi_n_1249);
  or csa_tree_add_51_79_groupi_g42551(csa_tree_add_51_79_groupi_n_3459 ,csa_tree_add_51_79_groupi_n_2710 ,csa_tree_add_51_79_groupi_n_1213);
  or csa_tree_add_51_79_groupi_g42552(csa_tree_add_51_79_groupi_n_3458 ,csa_tree_add_51_79_groupi_n_2639 ,csa_tree_add_51_79_groupi_n_1267);
  or csa_tree_add_51_79_groupi_g42553(csa_tree_add_51_79_groupi_n_3457 ,csa_tree_add_51_79_groupi_n_2182 ,csa_tree_add_51_79_groupi_n_1282);
  or csa_tree_add_51_79_groupi_g42554(csa_tree_add_51_79_groupi_n_3456 ,csa_tree_add_51_79_groupi_n_2055 ,csa_tree_add_51_79_groupi_n_1342);
  or csa_tree_add_51_79_groupi_g42555(csa_tree_add_51_79_groupi_n_3455 ,csa_tree_add_51_79_groupi_n_2152 ,csa_tree_add_51_79_groupi_n_658);
  or csa_tree_add_51_79_groupi_g42556(csa_tree_add_51_79_groupi_n_3454 ,csa_tree_add_51_79_groupi_n_2804 ,csa_tree_add_51_79_groupi_n_736);
  or csa_tree_add_51_79_groupi_g42557(csa_tree_add_51_79_groupi_n_3453 ,csa_tree_add_51_79_groupi_n_2847 ,csa_tree_add_51_79_groupi_n_1402);
  or csa_tree_add_51_79_groupi_g42558(csa_tree_add_51_79_groupi_n_3452 ,csa_tree_add_51_79_groupi_n_2196 ,csa_tree_add_51_79_groupi_n_700);
  or csa_tree_add_51_79_groupi_g42559(csa_tree_add_51_79_groupi_n_3451 ,csa_tree_add_51_79_groupi_n_2261 ,csa_tree_add_51_79_groupi_n_1285);
  or csa_tree_add_51_79_groupi_g42560(csa_tree_add_51_79_groupi_n_3450 ,csa_tree_add_51_79_groupi_n_2752 ,csa_tree_add_51_79_groupi_n_685);
  or csa_tree_add_51_79_groupi_g42561(csa_tree_add_51_79_groupi_n_3449 ,csa_tree_add_51_79_groupi_n_2845 ,csa_tree_add_51_79_groupi_n_1333);
  or csa_tree_add_51_79_groupi_g42562(csa_tree_add_51_79_groupi_n_3448 ,csa_tree_add_51_79_groupi_n_2158 ,csa_tree_add_51_79_groupi_n_697);
  or csa_tree_add_51_79_groupi_g42563(csa_tree_add_51_79_groupi_n_3447 ,csa_tree_add_51_79_groupi_n_2708 ,csa_tree_add_51_79_groupi_n_1366);
  or csa_tree_add_51_79_groupi_g42564(csa_tree_add_51_79_groupi_n_3446 ,csa_tree_add_51_79_groupi_n_2768 ,csa_tree_add_51_79_groupi_n_1399);
  or csa_tree_add_51_79_groupi_g42565(csa_tree_add_51_79_groupi_n_3445 ,csa_tree_add_51_79_groupi_n_2136 ,csa_tree_add_51_79_groupi_n_1438);
  or csa_tree_add_51_79_groupi_g42566(csa_tree_add_51_79_groupi_n_3444 ,csa_tree_add_51_79_groupi_n_2200 ,csa_tree_add_51_79_groupi_n_1282);
  or csa_tree_add_51_79_groupi_g42567(csa_tree_add_51_79_groupi_n_3443 ,csa_tree_add_51_79_groupi_n_2244 ,csa_tree_add_51_79_groupi_n_1372);
  or csa_tree_add_51_79_groupi_g42568(csa_tree_add_51_79_groupi_n_3442 ,csa_tree_add_51_79_groupi_n_2103 ,csa_tree_add_51_79_groupi_n_1306);
  or csa_tree_add_51_79_groupi_g42569(csa_tree_add_51_79_groupi_n_3441 ,csa_tree_add_51_79_groupi_n_2707 ,csa_tree_add_51_79_groupi_n_1444);
  or csa_tree_add_51_79_groupi_g42570(csa_tree_add_51_79_groupi_n_3440 ,csa_tree_add_51_79_groupi_n_2236 ,csa_tree_add_51_79_groupi_n_1318);
  or csa_tree_add_51_79_groupi_g42571(csa_tree_add_51_79_groupi_n_3439 ,csa_tree_add_51_79_groupi_n_2718 ,csa_tree_add_51_79_groupi_n_730);
  or csa_tree_add_51_79_groupi_g42572(csa_tree_add_51_79_groupi_n_3438 ,csa_tree_add_51_79_groupi_n_2586 ,csa_tree_add_51_79_groupi_n_1267);
  or csa_tree_add_51_79_groupi_g42573(csa_tree_add_51_79_groupi_n_3437 ,csa_tree_add_51_79_groupi_n_2638 ,csa_tree_add_51_79_groupi_n_1384);
  or csa_tree_add_51_79_groupi_g42574(csa_tree_add_51_79_groupi_n_3436 ,csa_tree_add_51_79_groupi_n_2802 ,csa_tree_add_51_79_groupi_n_1216);
  or csa_tree_add_51_79_groupi_g42575(csa_tree_add_51_79_groupi_n_3435 ,csa_tree_add_51_79_groupi_n_2163 ,csa_tree_add_51_79_groupi_n_1219);
  or csa_tree_add_51_79_groupi_g42576(csa_tree_add_51_79_groupi_n_3434 ,csa_tree_add_51_79_groupi_n_2593 ,csa_tree_add_51_79_groupi_n_1375);
  or csa_tree_add_51_79_groupi_g42577(csa_tree_add_51_79_groupi_n_3433 ,csa_tree_add_51_79_groupi_n_2197 ,csa_tree_add_51_79_groupi_n_1321);
  or csa_tree_add_51_79_groupi_g42578(csa_tree_add_51_79_groupi_n_3432 ,csa_tree_add_51_79_groupi_n_2243 ,csa_tree_add_51_79_groupi_n_1090);
  or csa_tree_add_51_79_groupi_g42579(csa_tree_add_51_79_groupi_n_3431 ,csa_tree_add_51_79_groupi_n_2582 ,csa_tree_add_51_79_groupi_n_1378);
  or csa_tree_add_51_79_groupi_g42580(csa_tree_add_51_79_groupi_n_3430 ,csa_tree_add_51_79_groupi_n_2270 ,csa_tree_add_51_79_groupi_n_1231);
  or csa_tree_add_51_79_groupi_g42581(csa_tree_add_51_79_groupi_n_3429 ,csa_tree_add_51_79_groupi_n_2221 ,csa_tree_add_51_79_groupi_n_1243);
  or csa_tree_add_51_79_groupi_g42582(csa_tree_add_51_79_groupi_n_3428 ,csa_tree_add_51_79_groupi_n_2064 ,csa_tree_add_51_79_groupi_n_1435);
  or csa_tree_add_51_79_groupi_g42583(csa_tree_add_51_79_groupi_n_3427 ,csa_tree_add_51_79_groupi_n_2664 ,csa_tree_add_51_79_groupi_n_1101);
  or csa_tree_add_51_79_groupi_g42584(csa_tree_add_51_79_groupi_n_3426 ,csa_tree_add_51_79_groupi_n_2039 ,csa_tree_add_51_79_groupi_n_1354);
  or csa_tree_add_51_79_groupi_g42585(csa_tree_add_51_79_groupi_n_3425 ,csa_tree_add_51_79_groupi_n_2865 ,csa_tree_add_51_79_groupi_n_1420);
  or csa_tree_add_51_79_groupi_g42586(csa_tree_add_51_79_groupi_n_3424 ,csa_tree_add_51_79_groupi_n_1783 ,csa_tree_add_51_79_groupi_n_2415);
  or csa_tree_add_51_79_groupi_g42587(csa_tree_add_51_79_groupi_n_3423 ,csa_tree_add_51_79_groupi_n_2045 ,csa_tree_add_51_79_groupi_n_1405);
  or csa_tree_add_51_79_groupi_g42588(csa_tree_add_51_79_groupi_n_3422 ,csa_tree_add_51_79_groupi_n_2074 ,csa_tree_add_51_79_groupi_n_724);
  or csa_tree_add_51_79_groupi_g42589(csa_tree_add_51_79_groupi_n_3421 ,csa_tree_add_51_79_groupi_n_2069 ,csa_tree_add_51_79_groupi_n_1273);
  or csa_tree_add_51_79_groupi_g42590(csa_tree_add_51_79_groupi_n_3420 ,csa_tree_add_51_79_groupi_n_2247 ,csa_tree_add_51_79_groupi_n_1303);
  or csa_tree_add_51_79_groupi_g42591(csa_tree_add_51_79_groupi_n_3419 ,csa_tree_add_51_79_groupi_n_2732 ,csa_tree_add_51_79_groupi_n_712);
  or csa_tree_add_51_79_groupi_g42592(csa_tree_add_51_79_groupi_n_3418 ,csa_tree_add_51_79_groupi_n_2730 ,csa_tree_add_51_79_groupi_n_1444);
  or csa_tree_add_51_79_groupi_g42593(csa_tree_add_51_79_groupi_n_3417 ,csa_tree_add_51_79_groupi_n_2672 ,csa_tree_add_51_79_groupi_n_1393);
  or csa_tree_add_51_79_groupi_g42594(csa_tree_add_51_79_groupi_n_3416 ,csa_tree_add_51_79_groupi_n_2690 ,csa_tree_add_51_79_groupi_n_1396);
  or csa_tree_add_51_79_groupi_g42595(csa_tree_add_51_79_groupi_n_3415 ,csa_tree_add_51_79_groupi_n_2280 ,csa_tree_add_51_79_groupi_n_1432);
  or csa_tree_add_51_79_groupi_g42596(csa_tree_add_51_79_groupi_n_3414 ,csa_tree_add_51_79_groupi_n_2141 ,csa_tree_add_51_79_groupi_n_1408);
  or csa_tree_add_51_79_groupi_g42597(csa_tree_add_51_79_groupi_n_3413 ,csa_tree_add_51_79_groupi_n_2788 ,csa_tree_add_51_79_groupi_n_1288);
  or csa_tree_add_51_79_groupi_g42598(csa_tree_add_51_79_groupi_n_3412 ,csa_tree_add_51_79_groupi_n_2275 ,csa_tree_add_51_79_groupi_n_751);
  or csa_tree_add_51_79_groupi_g42599(csa_tree_add_51_79_groupi_n_3411 ,csa_tree_add_51_79_groupi_n_2289 ,csa_tree_add_51_79_groupi_n_1330);
  or csa_tree_add_51_79_groupi_g42600(csa_tree_add_51_79_groupi_n_3410 ,csa_tree_add_51_79_groupi_n_2872 ,csa_tree_add_51_79_groupi_n_1429);
  or csa_tree_add_51_79_groupi_g42601(csa_tree_add_51_79_groupi_n_3409 ,csa_tree_add_51_79_groupi_n_2296 ,csa_tree_add_51_79_groupi_n_1405);
  nor csa_tree_add_51_79_groupi_g42602(csa_tree_add_51_79_groupi_n_3408 ,csa_tree_add_51_79_groupi_n_1694 ,csa_tree_add_51_79_groupi_n_2397);
  nor csa_tree_add_51_79_groupi_g42603(csa_tree_add_51_79_groupi_n_3407 ,csa_tree_add_51_79_groupi_n_1747 ,csa_tree_add_51_79_groupi_n_2414);
  nor csa_tree_add_51_79_groupi_g42604(csa_tree_add_51_79_groupi_n_3406 ,csa_tree_add_51_79_groupi_n_1699 ,csa_tree_add_51_79_groupi_n_2382);
  or csa_tree_add_51_79_groupi_g42605(csa_tree_add_51_79_groupi_n_3405 ,csa_tree_add_51_79_groupi_n_2871 ,csa_tree_add_51_79_groupi_n_751);
  or csa_tree_add_51_79_groupi_g42606(csa_tree_add_51_79_groupi_n_3404 ,csa_tree_add_51_79_groupi_n_2171 ,csa_tree_add_51_79_groupi_n_709);
  or csa_tree_add_51_79_groupi_g42607(csa_tree_add_51_79_groupi_n_3403 ,csa_tree_add_51_79_groupi_n_2239 ,csa_tree_add_51_79_groupi_n_1231);
  or csa_tree_add_51_79_groupi_g42608(csa_tree_add_51_79_groupi_n_3402 ,csa_tree_add_51_79_groupi_n_2204 ,csa_tree_add_51_79_groupi_n_700);
  or csa_tree_add_51_79_groupi_g42609(csa_tree_add_51_79_groupi_n_3401 ,csa_tree_add_51_79_groupi_n_2148 ,csa_tree_add_51_79_groupi_n_1369);
  or csa_tree_add_51_79_groupi_g42610(csa_tree_add_51_79_groupi_n_3400 ,csa_tree_add_51_79_groupi_n_2859 ,csa_tree_add_51_79_groupi_n_1252);
  or csa_tree_add_51_79_groupi_g42611(csa_tree_add_51_79_groupi_n_3399 ,csa_tree_add_51_79_groupi_n_2143 ,csa_tree_add_51_79_groupi_n_1243);
  or csa_tree_add_51_79_groupi_g42612(csa_tree_add_51_79_groupi_n_3398 ,csa_tree_add_51_79_groupi_n_2162 ,csa_tree_add_51_79_groupi_n_1300);
  or csa_tree_add_51_79_groupi_g42613(csa_tree_add_51_79_groupi_n_3397 ,csa_tree_add_51_79_groupi_n_2674 ,csa_tree_add_51_79_groupi_n_1216);
  or csa_tree_add_51_79_groupi_g42614(csa_tree_add_51_79_groupi_n_3396 ,csa_tree_add_51_79_groupi_n_2783 ,csa_tree_add_51_79_groupi_n_1096);
  or csa_tree_add_51_79_groupi_g42615(csa_tree_add_51_79_groupi_n_3395 ,csa_tree_add_51_79_groupi_n_2192 ,csa_tree_add_51_79_groupi_n_1273);
  or csa_tree_add_51_79_groupi_g42616(csa_tree_add_51_79_groupi_n_3394 ,csa_tree_add_51_79_groupi_n_2217 ,csa_tree_add_51_79_groupi_n_1258);
  nor csa_tree_add_51_79_groupi_g42617(csa_tree_add_51_79_groupi_n_3393 ,csa_tree_add_51_79_groupi_n_1738 ,csa_tree_add_51_79_groupi_n_2375);
  or csa_tree_add_51_79_groupi_g42618(csa_tree_add_51_79_groupi_n_3392 ,csa_tree_add_51_79_groupi_n_2205 ,csa_tree_add_51_79_groupi_n_1318);
  or csa_tree_add_51_79_groupi_g42619(csa_tree_add_51_79_groupi_n_3391 ,csa_tree_add_51_79_groupi_n_2133 ,csa_tree_add_51_79_groupi_n_1258);
  or csa_tree_add_51_79_groupi_g42620(csa_tree_add_51_79_groupi_n_3390 ,csa_tree_add_51_79_groupi_n_2242 ,csa_tree_add_51_79_groupi_n_658);
  nor csa_tree_add_51_79_groupi_g42621(csa_tree_add_51_79_groupi_n_3389 ,csa_tree_add_51_79_groupi_n_2543 ,csa_tree_add_51_79_groupi_n_2545);
  or csa_tree_add_51_79_groupi_g42622(csa_tree_add_51_79_groupi_n_3388 ,csa_tree_add_51_79_groupi_n_2833 ,csa_tree_add_51_79_groupi_n_1381);
  or csa_tree_add_51_79_groupi_g42623(csa_tree_add_51_79_groupi_n_3387 ,csa_tree_add_51_79_groupi_n_2702 ,csa_tree_add_51_79_groupi_n_745);
  or csa_tree_add_51_79_groupi_g42624(csa_tree_add_51_79_groupi_n_3386 ,csa_tree_add_51_79_groupi_n_2860 ,csa_tree_add_51_79_groupi_n_1345);
  or csa_tree_add_51_79_groupi_g42625(csa_tree_add_51_79_groupi_n_3385 ,csa_tree_add_51_79_groupi_n_2746 ,csa_tree_add_51_79_groupi_n_1414);
  or csa_tree_add_51_79_groupi_g42626(csa_tree_add_51_79_groupi_n_3384 ,csa_tree_add_51_79_groupi_n_2042 ,csa_tree_add_51_79_groupi_n_1103);
  or csa_tree_add_51_79_groupi_g42627(csa_tree_add_51_79_groupi_n_3383 ,csa_tree_add_51_79_groupi_n_2628 ,csa_tree_add_51_79_groupi_n_1438);
  nor csa_tree_add_51_79_groupi_g42628(csa_tree_add_51_79_groupi_n_3382 ,csa_tree_add_51_79_groupi_n_1679 ,csa_tree_add_51_79_groupi_n_2408);
  nor csa_tree_add_51_79_groupi_g42629(csa_tree_add_51_79_groupi_n_3381 ,csa_tree_add_51_79_groupi_n_1759 ,csa_tree_add_51_79_groupi_n_2433);
  or csa_tree_add_51_79_groupi_g42630(csa_tree_add_51_79_groupi_n_3380 ,csa_tree_add_51_79_groupi_n_2740 ,csa_tree_add_51_79_groupi_n_1255);
  or csa_tree_add_51_79_groupi_g42631(csa_tree_add_51_79_groupi_n_3379 ,csa_tree_add_51_79_groupi_n_2805 ,csa_tree_add_51_79_groupi_n_2478);
  or csa_tree_add_51_79_groupi_g42632(csa_tree_add_51_79_groupi_n_3378 ,csa_tree_add_51_79_groupi_n_2129 ,csa_tree_add_51_79_groupi_n_1098);
  or csa_tree_add_51_79_groupi_g42633(csa_tree_add_51_79_groupi_n_3377 ,csa_tree_add_51_79_groupi_n_2856 ,csa_tree_add_51_79_groupi_n_1360);
  or csa_tree_add_51_79_groupi_g42634(csa_tree_add_51_79_groupi_n_3376 ,csa_tree_add_51_79_groupi_n_2551 ,csa_tree_add_51_79_groupi_n_2549);
  and csa_tree_add_51_79_groupi_g42635(csa_tree_add_51_79_groupi_n_3375 ,csa_tree_add_51_79_groupi_n_2544 ,csa_tree_add_51_79_groupi_n_2547);
  or csa_tree_add_51_79_groupi_g42636(csa_tree_add_51_79_groupi_n_3374 ,csa_tree_add_51_79_groupi_n_2742 ,csa_tree_add_51_79_groupi_n_1092);
  or csa_tree_add_51_79_groupi_g42637(csa_tree_add_51_79_groupi_n_3872 ,csa_tree_add_51_79_groupi_n_2757 ,csa_tree_add_51_79_groupi_n_2466);
  and csa_tree_add_51_79_groupi_g42638(csa_tree_add_51_79_groupi_n_3870 ,csa_tree_add_51_79_groupi_n_2228 ,csa_tree_add_51_79_groupi_n_2487);
  or csa_tree_add_51_79_groupi_g42639(csa_tree_add_51_79_groupi_n_3869 ,csa_tree_add_51_79_groupi_n_2790 ,csa_tree_add_51_79_groupi_n_2457);
  or csa_tree_add_51_79_groupi_g42640(csa_tree_add_51_79_groupi_n_3868 ,csa_tree_add_51_79_groupi_n_2762 ,csa_tree_add_51_79_groupi_n_1363);
  and csa_tree_add_51_79_groupi_g42641(csa_tree_add_51_79_groupi_n_3866 ,csa_tree_add_51_79_groupi_n_2201 ,csa_tree_add_51_79_groupi_n_2434);
  or csa_tree_add_51_79_groupi_g42642(csa_tree_add_51_79_groupi_n_3865 ,csa_tree_add_51_79_groupi_n_2882 ,csa_tree_add_51_79_groupi_n_1348);
  or csa_tree_add_51_79_groupi_g42643(csa_tree_add_51_79_groupi_n_3864 ,csa_tree_add_51_79_groupi_n_2046 ,csa_tree_add_51_79_groupi_n_1970);
  or csa_tree_add_51_79_groupi_g42644(csa_tree_add_51_79_groupi_n_3863 ,csa_tree_add_51_79_groupi_n_2234 ,csa_tree_add_51_79_groupi_n_1099);
  or csa_tree_add_51_79_groupi_g42645(csa_tree_add_51_79_groupi_n_3862 ,csa_tree_add_51_79_groupi_n_2706 ,csa_tree_add_51_79_groupi_n_1333);
  or csa_tree_add_51_79_groupi_g42646(csa_tree_add_51_79_groupi_n_3861 ,csa_tree_add_51_79_groupi_n_2267 ,csa_tree_add_51_79_groupi_n_2497);
  or csa_tree_add_51_79_groupi_g42647(csa_tree_add_51_79_groupi_n_3860 ,csa_tree_add_51_79_groupi_n_592 ,csa_tree_add_51_79_groupi_n_2059);
  or csa_tree_add_51_79_groupi_g42648(csa_tree_add_51_79_groupi_n_3859 ,csa_tree_add_51_79_groupi_n_2607 ,csa_tree_add_51_79_groupi_n_1441);
  and csa_tree_add_51_79_groupi_g42649(csa_tree_add_51_79_groupi_n_3857 ,csa_tree_add_51_79_groupi_n_2166 ,csa_tree_add_51_79_groupi_n_2501);
  or csa_tree_add_51_79_groupi_g42650(csa_tree_add_51_79_groupi_n_3856 ,csa_tree_add_51_79_groupi_n_2617 ,csa_tree_add_51_79_groupi_n_1342);
  and csa_tree_add_51_79_groupi_g42651(csa_tree_add_51_79_groupi_n_3854 ,csa_tree_add_51_79_groupi_n_2772 ,csa_tree_add_51_79_groupi_n_1985);
  or csa_tree_add_51_79_groupi_g42652(csa_tree_add_51_79_groupi_n_3853 ,csa_tree_add_51_79_groupi_n_600 ,csa_tree_add_51_79_groupi_n_2759);
  or csa_tree_add_51_79_groupi_g42653(csa_tree_add_51_79_groupi_n_3852 ,csa_tree_add_51_79_groupi_n_2065 ,csa_tree_add_51_79_groupi_n_1294);
  or csa_tree_add_51_79_groupi_g42654(csa_tree_add_51_79_groupi_n_3851 ,csa_tree_add_51_79_groupi_n_2693 ,csa_tree_add_51_79_groupi_n_1111);
  and csa_tree_add_51_79_groupi_g42655(csa_tree_add_51_79_groupi_n_3849 ,csa_tree_add_51_79_groupi_n_2023 ,csa_tree_add_51_79_groupi_n_1989);
  or csa_tree_add_51_79_groupi_g42656(csa_tree_add_51_79_groupi_n_3848 ,csa_tree_add_51_79_groupi_n_2286 ,csa_tree_add_51_79_groupi_n_1435);
  and csa_tree_add_51_79_groupi_g42657(csa_tree_add_51_79_groupi_n_3846 ,csa_tree_add_51_79_groupi_n_2794 ,csa_tree_add_51_79_groupi_n_2511);
  or csa_tree_add_51_79_groupi_g42658(csa_tree_add_51_79_groupi_n_3845 ,csa_tree_add_51_79_groupi_n_2575 ,csa_tree_add_51_79_groupi_n_1366);
  or csa_tree_add_51_79_groupi_g42659(csa_tree_add_51_79_groupi_n_3844 ,csa_tree_add_51_79_groupi_n_871 ,csa_tree_add_51_79_groupi_n_2635);
  or csa_tree_add_51_79_groupi_g42660(csa_tree_add_51_79_groupi_n_3843 ,csa_tree_add_51_79_groupi_n_530 ,csa_tree_add_51_79_groupi_n_2671);
  or csa_tree_add_51_79_groupi_g42661(csa_tree_add_51_79_groupi_n_3842 ,csa_tree_add_51_79_groupi_n_2097 ,csa_tree_add_51_79_groupi_n_1995);
  or csa_tree_add_51_79_groupi_g42662(csa_tree_add_51_79_groupi_n_3841 ,csa_tree_add_51_79_groupi_n_551 ,csa_tree_add_51_79_groupi_n_2858);
  or csa_tree_add_51_79_groupi_g42663(csa_tree_add_51_79_groupi_n_3840 ,csa_tree_add_51_79_groupi_n_597 ,csa_tree_add_51_79_groupi_n_2027);
  or csa_tree_add_51_79_groupi_g42664(csa_tree_add_51_79_groupi_n_3839 ,csa_tree_add_51_79_groupi_n_864 ,csa_tree_add_51_79_groupi_n_2601);
  or csa_tree_add_51_79_groupi_g42665(csa_tree_add_51_79_groupi_n_3838 ,csa_tree_add_51_79_groupi_n_556 ,csa_tree_add_51_79_groupi_n_2603);
  or csa_tree_add_51_79_groupi_g42666(csa_tree_add_51_79_groupi_n_3837 ,csa_tree_add_51_79_groupi_n_543 ,csa_tree_add_51_79_groupi_n_2111);
  or csa_tree_add_51_79_groupi_g42667(csa_tree_add_51_79_groupi_n_3836 ,csa_tree_add_51_79_groupi_n_525 ,csa_tree_add_51_79_groupi_n_2653);
  or csa_tree_add_51_79_groupi_g42668(csa_tree_add_51_79_groupi_n_3835 ,csa_tree_add_51_79_groupi_n_535 ,csa_tree_add_51_79_groupi_n_2168);
  or csa_tree_add_51_79_groupi_g42669(csa_tree_add_51_79_groupi_n_3834 ,csa_tree_add_51_79_groupi_n_888 ,csa_tree_add_51_79_groupi_n_2611);
  and csa_tree_add_51_79_groupi_g42670(csa_tree_add_51_79_groupi_n_3833 ,csa_tree_add_51_79_groupi_n_1841 ,csa_tree_add_51_79_groupi_n_1450);
  and csa_tree_add_51_79_groupi_g42671(csa_tree_add_51_79_groupi_n_3832 ,csa_tree_add_51_79_groupi_n_1864 ,csa_tree_add_51_79_groupi_n_727);
  and csa_tree_add_51_79_groupi_g42672(csa_tree_add_51_79_groupi_n_3831 ,csa_tree_add_51_79_groupi_n_1920 ,csa_tree_add_51_79_groupi_n_1462);
  and csa_tree_add_51_79_groupi_g42673(csa_tree_add_51_79_groupi_n_3830 ,csa_tree_add_51_79_groupi_n_1858 ,csa_tree_add_51_79_groupi_n_727);
  and csa_tree_add_51_79_groupi_g42674(csa_tree_add_51_79_groupi_n_3828 ,csa_tree_add_51_79_groupi_n_1894 ,csa_tree_add_51_79_groupi_n_1459);
  and csa_tree_add_51_79_groupi_g42675(csa_tree_add_51_79_groupi_n_3827 ,csa_tree_add_51_79_groupi_n_1879 ,csa_tree_add_51_79_groupi_n_670);
  and csa_tree_add_51_79_groupi_g42676(csa_tree_add_51_79_groupi_n_3825 ,csa_tree_add_51_79_groupi_n_1868 ,csa_tree_add_51_79_groupi_n_1469);
  and csa_tree_add_51_79_groupi_g42677(csa_tree_add_51_79_groupi_n_3823 ,csa_tree_add_51_79_groupi_n_1918 ,csa_tree_add_51_79_groupi_n_1462);
  and csa_tree_add_51_79_groupi_g42678(csa_tree_add_51_79_groupi_n_3821 ,csa_tree_add_51_79_groupi_n_1886 ,csa_tree_add_51_79_groupi_n_1085);
  and csa_tree_add_51_79_groupi_g42679(csa_tree_add_51_79_groupi_n_3819 ,csa_tree_add_51_79_groupi_n_2569 ,csa_tree_add_51_79_groupi_n_2564);
  and csa_tree_add_51_79_groupi_g42680(csa_tree_add_51_79_groupi_n_3817 ,csa_tree_add_51_79_groupi_n_1939 ,csa_tree_add_51_79_groupi_n_2537);
  and csa_tree_add_51_79_groupi_g42681(csa_tree_add_51_79_groupi_n_3815 ,csa_tree_add_51_79_groupi_n_1875 ,csa_tree_add_51_79_groupi_n_1462);
  and csa_tree_add_51_79_groupi_g42682(csa_tree_add_51_79_groupi_n_3813 ,csa_tree_add_51_79_groupi_n_1897 ,csa_tree_add_51_79_groupi_n_2530);
  and csa_tree_add_51_79_groupi_g42683(csa_tree_add_51_79_groupi_n_3812 ,csa_tree_add_51_79_groupi_n_1861 ,csa_tree_add_51_79_groupi_n_1456);
  and csa_tree_add_51_79_groupi_g42684(csa_tree_add_51_79_groupi_n_3810 ,csa_tree_add_51_79_groupi_n_1883 ,csa_tree_add_51_79_groupi_n_718);
  and csa_tree_add_51_79_groupi_g42685(csa_tree_add_51_79_groupi_n_3808 ,csa_tree_add_51_79_groupi_n_1930 ,csa_tree_add_51_79_groupi_n_718);
  and csa_tree_add_51_79_groupi_g42686(csa_tree_add_51_79_groupi_n_3806 ,csa_tree_add_51_79_groupi_n_1941 ,csa_tree_add_51_79_groupi_n_1469);
  and csa_tree_add_51_79_groupi_g42687(csa_tree_add_51_79_groupi_n_3804 ,csa_tree_add_51_79_groupi_n_1839 ,csa_tree_add_51_79_groupi_n_1459);
  and csa_tree_add_51_79_groupi_g42688(csa_tree_add_51_79_groupi_n_3803 ,csa_tree_add_51_79_groupi_n_1963 ,csa_tree_add_51_79_groupi_n_1459);
  and csa_tree_add_51_79_groupi_g42689(csa_tree_add_51_79_groupi_n_3801 ,csa_tree_add_51_79_groupi_n_1842 ,csa_tree_add_51_79_groupi_n_1462);
  and csa_tree_add_51_79_groupi_g42690(csa_tree_add_51_79_groupi_n_3800 ,csa_tree_add_51_79_groupi_n_1937 ,csa_tree_add_51_79_groupi_n_742);
  and csa_tree_add_51_79_groupi_g42691(csa_tree_add_51_79_groupi_n_3799 ,csa_tree_add_51_79_groupi_n_1903 ,csa_tree_add_51_79_groupi_n_1469);
  and csa_tree_add_51_79_groupi_g42692(csa_tree_add_51_79_groupi_n_3797 ,csa_tree_add_51_79_groupi_n_1865 ,csa_tree_add_51_79_groupi_n_742);
  and csa_tree_add_51_79_groupi_g42693(csa_tree_add_51_79_groupi_n_3796 ,csa_tree_add_51_79_groupi_n_1851 ,csa_tree_add_51_79_groupi_n_670);
  and csa_tree_add_51_79_groupi_g42694(csa_tree_add_51_79_groupi_n_3795 ,csa_tree_add_51_79_groupi_n_1840 ,csa_tree_add_51_79_groupi_n_1083);
  and csa_tree_add_51_79_groupi_g42695(csa_tree_add_51_79_groupi_n_3794 ,csa_tree_add_51_79_groupi_n_1857 ,csa_tree_add_51_79_groupi_n_1456);
  and csa_tree_add_51_79_groupi_g42696(csa_tree_add_51_79_groupi_n_3792 ,csa_tree_add_51_79_groupi_n_1935 ,csa_tree_add_51_79_groupi_n_1459);
  and csa_tree_add_51_79_groupi_g42697(csa_tree_add_51_79_groupi_n_3790 ,csa_tree_add_51_79_groupi_n_1936 ,csa_tree_add_51_79_groupi_n_1079);
  and csa_tree_add_51_79_groupi_g42698(csa_tree_add_51_79_groupi_n_3789 ,csa_tree_add_51_79_groupi_n_1846 ,csa_tree_add_51_79_groupi_n_2537);
  and csa_tree_add_51_79_groupi_g42699(csa_tree_add_51_79_groupi_n_3787 ,csa_tree_add_51_79_groupi_n_1889 ,csa_tree_add_51_79_groupi_n_1450);
  and csa_tree_add_51_79_groupi_g42700(csa_tree_add_51_79_groupi_n_3786 ,csa_tree_add_51_79_groupi_n_1906 ,csa_tree_add_51_79_groupi_n_1124);
  and csa_tree_add_51_79_groupi_g42701(csa_tree_add_51_79_groupi_n_3785 ,csa_tree_add_51_79_groupi_n_1856 ,csa_tree_add_51_79_groupi_n_1459);
  and csa_tree_add_51_79_groupi_g42702(csa_tree_add_51_79_groupi_n_3783 ,csa_tree_add_51_79_groupi_n_1869 ,csa_tree_add_51_79_groupi_n_1081);
  and csa_tree_add_51_79_groupi_g42703(csa_tree_add_51_79_groupi_n_3781 ,csa_tree_add_51_79_groupi_n_1904 ,csa_tree_add_51_79_groupi_n_1081);
  and csa_tree_add_51_79_groupi_g42704(csa_tree_add_51_79_groupi_n_3780 ,csa_tree_add_51_79_groupi_n_1929 ,csa_tree_add_51_79_groupi_n_1469);
  and csa_tree_add_51_79_groupi_g42705(csa_tree_add_51_79_groupi_n_3778 ,csa_tree_add_51_79_groupi_n_1873 ,csa_tree_add_51_79_groupi_n_1124);
  and csa_tree_add_51_79_groupi_g42706(csa_tree_add_51_79_groupi_n_3776 ,csa_tree_add_51_79_groupi_n_1834 ,csa_tree_add_51_79_groupi_n_1079);
  and csa_tree_add_51_79_groupi_g42707(csa_tree_add_51_79_groupi_n_3775 ,csa_tree_add_51_79_groupi_n_1849 ,csa_tree_add_51_79_groupi_n_1456);
  and csa_tree_add_51_79_groupi_g42708(csa_tree_add_51_79_groupi_n_3773 ,csa_tree_add_51_79_groupi_n_1831 ,csa_tree_add_51_79_groupi_n_1469);
  and csa_tree_add_51_79_groupi_g42709(csa_tree_add_51_79_groupi_n_3771 ,csa_tree_add_51_79_groupi_n_1913 ,csa_tree_add_51_79_groupi_n_718);
  and csa_tree_add_51_79_groupi_g42710(csa_tree_add_51_79_groupi_n_3769 ,csa_tree_add_51_79_groupi_n_1960 ,csa_tree_add_51_79_groupi_n_718);
  and csa_tree_add_51_79_groupi_g42711(csa_tree_add_51_79_groupi_n_3767 ,csa_tree_add_51_79_groupi_n_1862 ,csa_tree_add_51_79_groupi_n_2530);
  and csa_tree_add_51_79_groupi_g42712(csa_tree_add_51_79_groupi_n_3765 ,csa_tree_add_51_79_groupi_n_1843 ,csa_tree_add_51_79_groupi_n_2537);
  and csa_tree_add_51_79_groupi_g42713(csa_tree_add_51_79_groupi_n_3763 ,csa_tree_add_51_79_groupi_n_1955 ,csa_tree_add_51_79_groupi_n_742);
  and csa_tree_add_51_79_groupi_g42714(csa_tree_add_51_79_groupi_n_3762 ,csa_tree_add_51_79_groupi_n_1835 ,csa_tree_add_51_79_groupi_n_2530);
  and csa_tree_add_51_79_groupi_g42715(csa_tree_add_51_79_groupi_n_3760 ,csa_tree_add_51_79_groupi_n_1914 ,csa_tree_add_51_79_groupi_n_1085);
  and csa_tree_add_51_79_groupi_g42716(csa_tree_add_51_79_groupi_n_3758 ,csa_tree_add_51_79_groupi_n_1854 ,csa_tree_add_51_79_groupi_n_2518);
  and csa_tree_add_51_79_groupi_g42717(csa_tree_add_51_79_groupi_n_3757 ,csa_tree_add_51_79_groupi_n_1859 ,csa_tree_add_51_79_groupi_n_1124);
  and csa_tree_add_51_79_groupi_g42718(csa_tree_add_51_79_groupi_n_3755 ,csa_tree_add_51_79_groupi_n_1945 ,csa_tree_add_51_79_groupi_n_742);
  and csa_tree_add_51_79_groupi_g42719(csa_tree_add_51_79_groupi_n_3753 ,csa_tree_add_51_79_groupi_n_1838 ,csa_tree_add_51_79_groupi_n_1459);
  and csa_tree_add_51_79_groupi_g42720(csa_tree_add_51_79_groupi_n_3752 ,csa_tree_add_51_79_groupi_n_1943 ,csa_tree_add_51_79_groupi_n_1124);
  and csa_tree_add_51_79_groupi_g42721(csa_tree_add_51_79_groupi_n_3750 ,csa_tree_add_51_79_groupi_n_1845 ,csa_tree_add_51_79_groupi_n_1124);
  and csa_tree_add_51_79_groupi_g42722(csa_tree_add_51_79_groupi_n_3748 ,csa_tree_add_51_79_groupi_n_1951 ,csa_tree_add_51_79_groupi_n_2515);
  and csa_tree_add_51_79_groupi_g42723(csa_tree_add_51_79_groupi_n_3746 ,csa_tree_add_51_79_groupi_n_1934 ,csa_tree_add_51_79_groupi_n_1083);
  and csa_tree_add_51_79_groupi_g42724(csa_tree_add_51_79_groupi_n_3744 ,csa_tree_add_51_79_groupi_n_1946 ,csa_tree_add_51_79_groupi_n_742);
  and csa_tree_add_51_79_groupi_g42725(csa_tree_add_51_79_groupi_n_3743 ,csa_tree_add_51_79_groupi_n_1878 ,csa_tree_add_51_79_groupi_n_727);
  and csa_tree_add_51_79_groupi_g42726(csa_tree_add_51_79_groupi_n_3742 ,csa_tree_add_51_79_groupi_n_1885 ,csa_tree_add_51_79_groupi_n_718);
  and csa_tree_add_51_79_groupi_g42727(csa_tree_add_51_79_groupi_n_3740 ,csa_tree_add_51_79_groupi_n_1828 ,csa_tree_add_51_79_groupi_n_1456);
  and csa_tree_add_51_79_groupi_g42728(csa_tree_add_51_79_groupi_n_3739 ,csa_tree_add_51_79_groupi_n_1962 ,csa_tree_add_51_79_groupi_n_670);
  and csa_tree_add_51_79_groupi_g42729(csa_tree_add_51_79_groupi_n_3738 ,csa_tree_add_51_79_groupi_n_1915 ,csa_tree_add_51_79_groupi_n_742);
  and csa_tree_add_51_79_groupi_g42730(csa_tree_add_51_79_groupi_n_3737 ,csa_tree_add_51_79_groupi_n_1942 ,csa_tree_add_51_79_groupi_n_1450);
  and csa_tree_add_51_79_groupi_g42731(csa_tree_add_51_79_groupi_n_3735 ,csa_tree_add_51_79_groupi_n_1880 ,csa_tree_add_51_79_groupi_n_670);
  and csa_tree_add_51_79_groupi_g42732(csa_tree_add_51_79_groupi_n_3734 ,csa_tree_add_51_79_groupi_n_1922 ,csa_tree_add_51_79_groupi_n_2537);
  or csa_tree_add_51_79_groupi_g42733(csa_tree_add_51_79_groupi_n_3732 ,csa_tree_add_51_79_groupi_n_2321 ,csa_tree_add_51_79_groupi_n_1286);
  or csa_tree_add_51_79_groupi_g42734(csa_tree_add_51_79_groupi_n_3731 ,csa_tree_add_51_79_groupi_n_1802 ,csa_tree_add_51_79_groupi_n_1232);
  or csa_tree_add_51_79_groupi_g42735(csa_tree_add_51_79_groupi_n_3730 ,csa_tree_add_51_79_groupi_n_2338 ,csa_tree_add_51_79_groupi_n_1292);
  or csa_tree_add_51_79_groupi_g42736(csa_tree_add_51_79_groupi_n_3729 ,csa_tree_add_51_79_groupi_n_2333 ,csa_tree_add_51_79_groupi_n_1340);
  or csa_tree_add_51_79_groupi_g42737(csa_tree_add_51_79_groupi_n_3728 ,csa_tree_add_51_79_groupi_n_2332 ,csa_tree_add_51_79_groupi_n_1358);
  or csa_tree_add_51_79_groupi_g42738(csa_tree_add_51_79_groupi_n_3727 ,csa_tree_add_51_79_groupi_n_1810 ,csa_tree_add_51_79_groupi_n_2506);
  or csa_tree_add_51_79_groupi_g42739(csa_tree_add_51_79_groupi_n_3726 ,in22[0] ,csa_tree_add_51_79_groupi_n_1539);
  or csa_tree_add_51_79_groupi_g42740(csa_tree_add_51_79_groupi_n_3725 ,in14[0] ,csa_tree_add_51_79_groupi_n_1550);
  or csa_tree_add_51_79_groupi_g42741(csa_tree_add_51_79_groupi_n_3724 ,in24[0] ,csa_tree_add_51_79_groupi_n_1542);
  or csa_tree_add_51_79_groupi_g42742(csa_tree_add_51_79_groupi_n_3723 ,csa_tree_add_51_79_groupi_n_2360 ,csa_tree_add_51_79_groupi_n_1388);
  or csa_tree_add_51_79_groupi_g42743(csa_tree_add_51_79_groupi_n_3722 ,csa_tree_add_51_79_groupi_n_2339 ,csa_tree_add_51_79_groupi_n_1214);
  or csa_tree_add_51_79_groupi_g42744(csa_tree_add_51_79_groupi_n_3721 ,csa_tree_add_51_79_groupi_n_2329 ,csa_tree_add_51_79_groupi_n_1334);
  or csa_tree_add_51_79_groupi_g42745(csa_tree_add_51_79_groupi_n_3720 ,in12[0] ,csa_tree_add_51_79_groupi_n_1540);
  or csa_tree_add_51_79_groupi_g42746(csa_tree_add_51_79_groupi_n_3719 ,csa_tree_add_51_79_groupi_n_2365 ,csa_tree_add_51_79_groupi_n_1271);
  or csa_tree_add_51_79_groupi_g42747(csa_tree_add_51_79_groupi_n_3718 ,csa_tree_add_51_79_groupi_n_1853 ,csa_tree_add_51_79_groupi_n_1274);
  or csa_tree_add_51_79_groupi_g42748(csa_tree_add_51_79_groupi_n_3717 ,csa_tree_add_51_79_groupi_n_1921 ,csa_tree_add_51_79_groupi_n_1382);
  or csa_tree_add_51_79_groupi_g42749(csa_tree_add_51_79_groupi_n_3716 ,in20[0] ,csa_tree_add_51_79_groupi_n_1599);
  or csa_tree_add_51_79_groupi_g42750(csa_tree_add_51_79_groupi_n_3715 ,csa_tree_add_51_79_groupi_n_1795 ,csa_tree_add_51_79_groupi_n_1367);
  or csa_tree_add_51_79_groupi_g42751(csa_tree_add_51_79_groupi_n_3714 ,csa_tree_add_51_79_groupi_n_2347 ,csa_tree_add_51_79_groupi_n_1364);
  or csa_tree_add_51_79_groupi_g42752(csa_tree_add_51_79_groupi_n_3713 ,csa_tree_add_51_79_groupi_n_1801 ,csa_tree_add_51_79_groupi_n_1415);
  or csa_tree_add_51_79_groupi_g42753(csa_tree_add_51_79_groupi_n_3712 ,csa_tree_add_51_79_groupi_n_2354 ,csa_tree_add_51_79_groupi_n_1352);
  or csa_tree_add_51_79_groupi_g42754(csa_tree_add_51_79_groupi_n_3711 ,csa_tree_add_51_79_groupi_n_2403 ,csa_tree_add_51_79_groupi_n_1391);
  or csa_tree_add_51_79_groupi_g42755(csa_tree_add_51_79_groupi_n_3710 ,csa_tree_add_51_79_groupi_n_1791 ,csa_tree_add_51_79_groupi_n_1304);
  or csa_tree_add_51_79_groupi_g42756(csa_tree_add_51_79_groupi_n_3709 ,csa_tree_add_51_79_groupi_n_1796 ,csa_tree_add_51_79_groupi_n_1217);
  or csa_tree_add_51_79_groupi_g42757(csa_tree_add_51_79_groupi_n_3708 ,in4[0] ,csa_tree_add_51_79_groupi_n_1606);
  or csa_tree_add_51_79_groupi_g42758(csa_tree_add_51_79_groupi_n_3707 ,csa_tree_add_51_79_groupi_n_1789 ,csa_tree_add_51_79_groupi_n_1409);
  or csa_tree_add_51_79_groupi_g42759(csa_tree_add_51_79_groupi_n_3706 ,csa_tree_add_51_79_groupi_n_2323 ,csa_tree_add_51_79_groupi_n_1427);
  or csa_tree_add_51_79_groupi_g42760(csa_tree_add_51_79_groupi_n_3705 ,csa_tree_add_51_79_groupi_n_2331 ,csa_tree_add_51_79_groupi_n_1250);
  not csa_tree_add_51_79_groupi_g42761(csa_tree_add_51_79_groupi_n_3371 ,csa_tree_add_51_79_groupi_n_3370);
  not csa_tree_add_51_79_groupi_g42762(csa_tree_add_51_79_groupi_n_3369 ,csa_tree_add_51_79_groupi_n_3368);
  not csa_tree_add_51_79_groupi_g42763(csa_tree_add_51_79_groupi_n_3367 ,csa_tree_add_51_79_groupi_n_3366);
  not csa_tree_add_51_79_groupi_g42764(csa_tree_add_51_79_groupi_n_3365 ,csa_tree_add_51_79_groupi_n_3364);
  not csa_tree_add_51_79_groupi_g42765(csa_tree_add_51_79_groupi_n_3363 ,csa_tree_add_51_79_groupi_n_3362);
  not csa_tree_add_51_79_groupi_g42766(csa_tree_add_51_79_groupi_n_3361 ,csa_tree_add_51_79_groupi_n_3360);
  not csa_tree_add_51_79_groupi_g42767(csa_tree_add_51_79_groupi_n_3359 ,csa_tree_add_51_79_groupi_n_3358);
  not csa_tree_add_51_79_groupi_g42768(csa_tree_add_51_79_groupi_n_3355 ,csa_tree_add_51_79_groupi_n_3354);
  not csa_tree_add_51_79_groupi_g42769(csa_tree_add_51_79_groupi_n_3353 ,csa_tree_add_51_79_groupi_n_3352);
  not csa_tree_add_51_79_groupi_g42770(csa_tree_add_51_79_groupi_n_3347 ,csa_tree_add_51_79_groupi_n_3346);
  not csa_tree_add_51_79_groupi_g42771(csa_tree_add_51_79_groupi_n_3341 ,csa_tree_add_51_79_groupi_n_3340);
  not csa_tree_add_51_79_groupi_g42772(csa_tree_add_51_79_groupi_n_3336 ,csa_tree_add_51_79_groupi_n_3335);
  not csa_tree_add_51_79_groupi_g42774(csa_tree_add_51_79_groupi_n_3309 ,csa_tree_add_51_79_groupi_n_3308);
  not csa_tree_add_51_79_groupi_g42775(csa_tree_add_51_79_groupi_n_3306 ,csa_tree_add_51_79_groupi_n_3305);
  not csa_tree_add_51_79_groupi_g42776(csa_tree_add_51_79_groupi_n_3304 ,csa_tree_add_51_79_groupi_n_3303);
  not csa_tree_add_51_79_groupi_g42777(csa_tree_add_51_79_groupi_n_3302 ,csa_tree_add_51_79_groupi_n_3301);
  not csa_tree_add_51_79_groupi_g42778(csa_tree_add_51_79_groupi_n_3300 ,csa_tree_add_51_79_groupi_n_3299);
  not csa_tree_add_51_79_groupi_g42779(csa_tree_add_51_79_groupi_n_3296 ,csa_tree_add_51_79_groupi_n_3295);
  not csa_tree_add_51_79_groupi_g42780(csa_tree_add_51_79_groupi_n_3292 ,csa_tree_add_51_79_groupi_n_3291);
  not csa_tree_add_51_79_groupi_g42781(csa_tree_add_51_79_groupi_n_3286 ,csa_tree_add_51_79_groupi_n_3285);
  not csa_tree_add_51_79_groupi_g42782(csa_tree_add_51_79_groupi_n_3284 ,csa_tree_add_51_79_groupi_n_3283);
  not csa_tree_add_51_79_groupi_g42783(csa_tree_add_51_79_groupi_n_3279 ,csa_tree_add_51_79_groupi_n_3278);
  not csa_tree_add_51_79_groupi_g42784(csa_tree_add_51_79_groupi_n_3276 ,csa_tree_add_51_79_groupi_n_3275);
  not csa_tree_add_51_79_groupi_g42786(csa_tree_add_51_79_groupi_n_3272 ,csa_tree_add_51_79_groupi_n_3271);
  not csa_tree_add_51_79_groupi_g42788(csa_tree_add_51_79_groupi_n_3260 ,csa_tree_add_51_79_groupi_n_3259);
  not csa_tree_add_51_79_groupi_g42790(csa_tree_add_51_79_groupi_n_3255 ,csa_tree_add_51_79_groupi_n_3254);
  not csa_tree_add_51_79_groupi_g42791(csa_tree_add_51_79_groupi_n_3252 ,csa_tree_add_51_79_groupi_n_3251);
  not csa_tree_add_51_79_groupi_g42792(csa_tree_add_51_79_groupi_n_3249 ,csa_tree_add_51_79_groupi_n_3248);
  not csa_tree_add_51_79_groupi_g42793(csa_tree_add_51_79_groupi_n_3241 ,csa_tree_add_51_79_groupi_n_3240);
  not csa_tree_add_51_79_groupi_g42795(csa_tree_add_51_79_groupi_n_3238 ,csa_tree_add_51_79_groupi_n_3237);
  not csa_tree_add_51_79_groupi_g42796(csa_tree_add_51_79_groupi_n_3235 ,csa_tree_add_51_79_groupi_n_3234);
  not csa_tree_add_51_79_groupi_g42797(csa_tree_add_51_79_groupi_n_3232 ,csa_tree_add_51_79_groupi_n_3231);
  not csa_tree_add_51_79_groupi_g42798(csa_tree_add_51_79_groupi_n_3229 ,csa_tree_add_51_79_groupi_n_3228);
  not csa_tree_add_51_79_groupi_g42799(csa_tree_add_51_79_groupi_n_3227 ,csa_tree_add_51_79_groupi_n_3226);
  not csa_tree_add_51_79_groupi_g42800(csa_tree_add_51_79_groupi_n_3215 ,csa_tree_add_51_79_groupi_n_3214);
  not csa_tree_add_51_79_groupi_g42801(csa_tree_add_51_79_groupi_n_3213 ,csa_tree_add_51_79_groupi_n_3212);
  not csa_tree_add_51_79_groupi_g42802(csa_tree_add_51_79_groupi_n_3197 ,csa_tree_add_51_79_groupi_n_3196);
  or csa_tree_add_51_79_groupi_g42803(csa_tree_add_51_79_groupi_n_3158 ,csa_tree_add_51_79_groupi_n_2090 ,csa_tree_add_51_79_groupi_n_748);
  nor csa_tree_add_51_79_groupi_g42804(csa_tree_add_51_79_groupi_n_3157 ,csa_tree_add_51_79_groupi_n_1687 ,csa_tree_add_51_79_groupi_n_2412);
  or csa_tree_add_51_79_groupi_g42805(csa_tree_add_51_79_groupi_n_3156 ,csa_tree_add_51_79_groupi_n_2193 ,csa_tree_add_51_79_groupi_n_1110);
  or csa_tree_add_51_79_groupi_g42806(csa_tree_add_51_79_groupi_n_3155 ,csa_tree_add_51_79_groupi_n_2738 ,csa_tree_add_51_79_groupi_n_2510);
  or csa_tree_add_51_79_groupi_g42807(csa_tree_add_51_79_groupi_n_3154 ,csa_tree_add_51_79_groupi_n_2093 ,csa_tree_add_51_79_groupi_n_1246);
  or csa_tree_add_51_79_groupi_g42808(csa_tree_add_51_79_groupi_n_3153 ,csa_tree_add_51_79_groupi_n_2318 ,csa_tree_add_51_79_groupi_n_706);
  or csa_tree_add_51_79_groupi_g42809(csa_tree_add_51_79_groupi_n_3152 ,csa_tree_add_51_79_groupi_n_2855 ,csa_tree_add_51_79_groupi_n_736);
  or csa_tree_add_51_79_groupi_g42810(csa_tree_add_51_79_groupi_n_3151 ,csa_tree_add_51_79_groupi_n_2780 ,csa_tree_add_51_79_groupi_n_724);
  or csa_tree_add_51_79_groupi_g42811(csa_tree_add_51_79_groupi_n_3150 ,csa_tree_add_51_79_groupi_n_2109 ,csa_tree_add_51_79_groupi_n_1097);
  or csa_tree_add_51_79_groupi_g42812(csa_tree_add_51_79_groupi_n_3149 ,csa_tree_add_51_79_groupi_n_2765 ,csa_tree_add_51_79_groupi_n_1399);
  or csa_tree_add_51_79_groupi_g42813(csa_tree_add_51_79_groupi_n_3148 ,csa_tree_add_51_79_groupi_n_2086 ,csa_tree_add_51_79_groupi_n_1357);
  or csa_tree_add_51_79_groupi_g42814(csa_tree_add_51_79_groupi_n_3147 ,csa_tree_add_51_79_groupi_n_2652 ,csa_tree_add_51_79_groupi_n_1270);
  or csa_tree_add_51_79_groupi_g42815(csa_tree_add_51_79_groupi_n_3146 ,csa_tree_add_51_79_groupi_n_2626 ,csa_tree_add_51_79_groupi_n_1309);
  or csa_tree_add_51_79_groupi_g42816(csa_tree_add_51_79_groupi_n_3145 ,csa_tree_add_51_79_groupi_n_2754 ,csa_tree_add_51_79_groupi_n_1423);
  or csa_tree_add_51_79_groupi_g42817(csa_tree_add_51_79_groupi_n_3144 ,csa_tree_add_51_79_groupi_n_2135 ,csa_tree_add_51_79_groupi_n_1261);
  or csa_tree_add_51_79_groupi_g42818(csa_tree_add_51_79_groupi_n_3143 ,csa_tree_add_51_79_groupi_n_2800 ,csa_tree_add_51_79_groupi_n_1402);
  nor csa_tree_add_51_79_groupi_g42819(csa_tree_add_51_79_groupi_n_3142 ,csa_tree_add_51_79_groupi_n_1752 ,csa_tree_add_51_79_groupi_n_2373);
  or csa_tree_add_51_79_groupi_g42820(csa_tree_add_51_79_groupi_n_3141 ,csa_tree_add_51_79_groupi_n_2637 ,csa_tree_add_51_79_groupi_n_1330);
  or csa_tree_add_51_79_groupi_g42821(csa_tree_add_51_79_groupi_n_3140 ,csa_tree_add_51_79_groupi_n_2862 ,csa_tree_add_51_79_groupi_n_1339);
  or csa_tree_add_51_79_groupi_g42822(csa_tree_add_51_79_groupi_n_3139 ,csa_tree_add_51_79_groupi_n_2724 ,csa_tree_add_51_79_groupi_n_1105);
  or csa_tree_add_51_79_groupi_g42823(csa_tree_add_51_79_groupi_n_3138 ,csa_tree_add_51_79_groupi_n_2620 ,csa_tree_add_51_79_groupi_n_1225);
  or csa_tree_add_51_79_groupi_g42824(csa_tree_add_51_79_groupi_n_3137 ,csa_tree_add_51_79_groupi_n_2206 ,csa_tree_add_51_79_groupi_n_676);
  or csa_tree_add_51_79_groupi_g42825(csa_tree_add_51_79_groupi_n_3136 ,csa_tree_add_51_79_groupi_n_2867 ,csa_tree_add_51_79_groupi_n_682);
  or csa_tree_add_51_79_groupi_g42826(csa_tree_add_51_79_groupi_n_3135 ,csa_tree_add_51_79_groupi_n_2145 ,csa_tree_add_51_79_groupi_n_2463);
  or csa_tree_add_51_79_groupi_g42827(csa_tree_add_51_79_groupi_n_3134 ,csa_tree_add_51_79_groupi_n_2050 ,csa_tree_add_51_79_groupi_n_1306);
  or csa_tree_add_51_79_groupi_g42828(csa_tree_add_51_79_groupi_n_3133 ,csa_tree_add_51_79_groupi_n_2648 ,csa_tree_add_51_79_groupi_n_1432);
  or csa_tree_add_51_79_groupi_g42829(csa_tree_add_51_79_groupi_n_3132 ,csa_tree_add_51_79_groupi_n_2210 ,csa_tree_add_51_79_groupi_n_697);
  or csa_tree_add_51_79_groupi_g42830(csa_tree_add_51_79_groupi_n_3131 ,csa_tree_add_51_79_groupi_n_2317 ,csa_tree_add_51_79_groupi_n_1411);
  nor csa_tree_add_51_79_groupi_g42831(csa_tree_add_51_79_groupi_n_3130 ,csa_tree_add_51_79_groupi_n_1701 ,csa_tree_add_51_79_groupi_n_2395);
  or csa_tree_add_51_79_groupi_g42832(csa_tree_add_51_79_groupi_n_3129 ,csa_tree_add_51_79_groupi_n_2303 ,csa_tree_add_51_79_groupi_n_1375);
  or csa_tree_add_51_79_groupi_g42833(csa_tree_add_51_79_groupi_n_3128 ,csa_tree_add_51_79_groupi_n_2843 ,csa_tree_add_51_79_groupi_n_1336);
  or csa_tree_add_51_79_groupi_g42834(csa_tree_add_51_79_groupi_n_3127 ,csa_tree_add_51_79_groupi_n_2131 ,csa_tree_add_51_79_groupi_n_1093);
  or csa_tree_add_51_79_groupi_g42835(csa_tree_add_51_79_groupi_n_3126 ,csa_tree_add_51_79_groupi_n_2252 ,csa_tree_add_51_79_groupi_n_1366);
  or csa_tree_add_51_79_groupi_g42836(csa_tree_add_51_79_groupi_n_3125 ,csa_tree_add_51_79_groupi_n_2665 ,csa_tree_add_51_79_groupi_n_1276);
  or csa_tree_add_51_79_groupi_g42837(csa_tree_add_51_79_groupi_n_3124 ,csa_tree_add_51_79_groupi_n_2669 ,csa_tree_add_51_79_groupi_n_1393);
  or csa_tree_add_51_79_groupi_g42838(csa_tree_add_51_79_groupi_n_3123 ,csa_tree_add_51_79_groupi_n_2791 ,csa_tree_add_51_79_groupi_n_1086);
  or csa_tree_add_51_79_groupi_g42839(csa_tree_add_51_79_groupi_n_3122 ,csa_tree_add_51_79_groupi_n_2249 ,csa_tree_add_51_79_groupi_n_1267);
  or csa_tree_add_51_79_groupi_g42840(csa_tree_add_51_79_groupi_n_3121 ,csa_tree_add_51_79_groupi_n_2189 ,csa_tree_add_51_79_groupi_n_1303);
  or csa_tree_add_51_79_groupi_g42841(csa_tree_add_51_79_groupi_n_3120 ,csa_tree_add_51_79_groupi_n_2238 ,csa_tree_add_51_79_groupi_n_2005);
  or csa_tree_add_51_79_groupi_g42842(csa_tree_add_51_79_groupi_n_3119 ,csa_tree_add_51_79_groupi_n_2581 ,csa_tree_add_51_79_groupi_n_745);
  or csa_tree_add_51_79_groupi_g42843(csa_tree_add_51_79_groupi_n_3118 ,csa_tree_add_51_79_groupi_n_2276 ,csa_tree_add_51_79_groupi_n_1112);
  or csa_tree_add_51_79_groupi_g42844(csa_tree_add_51_79_groupi_n_3117 ,csa_tree_add_51_79_groupi_n_2116 ,csa_tree_add_51_79_groupi_n_685);
  or csa_tree_add_51_79_groupi_g42845(csa_tree_add_51_79_groupi_n_3116 ,csa_tree_add_51_79_groupi_n_2020 ,csa_tree_add_51_79_groupi_n_1315);
  or csa_tree_add_51_79_groupi_g42846(csa_tree_add_51_79_groupi_n_3115 ,csa_tree_add_51_79_groupi_n_2144 ,csa_tree_add_51_79_groupi_n_709);
  or csa_tree_add_51_79_groupi_g42847(csa_tree_add_51_79_groupi_n_3114 ,csa_tree_add_51_79_groupi_n_2030 ,csa_tree_add_51_79_groupi_n_1213);
  or csa_tree_add_51_79_groupi_g42848(csa_tree_add_51_79_groupi_n_3113 ,csa_tree_add_51_79_groupi_n_2846 ,csa_tree_add_51_79_groupi_n_1222);
  or csa_tree_add_51_79_groupi_g42849(csa_tree_add_51_79_groupi_n_3112 ,csa_tree_add_51_79_groupi_n_2722 ,csa_tree_add_51_79_groupi_n_1225);
  or csa_tree_add_51_79_groupi_g42850(csa_tree_add_51_79_groupi_n_3111 ,csa_tree_add_51_79_groupi_n_2208 ,csa_tree_add_51_79_groupi_n_1285);
  nor csa_tree_add_51_79_groupi_g42851(csa_tree_add_51_79_groupi_n_3110 ,csa_tree_add_51_79_groupi_n_1727 ,csa_tree_add_51_79_groupi_n_2379);
  or csa_tree_add_51_79_groupi_g42852(csa_tree_add_51_79_groupi_n_3109 ,csa_tree_add_51_79_groupi_n_2250 ,csa_tree_add_51_79_groupi_n_712);
  or csa_tree_add_51_79_groupi_g42853(csa_tree_add_51_79_groupi_n_3108 ,csa_tree_add_51_79_groupi_n_2764 ,csa_tree_add_51_79_groupi_n_1114);
  or csa_tree_add_51_79_groupi_g42854(csa_tree_add_51_79_groupi_n_3107 ,csa_tree_add_51_79_groupi_n_2723 ,csa_tree_add_51_79_groupi_n_2452);
  or csa_tree_add_51_79_groupi_g42855(csa_tree_add_51_79_groupi_n_3106 ,csa_tree_add_51_79_groupi_n_2265 ,csa_tree_add_51_79_groupi_n_2444);
  or csa_tree_add_51_79_groupi_g42856(csa_tree_add_51_79_groupi_n_3105 ,csa_tree_add_51_79_groupi_n_2188 ,csa_tree_add_51_79_groupi_n_694);
  or csa_tree_add_51_79_groupi_g42857(csa_tree_add_51_79_groupi_n_3104 ,csa_tree_add_51_79_groupi_n_2057 ,csa_tree_add_51_79_groupi_n_1408);
  or csa_tree_add_51_79_groupi_g42858(csa_tree_add_51_79_groupi_n_3103 ,csa_tree_add_51_79_groupi_n_2066 ,csa_tree_add_51_79_groupi_n_745);
  or csa_tree_add_51_79_groupi_g42859(csa_tree_add_51_79_groupi_n_3102 ,csa_tree_add_51_79_groupi_n_2299 ,csa_tree_add_51_79_groupi_n_1237);
  or csa_tree_add_51_79_groupi_g42860(csa_tree_add_51_79_groupi_n_3101 ,csa_tree_add_51_79_groupi_n_2186 ,csa_tree_add_51_79_groupi_n_1234);
  or csa_tree_add_51_79_groupi_g42861(csa_tree_add_51_79_groupi_n_3100 ,csa_tree_add_51_79_groupi_n_2232 ,csa_tree_add_51_79_groupi_n_1300);
  or csa_tree_add_51_79_groupi_g42862(csa_tree_add_51_79_groupi_n_3099 ,csa_tree_add_51_79_groupi_n_2673 ,csa_tree_add_51_79_groupi_n_1264);
  or csa_tree_add_51_79_groupi_g42863(csa_tree_add_51_79_groupi_n_3098 ,csa_tree_add_51_79_groupi_n_2096 ,csa_tree_add_51_79_groupi_n_1237);
  or csa_tree_add_51_79_groupi_g42864(csa_tree_add_51_79_groupi_n_3097 ,csa_tree_add_51_79_groupi_n_2268 ,csa_tree_add_51_79_groupi_n_658);
  or csa_tree_add_51_79_groupi_g42865(csa_tree_add_51_79_groupi_n_3096 ,csa_tree_add_51_79_groupi_n_2040 ,csa_tree_add_51_79_groupi_n_1390);
  or csa_tree_add_51_79_groupi_g42866(csa_tree_add_51_79_groupi_n_3095 ,csa_tree_add_51_79_groupi_n_2043 ,csa_tree_add_51_79_groupi_n_706);
  or csa_tree_add_51_79_groupi_g42867(csa_tree_add_51_79_groupi_n_3094 ,csa_tree_add_51_79_groupi_n_2078 ,csa_tree_add_51_79_groupi_n_1115);
  or csa_tree_add_51_79_groupi_g42868(csa_tree_add_51_79_groupi_n_3093 ,csa_tree_add_51_79_groupi_n_2668 ,csa_tree_add_51_79_groupi_n_1360);
  or csa_tree_add_51_79_groupi_g42869(csa_tree_add_51_79_groupi_n_3092 ,csa_tree_add_51_79_groupi_n_2156 ,csa_tree_add_51_79_groupi_n_694);
  or csa_tree_add_51_79_groupi_g42870(csa_tree_add_51_79_groupi_n_3091 ,csa_tree_add_51_79_groupi_n_2573 ,csa_tree_add_51_79_groupi_n_1240);
  or csa_tree_add_51_79_groupi_g42871(csa_tree_add_51_79_groupi_n_3090 ,csa_tree_add_51_79_groupi_n_2756 ,csa_tree_add_51_79_groupi_n_1222);
  or csa_tree_add_51_79_groupi_g42872(csa_tree_add_51_79_groupi_n_3089 ,csa_tree_add_51_79_groupi_n_2622 ,csa_tree_add_51_79_groupi_n_1378);
  nor csa_tree_add_51_79_groupi_g42873(csa_tree_add_51_79_groupi_n_3088 ,csa_tree_add_51_79_groupi_n_1717 ,csa_tree_add_51_79_groupi_n_2386);
  or csa_tree_add_51_79_groupi_g42874(csa_tree_add_51_79_groupi_n_3087 ,csa_tree_add_51_79_groupi_n_2624 ,csa_tree_add_51_79_groupi_n_685);
  or csa_tree_add_51_79_groupi_g42875(csa_tree_add_51_79_groupi_n_3086 ,csa_tree_add_51_79_groupi_n_2736 ,csa_tree_add_51_79_groupi_n_1420);
  or csa_tree_add_51_79_groupi_g42876(csa_tree_add_51_79_groupi_n_3085 ,csa_tree_add_51_79_groupi_n_2837 ,csa_tree_add_51_79_groupi_n_1252);
  or csa_tree_add_51_79_groupi_g42877(csa_tree_add_51_79_groupi_n_3084 ,csa_tree_add_51_79_groupi_n_2835 ,csa_tree_add_51_79_groupi_n_1291);
  or csa_tree_add_51_79_groupi_g42878(csa_tree_add_51_79_groupi_n_3083 ,csa_tree_add_51_79_groupi_n_2583 ,csa_tree_add_51_79_groupi_n_1312);
  or csa_tree_add_51_79_groupi_g42879(csa_tree_add_51_79_groupi_n_3082 ,csa_tree_add_51_79_groupi_n_2854 ,csa_tree_add_51_79_groupi_n_1288);
  or csa_tree_add_51_79_groupi_g42880(csa_tree_add_51_79_groupi_n_3081 ,csa_tree_add_51_79_groupi_n_2149 ,csa_tree_add_51_79_groupi_n_1321);
  or csa_tree_add_51_79_groupi_g42881(csa_tree_add_51_79_groupi_n_3080 ,csa_tree_add_51_79_groupi_n_2301 ,csa_tree_add_51_79_groupi_n_1264);
  or csa_tree_add_51_79_groupi_g42882(csa_tree_add_51_79_groupi_n_3079 ,csa_tree_add_51_79_groupi_n_2079 ,csa_tree_add_51_79_groupi_n_739);
  or csa_tree_add_51_79_groupi_g42883(csa_tree_add_51_79_groupi_n_3078 ,csa_tree_add_51_79_groupi_n_2233 ,csa_tree_add_51_79_groupi_n_673);
  or csa_tree_add_51_79_groupi_g42884(csa_tree_add_51_79_groupi_n_3077 ,csa_tree_add_51_79_groupi_n_2128 ,csa_tree_add_51_79_groupi_n_1426);
  or csa_tree_add_51_79_groupi_g42885(csa_tree_add_51_79_groupi_n_3076 ,csa_tree_add_51_79_groupi_n_2715 ,csa_tree_add_51_79_groupi_n_1354);
  or csa_tree_add_51_79_groupi_g42886(csa_tree_add_51_79_groupi_n_3075 ,csa_tree_add_51_79_groupi_n_2056 ,csa_tree_add_51_79_groupi_n_1291);
  nor csa_tree_add_51_79_groupi_g42887(csa_tree_add_51_79_groupi_n_3074 ,csa_tree_add_51_79_groupi_n_1767 ,csa_tree_add_51_79_groupi_n_2374);
  or csa_tree_add_51_79_groupi_g42888(csa_tree_add_51_79_groupi_n_3073 ,csa_tree_add_51_79_groupi_n_2719 ,csa_tree_add_51_79_groupi_n_1240);
  or csa_tree_add_51_79_groupi_g42889(csa_tree_add_51_79_groupi_n_3072 ,csa_tree_add_51_79_groupi_n_2260 ,csa_tree_add_51_79_groupi_n_1106);
  or csa_tree_add_51_79_groupi_g42890(csa_tree_add_51_79_groupi_n_3071 ,csa_tree_add_51_79_groupi_n_2633 ,csa_tree_add_51_79_groupi_n_1351);
  nor csa_tree_add_51_79_groupi_g42891(csa_tree_add_51_79_groupi_n_3070 ,csa_tree_add_51_79_groupi_n_1750 ,csa_tree_add_51_79_groupi_n_2385);
  nor csa_tree_add_51_79_groupi_g42892(csa_tree_add_51_79_groupi_n_3069 ,csa_tree_add_51_79_groupi_n_1676 ,csa_tree_add_51_79_groupi_n_2407);
  or csa_tree_add_51_79_groupi_g42893(csa_tree_add_51_79_groupi_n_3068 ,csa_tree_add_51_79_groupi_n_2775 ,csa_tree_add_51_79_groupi_n_1096);
  nor csa_tree_add_51_79_groupi_g42894(csa_tree_add_51_79_groupi_n_3067 ,csa_tree_add_51_79_groupi_n_1705 ,csa_tree_add_51_79_groupi_n_2402);
  nor csa_tree_add_51_79_groupi_g42895(csa_tree_add_51_79_groupi_n_3066 ,csa_tree_add_51_79_groupi_n_1730 ,csa_tree_add_51_79_groupi_n_2432);
  or csa_tree_add_51_79_groupi_g42896(csa_tree_add_51_79_groupi_n_3065 ,csa_tree_add_51_79_groupi_n_2789 ,csa_tree_add_51_79_groupi_n_1315);
  or csa_tree_add_51_79_groupi_g42897(csa_tree_add_51_79_groupi_n_3064 ,csa_tree_add_51_79_groupi_n_2834 ,csa_tree_add_51_79_groupi_n_2486);
  or csa_tree_add_51_79_groupi_g42898(csa_tree_add_51_79_groupi_n_3063 ,csa_tree_add_51_79_groupi_n_2817 ,csa_tree_add_51_79_groupi_n_1094);
  nor csa_tree_add_51_79_groupi_g42899(csa_tree_add_51_79_groupi_n_3062 ,csa_tree_add_51_79_groupi_n_1710 ,csa_tree_add_51_79_groupi_n_2388);
  or csa_tree_add_51_79_groupi_g42900(csa_tree_add_51_79_groupi_n_3061 ,csa_tree_add_51_79_groupi_n_2036 ,csa_tree_add_51_79_groupi_n_1387);
  or csa_tree_add_51_79_groupi_g42901(csa_tree_add_51_79_groupi_n_3060 ,csa_tree_add_51_79_groupi_n_2579 ,csa_tree_add_51_79_groupi_n_1104);
  or csa_tree_add_51_79_groupi_g42902(csa_tree_add_51_79_groupi_n_3059 ,csa_tree_add_51_79_groupi_n_2658 ,csa_tree_add_51_79_groupi_n_1246);
  or csa_tree_add_51_79_groupi_g42903(csa_tree_add_51_79_groupi_n_3058 ,csa_tree_add_51_79_groupi_n_2226 ,csa_tree_add_51_79_groupi_n_748);
  nor csa_tree_add_51_79_groupi_g42904(csa_tree_add_51_79_groupi_n_3057 ,csa_tree_add_51_79_groupi_n_1691 ,csa_tree_add_51_79_groupi_n_2423);
  or csa_tree_add_51_79_groupi_g42905(csa_tree_add_51_79_groupi_n_3056 ,csa_tree_add_51_79_groupi_n_2085 ,csa_tree_add_51_79_groupi_n_1089);
  or csa_tree_add_51_79_groupi_g42906(csa_tree_add_51_79_groupi_n_3055 ,csa_tree_add_51_79_groupi_n_2650 ,csa_tree_add_51_79_groupi_n_1246);
  or csa_tree_add_51_79_groupi_g42907(csa_tree_add_51_79_groupi_n_3054 ,csa_tree_add_51_79_groupi_n_2115 ,csa_tree_add_51_79_groupi_n_1297);
  nor csa_tree_add_51_79_groupi_g42908(csa_tree_add_51_79_groupi_n_3053 ,csa_tree_add_51_79_groupi_n_1725 ,csa_tree_add_51_79_groupi_n_2411);
  or csa_tree_add_51_79_groupi_g42909(csa_tree_add_51_79_groupi_n_3052 ,csa_tree_add_51_79_groupi_n_2826 ,csa_tree_add_51_79_groupi_n_1381);
  or csa_tree_add_51_79_groupi_g42910(csa_tree_add_51_79_groupi_n_3051 ,csa_tree_add_51_79_groupi_n_2304 ,csa_tree_add_51_79_groupi_n_730);
  or csa_tree_add_51_79_groupi_g42911(csa_tree_add_51_79_groupi_n_3050 ,csa_tree_add_51_79_groupi_n_2295 ,csa_tree_add_51_79_groupi_n_1091);
  nor csa_tree_add_51_79_groupi_g42912(csa_tree_add_51_79_groupi_n_3049 ,csa_tree_add_51_79_groupi_n_1683 ,csa_tree_add_51_79_groupi_n_2387);
  or csa_tree_add_51_79_groupi_g42913(csa_tree_add_51_79_groupi_n_3048 ,csa_tree_add_51_79_groupi_n_2122 ,csa_tree_add_51_79_groupi_n_1234);
  or csa_tree_add_51_79_groupi_g42914(csa_tree_add_51_79_groupi_n_3047 ,csa_tree_add_51_79_groupi_n_2044 ,csa_tree_add_51_79_groupi_n_2460);
  nor csa_tree_add_51_79_groupi_g42915(csa_tree_add_51_79_groupi_n_3046 ,csa_tree_add_51_79_groupi_n_1735 ,csa_tree_add_51_79_groupi_n_2391);
  nor csa_tree_add_51_79_groupi_g42916(csa_tree_add_51_79_groupi_n_3045 ,csa_tree_add_51_79_groupi_n_1719 ,csa_tree_add_51_79_groupi_n_2427);
  or csa_tree_add_51_79_groupi_g42917(csa_tree_add_51_79_groupi_n_3044 ,csa_tree_add_51_79_groupi_n_2731 ,csa_tree_add_51_79_groupi_n_682);
  or csa_tree_add_51_79_groupi_g42918(csa_tree_add_51_79_groupi_n_3043 ,csa_tree_add_51_79_groupi_n_2049 ,csa_tree_add_51_79_groupi_n_2491);
  nor csa_tree_add_51_79_groupi_g42919(csa_tree_add_51_79_groupi_n_3042 ,csa_tree_add_51_79_groupi_n_1746 ,csa_tree_add_51_79_groupi_n_2410);
  or csa_tree_add_51_79_groupi_g42920(csa_tree_add_51_79_groupi_n_3041 ,csa_tree_add_51_79_groupi_n_2684 ,csa_tree_add_51_79_groupi_n_1228);
  or csa_tree_add_51_79_groupi_g42921(csa_tree_add_51_79_groupi_n_3040 ,csa_tree_add_51_79_groupi_n_2235 ,csa_tree_add_51_79_groupi_n_730);
  nor csa_tree_add_51_79_groupi_g42922(csa_tree_add_51_79_groupi_n_3039 ,csa_tree_add_51_79_groupi_n_1715 ,csa_tree_add_51_79_groupi_n_2396);
  or csa_tree_add_51_79_groupi_g42923(csa_tree_add_51_79_groupi_n_3038 ,csa_tree_add_51_79_groupi_n_2222 ,csa_tree_add_51_79_groupi_n_1249);
  or csa_tree_add_51_79_groupi_g42924(csa_tree_add_51_79_groupi_n_3037 ,csa_tree_add_51_79_groupi_n_2642 ,csa_tree_add_51_79_groupi_n_706);
  nor csa_tree_add_51_79_groupi_g42925(csa_tree_add_51_79_groupi_n_3036 ,csa_tree_add_51_79_groupi_n_1731 ,csa_tree_add_51_79_groupi_n_2398);
  or csa_tree_add_51_79_groupi_g42926(csa_tree_add_51_79_groupi_n_3035 ,csa_tree_add_51_79_groupi_n_2021 ,csa_tree_add_51_79_groupi_n_1375);
  or csa_tree_add_51_79_groupi_g42927(csa_tree_add_51_79_groupi_n_3034 ,csa_tree_add_51_79_groupi_n_2292 ,csa_tree_add_51_79_groupi_n_1429);
  or csa_tree_add_51_79_groupi_g42928(csa_tree_add_51_79_groupi_n_3033 ,csa_tree_add_51_79_groupi_n_2680 ,csa_tree_add_51_79_groupi_n_1255);
  or csa_tree_add_51_79_groupi_g42929(csa_tree_add_51_79_groupi_n_3032 ,csa_tree_add_51_79_groupi_n_2728 ,csa_tree_add_51_79_groupi_n_2002);
  nor csa_tree_add_51_79_groupi_g42930(csa_tree_add_51_79_groupi_n_3031 ,csa_tree_add_51_79_groupi_n_1770 ,csa_tree_add_51_79_groupi_n_2409);
  or csa_tree_add_51_79_groupi_g42931(csa_tree_add_51_79_groupi_n_3030 ,csa_tree_add_51_79_groupi_n_2827 ,csa_tree_add_51_79_groupi_n_736);
  or csa_tree_add_51_79_groupi_g42932(csa_tree_add_51_79_groupi_n_3029 ,csa_tree_add_51_79_groupi_n_2786 ,csa_tree_add_51_79_groupi_n_1100);
  or csa_tree_add_51_79_groupi_g42933(csa_tree_add_51_79_groupi_n_3028 ,csa_tree_add_51_79_groupi_n_2165 ,csa_tree_add_51_79_groupi_n_697);
  or csa_tree_add_51_79_groupi_g42934(csa_tree_add_51_79_groupi_n_3027 ,csa_tree_add_51_79_groupi_n_2749 ,csa_tree_add_51_79_groupi_n_1294);
  or csa_tree_add_51_79_groupi_g42935(csa_tree_add_51_79_groupi_n_3026 ,csa_tree_add_51_79_groupi_n_2662 ,csa_tree_add_51_79_groupi_n_1333);
  or csa_tree_add_51_79_groupi_g42936(csa_tree_add_51_79_groupi_n_3025 ,csa_tree_add_51_79_groupi_n_2678 ,csa_tree_add_51_79_groupi_n_1348);
  or csa_tree_add_51_79_groupi_g42937(csa_tree_add_51_79_groupi_n_3024 ,csa_tree_add_51_79_groupi_n_2868 ,csa_tree_add_51_79_groupi_n_1107);
  or csa_tree_add_51_79_groupi_g42938(csa_tree_add_51_79_groupi_n_3023 ,csa_tree_add_51_79_groupi_n_2599 ,csa_tree_add_51_79_groupi_n_1279);
  or csa_tree_add_51_79_groupi_g42939(csa_tree_add_51_79_groupi_n_3022 ,csa_tree_add_51_79_groupi_n_2203 ,csa_tree_add_51_79_groupi_n_709);
  or csa_tree_add_51_79_groupi_g42940(csa_tree_add_51_79_groupi_n_3021 ,csa_tree_add_51_79_groupi_n_2302 ,csa_tree_add_51_79_groupi_n_1312);
  or csa_tree_add_51_79_groupi_g42941(csa_tree_add_51_79_groupi_n_3020 ,csa_tree_add_51_79_groupi_n_2709 ,csa_tree_add_51_79_groupi_n_748);
  or csa_tree_add_51_79_groupi_g42942(csa_tree_add_51_79_groupi_n_3019 ,csa_tree_add_51_79_groupi_n_2763 ,csa_tree_add_51_79_groupi_n_1108);
  or csa_tree_add_51_79_groupi_g42943(csa_tree_add_51_79_groupi_n_3018 ,csa_tree_add_51_79_groupi_n_2592 ,csa_tree_add_51_79_groupi_n_1405);
  or csa_tree_add_51_79_groupi_g42944(csa_tree_add_51_79_groupi_n_3017 ,csa_tree_add_51_79_groupi_n_2842 ,csa_tree_add_51_79_groupi_n_1276);
  or csa_tree_add_51_79_groupi_g42945(csa_tree_add_51_79_groupi_n_3016 ,csa_tree_add_51_79_groupi_n_2150 ,csa_tree_add_51_79_groupi_n_1288);
  or csa_tree_add_51_79_groupi_g42946(csa_tree_add_51_79_groupi_n_3015 ,csa_tree_add_51_79_groupi_n_2179 ,csa_tree_add_51_79_groupi_n_1282);
  or csa_tree_add_51_79_groupi_g42947(csa_tree_add_51_79_groupi_n_3014 ,csa_tree_add_51_79_groupi_n_2542 ,csa_tree_add_51_79_groupi_n_2546);
  or csa_tree_add_51_79_groupi_g42948(csa_tree_add_51_79_groupi_n_3013 ,csa_tree_add_51_79_groupi_n_2816 ,csa_tree_add_51_79_groupi_n_724);
  or csa_tree_add_51_79_groupi_g42949(csa_tree_add_51_79_groupi_n_3012 ,csa_tree_add_51_79_groupi_n_2647 ,csa_tree_add_51_79_groupi_n_2494);
  or csa_tree_add_51_79_groupi_g42950(csa_tree_add_51_79_groupi_n_3011 ,csa_tree_add_51_79_groupi_n_2068 ,csa_tree_add_51_79_groupi_n_2483);
  or csa_tree_add_51_79_groupi_g42951(csa_tree_add_51_79_groupi_n_3010 ,csa_tree_add_51_79_groupi_n_2819 ,csa_tree_add_51_79_groupi_n_706);
  or csa_tree_add_51_79_groupi_g42952(csa_tree_add_51_79_groupi_n_3009 ,csa_tree_add_51_79_groupi_n_2225 ,csa_tree_add_51_79_groupi_n_709);
  or csa_tree_add_51_79_groupi_g42953(csa_tree_add_51_79_groupi_n_3008 ,csa_tree_add_51_79_groupi_n_2557 ,csa_tree_add_51_79_groupi_n_2556);
  and csa_tree_add_51_79_groupi_g42954(csa_tree_add_51_79_groupi_n_3007 ,csa_tree_add_51_79_groupi_n_2557 ,csa_tree_add_51_79_groupi_n_2556);
  or csa_tree_add_51_79_groupi_g42955(csa_tree_add_51_79_groupi_n_3006 ,csa_tree_add_51_79_groupi_n_2311 ,csa_tree_add_51_79_groupi_n_682);
  or csa_tree_add_51_79_groupi_g42956(csa_tree_add_51_79_groupi_n_3005 ,csa_tree_add_51_79_groupi_n_2801 ,csa_tree_add_51_79_groupi_n_1976);
  or csa_tree_add_51_79_groupi_g42957(csa_tree_add_51_79_groupi_n_3004 ,csa_tree_add_51_79_groupi_n_2878 ,csa_tree_add_51_79_groupi_n_1088);
  nor csa_tree_add_51_79_groupi_g42958(csa_tree_add_51_79_groupi_n_3003 ,csa_tree_add_51_79_groupi_n_2544 ,csa_tree_add_51_79_groupi_n_2547);
  or csa_tree_add_51_79_groupi_g42959(csa_tree_add_51_79_groupi_n_3002 ,csa_tree_add_51_79_groupi_n_2274 ,csa_tree_add_51_79_groupi_n_1113);
  or csa_tree_add_51_79_groupi_g42960(csa_tree_add_51_79_groupi_n_3001 ,csa_tree_add_51_79_groupi_n_2787 ,csa_tree_add_51_79_groupi_n_1255);
  or csa_tree_add_51_79_groupi_g42961(csa_tree_add_51_79_groupi_n_3000 ,csa_tree_add_51_79_groupi_n_2123 ,csa_tree_add_51_79_groupi_n_2014);
  or csa_tree_add_51_79_groupi_g42962(csa_tree_add_51_79_groupi_n_2999 ,csa_tree_add_51_79_groupi_n_2829 ,csa_tree_add_51_79_groupi_n_1444);
  or csa_tree_add_51_79_groupi_g42963(csa_tree_add_51_79_groupi_n_2998 ,csa_tree_add_51_79_groupi_n_2850 ,csa_tree_add_51_79_groupi_n_1384);
  or csa_tree_add_51_79_groupi_g42964(csa_tree_add_51_79_groupi_n_2997 ,csa_tree_add_51_79_groupi_n_2185 ,csa_tree_add_51_79_groupi_n_1095);
  or csa_tree_add_51_79_groupi_g42965(csa_tree_add_51_79_groupi_n_2996 ,csa_tree_add_51_79_groupi_n_2839 ,csa_tree_add_51_79_groupi_n_685);
  or csa_tree_add_51_79_groupi_g42966(csa_tree_add_51_79_groupi_n_2995 ,csa_tree_add_51_79_groupi_n_2840 ,csa_tree_add_51_79_groupi_n_1228);
  or csa_tree_add_51_79_groupi_g42967(csa_tree_add_51_79_groupi_n_2994 ,csa_tree_add_51_79_groupi_n_2704 ,csa_tree_add_51_79_groupi_n_2438);
  or csa_tree_add_51_79_groupi_g42968(csa_tree_add_51_79_groupi_n_2993 ,csa_tree_add_51_79_groupi_n_2306 ,csa_tree_add_51_79_groupi_n_1345);
  or csa_tree_add_51_79_groupi_g42969(csa_tree_add_51_79_groupi_n_2992 ,csa_tree_add_51_79_groupi_n_2125 ,csa_tree_add_51_79_groupi_n_1303);
  or csa_tree_add_51_79_groupi_g42970(csa_tree_add_51_79_groupi_n_2991 ,csa_tree_add_51_79_groupi_n_2660 ,csa_tree_add_51_79_groupi_n_1102);
  and csa_tree_add_51_79_groupi_g42971(csa_tree_add_51_79_groupi_n_2990 ,csa_tree_add_51_79_groupi_n_2553 ,csa_tree_add_51_79_groupi_n_2554);
  or csa_tree_add_51_79_groupi_g42972(csa_tree_add_51_79_groupi_n_2989 ,csa_tree_add_51_79_groupi_n_2613 ,csa_tree_add_51_79_groupi_n_739);
  or csa_tree_add_51_79_groupi_g42973(csa_tree_add_51_79_groupi_n_2988 ,csa_tree_add_51_79_groupi_n_2070 ,csa_tree_add_51_79_groupi_n_2505);
  or csa_tree_add_51_79_groupi_g42974(csa_tree_add_51_79_groupi_n_2987 ,csa_tree_add_51_79_groupi_n_2124 ,csa_tree_add_51_79_groupi_n_676);
  or csa_tree_add_51_79_groupi_g42975(csa_tree_add_51_79_groupi_n_2986 ,csa_tree_add_51_79_groupi_n_2720 ,csa_tree_add_51_79_groupi_n_1098);
  or csa_tree_add_51_79_groupi_g42976(csa_tree_add_51_79_groupi_n_2985 ,csa_tree_add_51_79_groupi_n_2246 ,csa_tree_add_51_79_groupi_n_2472);
  or csa_tree_add_51_79_groupi_g42977(csa_tree_add_51_79_groupi_n_2984 ,csa_tree_add_51_79_groupi_n_2861 ,csa_tree_add_51_79_groupi_n_745);
  or csa_tree_add_51_79_groupi_g42978(csa_tree_add_51_79_groupi_n_2983 ,csa_tree_add_51_79_groupi_n_2294 ,csa_tree_add_51_79_groupi_n_2441);
  or csa_tree_add_51_79_groupi_g42979(csa_tree_add_51_79_groupi_n_2982 ,csa_tree_add_51_79_groupi_n_2207 ,csa_tree_add_51_79_groupi_n_1300);
  or csa_tree_add_51_79_groupi_g42980(csa_tree_add_51_79_groupi_n_2981 ,csa_tree_add_51_79_groupi_n_2190 ,csa_tree_add_51_79_groupi_n_1417);
  nor csa_tree_add_51_79_groupi_g42981(csa_tree_add_51_79_groupi_n_2980 ,csa_tree_add_51_79_groupi_n_1689 ,csa_tree_add_51_79_groupi_n_2390);
  or csa_tree_add_51_79_groupi_g42982(csa_tree_add_51_79_groupi_n_2979 ,csa_tree_add_51_79_groupi_n_2105 ,csa_tree_add_51_79_groupi_n_724);
  or csa_tree_add_51_79_groupi_g42983(csa_tree_add_51_79_groupi_n_2978 ,csa_tree_add_51_79_groupi_n_2198 ,csa_tree_add_51_79_groupi_n_2500);
  or csa_tree_add_51_79_groupi_g42984(csa_tree_add_51_79_groupi_n_2977 ,csa_tree_add_51_79_groupi_n_2241 ,csa_tree_add_51_79_groupi_n_1372);
  or csa_tree_add_51_79_groupi_g42985(csa_tree_add_51_79_groupi_n_2976 ,csa_tree_add_51_79_groupi_n_2160 ,csa_tree_add_51_79_groupi_n_1261);
  or csa_tree_add_51_79_groupi_g42986(csa_tree_add_51_79_groupi_n_2975 ,csa_tree_add_51_79_groupi_n_2739 ,csa_tree_add_51_79_groupi_n_1087);
  or csa_tree_add_51_79_groupi_g42987(csa_tree_add_51_79_groupi_n_2974 ,csa_tree_add_51_79_groupi_n_2180 ,csa_tree_add_51_79_groupi_n_1234);
  or csa_tree_add_51_79_groupi_g42988(csa_tree_add_51_79_groupi_n_2973 ,csa_tree_add_51_79_groupi_n_2714 ,csa_tree_add_51_79_groupi_n_1213);
  or csa_tree_add_51_79_groupi_g42989(csa_tree_add_51_79_groupi_n_2972 ,csa_tree_add_51_79_groupi_n_2258 ,csa_tree_add_51_79_groupi_n_1369);
  or csa_tree_add_51_79_groupi_g42990(csa_tree_add_51_79_groupi_n_2971 ,csa_tree_add_51_79_groupi_n_2705 ,csa_tree_add_51_79_groupi_n_1435);
  or csa_tree_add_51_79_groupi_g42991(csa_tree_add_51_79_groupi_n_2970 ,csa_tree_add_51_79_groupi_n_2088 ,csa_tree_add_51_79_groupi_n_712);
  or csa_tree_add_51_79_groupi_g42992(csa_tree_add_51_79_groupi_n_2969 ,csa_tree_add_51_79_groupi_n_2161 ,csa_tree_add_51_79_groupi_n_700);
  or csa_tree_add_51_79_groupi_g42993(csa_tree_add_51_79_groupi_n_2968 ,csa_tree_add_51_79_groupi_n_2733 ,csa_tree_add_51_79_groupi_n_1273);
  or csa_tree_add_51_79_groupi_g42994(csa_tree_add_51_79_groupi_n_2967 ,csa_tree_add_51_79_groupi_n_2223 ,csa_tree_add_51_79_groupi_n_739);
  or csa_tree_add_51_79_groupi_g42995(csa_tree_add_51_79_groupi_n_2966 ,csa_tree_add_51_79_groupi_n_2832 ,csa_tree_add_51_79_groupi_n_1414);
  and csa_tree_add_51_79_groupi_g42996(csa_tree_add_51_79_groupi_n_2965 ,csa_tree_add_51_79_groupi_n_2551 ,csa_tree_add_51_79_groupi_n_2549);
  or csa_tree_add_51_79_groupi_g42997(csa_tree_add_51_79_groupi_n_2964 ,csa_tree_add_51_79_groupi_n_2670 ,csa_tree_add_51_79_groupi_n_1109);
  or csa_tree_add_51_79_groupi_g42998(csa_tree_add_51_79_groupi_n_2963 ,csa_tree_add_51_79_groupi_n_2598 ,csa_tree_add_51_79_groupi_n_2475);
  or csa_tree_add_51_79_groupi_g42999(csa_tree_add_51_79_groupi_n_2962 ,csa_tree_add_51_79_groupi_n_2701 ,csa_tree_add_51_79_groupi_n_1973);
  or csa_tree_add_51_79_groupi_g43000(csa_tree_add_51_79_groupi_n_2961 ,csa_tree_add_51_79_groupi_n_2269 ,csa_tree_add_51_79_groupi_n_1099);
  or csa_tree_add_51_79_groupi_g43001(csa_tree_add_51_79_groupi_n_2960 ,csa_tree_add_51_79_groupi_n_2616 ,csa_tree_add_51_79_groupi_n_1309);
  or csa_tree_add_51_79_groupi_g43002(csa_tree_add_51_79_groupi_n_2959 ,csa_tree_add_51_79_groupi_n_2054 ,csa_tree_add_51_79_groupi_n_1342);
  or csa_tree_add_51_79_groupi_g43003(csa_tree_add_51_79_groupi_n_2958 ,csa_tree_add_51_79_groupi_n_2284 ,csa_tree_add_51_79_groupi_n_2449);
  or csa_tree_add_51_79_groupi_g43004(csa_tree_add_51_79_groupi_n_2957 ,csa_tree_add_51_79_groupi_n_2287 ,csa_tree_add_51_79_groupi_n_1315);
  or csa_tree_add_51_79_groupi_g43005(csa_tree_add_51_79_groupi_n_2956 ,csa_tree_add_51_79_groupi_n_2796 ,csa_tree_add_51_79_groupi_n_2469);
  or csa_tree_add_51_79_groupi_g43006(csa_tree_add_51_79_groupi_n_2955 ,csa_tree_add_51_79_groupi_n_2769 ,csa_tree_add_51_79_groupi_n_1216);
  or csa_tree_add_51_79_groupi_g43007(csa_tree_add_51_79_groupi_n_2954 ,csa_tree_add_51_79_groupi_n_2881 ,csa_tree_add_51_79_groupi_n_1423);
  or csa_tree_add_51_79_groupi_g43008(csa_tree_add_51_79_groupi_n_2953 ,csa_tree_add_51_79_groupi_n_2869 ,csa_tree_add_51_79_groupi_n_2008);
  or csa_tree_add_51_79_groupi_g43009(csa_tree_add_51_79_groupi_n_2952 ,csa_tree_add_51_79_groupi_n_2836 ,csa_tree_add_51_79_groupi_n_1438);
  or csa_tree_add_51_79_groupi_g43010(csa_tree_add_51_79_groupi_n_2951 ,csa_tree_add_51_79_groupi_n_2015 ,csa_tree_add_51_79_groupi_n_1097);
  or csa_tree_add_51_79_groupi_g43011(csa_tree_add_51_79_groupi_n_2950 ,csa_tree_add_51_79_groupi_n_2602 ,csa_tree_add_51_79_groupi_n_1399);
  or csa_tree_add_51_79_groupi_g43012(csa_tree_add_51_79_groupi_n_2949 ,csa_tree_add_51_79_groupi_n_2081 ,csa_tree_add_51_79_groupi_n_1363);
  or csa_tree_add_51_79_groupi_g43013(csa_tree_add_51_79_groupi_n_2948 ,csa_tree_add_51_79_groupi_n_2779 ,csa_tree_add_51_79_groupi_n_1429);
  or csa_tree_add_51_79_groupi_g43014(csa_tree_add_51_79_groupi_n_2947 ,csa_tree_add_51_79_groupi_n_2191 ,csa_tree_add_51_79_groupi_n_673);
  or csa_tree_add_51_79_groupi_g43015(csa_tree_add_51_79_groupi_n_2946 ,csa_tree_add_51_79_groupi_n_2215 ,csa_tree_add_51_79_groupi_n_1231);
  or csa_tree_add_51_79_groupi_g43016(csa_tree_add_51_79_groupi_n_2945 ,csa_tree_add_51_79_groupi_n_2605 ,csa_tree_add_51_79_groupi_n_1402);
  or csa_tree_add_51_79_groupi_g43017(csa_tree_add_51_79_groupi_n_2944 ,csa_tree_add_51_79_groupi_n_2694 ,csa_tree_add_51_79_groupi_n_1222);
  or csa_tree_add_51_79_groupi_g43018(csa_tree_add_51_79_groupi_n_2943 ,csa_tree_add_51_79_groupi_n_2828 ,csa_tree_add_51_79_groupi_n_2011);
  or csa_tree_add_51_79_groupi_g43019(csa_tree_add_51_79_groupi_n_2942 ,csa_tree_add_51_79_groupi_n_2634 ,csa_tree_add_51_79_groupi_n_1111);
  or csa_tree_add_51_79_groupi_g43020(csa_tree_add_51_79_groupi_n_2941 ,csa_tree_add_51_79_groupi_n_2809 ,csa_tree_add_51_79_groupi_n_1441);
  or csa_tree_add_51_79_groupi_g43021(csa_tree_add_51_79_groupi_n_2940 ,csa_tree_add_51_79_groupi_n_2712 ,csa_tree_add_51_79_groupi_n_685);
  or csa_tree_add_51_79_groupi_g43022(csa_tree_add_51_79_groupi_n_2939 ,csa_tree_add_51_79_groupi_n_2596 ,csa_tree_add_51_79_groupi_n_1396);
  or csa_tree_add_51_79_groupi_g43023(csa_tree_add_51_79_groupi_n_2938 ,csa_tree_add_51_79_groupi_n_2699 ,csa_tree_add_51_79_groupi_n_1312);
  or csa_tree_add_51_79_groupi_g43024(csa_tree_add_51_79_groupi_n_2937 ,csa_tree_add_51_79_groupi_n_2091 ,csa_tree_add_51_79_groupi_n_1270);
  or csa_tree_add_51_79_groupi_g43025(csa_tree_add_51_79_groupi_n_2936 ,csa_tree_add_51_79_groupi_n_2017 ,csa_tree_add_51_79_groupi_n_1420);
  or csa_tree_add_51_79_groupi_g43026(csa_tree_add_51_79_groupi_n_2935 ,csa_tree_add_51_79_groupi_n_2864 ,csa_tree_add_51_79_groupi_n_1108);
  or csa_tree_add_51_79_groupi_g43027(csa_tree_add_51_79_groupi_n_2934 ,csa_tree_add_51_79_groupi_n_2663 ,csa_tree_add_51_79_groupi_n_1366);
  or csa_tree_add_51_79_groupi_g43028(csa_tree_add_51_79_groupi_n_2933 ,csa_tree_add_51_79_groupi_n_2863 ,csa_tree_add_51_79_groupi_n_1104);
  or csa_tree_add_51_79_groupi_g43029(csa_tree_add_51_79_groupi_n_2932 ,csa_tree_add_51_79_groupi_n_2272 ,csa_tree_add_51_79_groupi_n_1318);
  or csa_tree_add_51_79_groupi_g43030(csa_tree_add_51_79_groupi_n_2931 ,csa_tree_add_51_79_groupi_n_2187 ,csa_tree_add_51_79_groupi_n_1249);
  or csa_tree_add_51_79_groupi_g43031(csa_tree_add_51_79_groupi_n_2930 ,csa_tree_add_51_79_groupi_n_2806 ,csa_tree_add_51_79_groupi_n_1228);
  or csa_tree_add_51_79_groupi_g43032(csa_tree_add_51_79_groupi_n_2929 ,csa_tree_add_51_79_groupi_n_2279 ,csa_tree_add_51_79_groupi_n_1306);
  or csa_tree_add_51_79_groupi_g43033(csa_tree_add_51_79_groupi_n_2928 ,csa_tree_add_51_79_groupi_n_2797 ,csa_tree_add_51_79_groupi_n_1246);
  or csa_tree_add_51_79_groupi_g43034(csa_tree_add_51_79_groupi_n_2927 ,csa_tree_add_51_79_groupi_n_2777 ,csa_tree_add_51_79_groupi_n_1086);
  or csa_tree_add_51_79_groupi_g43035(csa_tree_add_51_79_groupi_n_2926 ,csa_tree_add_51_79_groupi_n_2176 ,csa_tree_add_51_79_groupi_n_700);
  or csa_tree_add_51_79_groupi_g43036(csa_tree_add_51_79_groupi_n_2925 ,csa_tree_add_51_79_groupi_n_2089 ,csa_tree_add_51_79_groupi_n_1330);
  or csa_tree_add_51_79_groupi_g43037(csa_tree_add_51_79_groupi_n_2924 ,csa_tree_add_51_79_groupi_n_2154 ,csa_tree_add_51_79_groupi_n_694);
  or csa_tree_add_51_79_groupi_g43038(csa_tree_add_51_79_groupi_n_2923 ,csa_tree_add_51_79_groupi_n_2687 ,csa_tree_add_51_79_groupi_n_751);
  or csa_tree_add_51_79_groupi_g43039(csa_tree_add_51_79_groupi_n_2922 ,csa_tree_add_51_79_groupi_n_2770 ,csa_tree_add_51_79_groupi_n_1411);
  or csa_tree_add_51_79_groupi_g43040(csa_tree_add_51_79_groupi_n_2921 ,csa_tree_add_51_79_groupi_n_2273 ,csa_tree_add_51_79_groupi_n_694);
  or csa_tree_add_51_79_groupi_g43041(csa_tree_add_51_79_groupi_n_2920 ,csa_tree_add_51_79_groupi_n_2697 ,csa_tree_add_51_79_groupi_n_751);
  or csa_tree_add_51_79_groupi_g43042(csa_tree_add_51_79_groupi_n_2919 ,csa_tree_add_51_79_groupi_n_2692 ,csa_tree_add_51_79_groupi_n_1213);
  or csa_tree_add_51_79_groupi_g43043(csa_tree_add_51_79_groupi_n_2918 ,csa_tree_add_51_79_groupi_n_2645 ,csa_tree_add_51_79_groupi_n_745);
  or csa_tree_add_51_79_groupi_g43044(csa_tree_add_51_79_groupi_n_2917 ,csa_tree_add_51_79_groupi_n_2717 ,csa_tree_add_51_79_groupi_n_1297);
  and csa_tree_add_51_79_groupi_g43045(csa_tree_add_51_79_groupi_n_2916 ,csa_tree_add_51_79_groupi_n_2558 ,csa_tree_add_51_79_groupi_n_2552);
  or csa_tree_add_51_79_groupi_g43046(csa_tree_add_51_79_groupi_n_2915 ,csa_tree_add_51_79_groupi_n_2230 ,csa_tree_add_51_79_groupi_n_1243);
  or csa_tree_add_51_79_groupi_g43047(csa_tree_add_51_79_groupi_n_2914 ,csa_tree_add_51_79_groupi_n_2087 ,csa_tree_add_51_79_groupi_n_1112);
  or csa_tree_add_51_79_groupi_g43048(csa_tree_add_51_79_groupi_n_2913 ,csa_tree_add_51_79_groupi_n_2159 ,csa_tree_add_51_79_groupi_n_1258);
  or csa_tree_add_51_79_groupi_g43049(csa_tree_add_51_79_groupi_n_2912 ,csa_tree_add_51_79_groupi_n_2849 ,csa_tree_add_51_79_groupi_n_1103);
  or csa_tree_add_51_79_groupi_g43050(csa_tree_add_51_79_groupi_n_2911 ,csa_tree_add_51_79_groupi_n_2666 ,csa_tree_add_51_79_groupi_n_1294);
  or csa_tree_add_51_79_groupi_g43051(csa_tree_add_51_79_groupi_n_2910 ,csa_tree_add_51_79_groupi_n_2811 ,csa_tree_add_51_79_groupi_n_1240);
  or csa_tree_add_51_79_groupi_g43052(csa_tree_add_51_79_groupi_n_2909 ,csa_tree_add_51_79_groupi_n_2067 ,csa_tree_add_51_79_groupi_n_1393);
  or csa_tree_add_51_79_groupi_g43053(csa_tree_add_51_79_groupi_n_2908 ,csa_tree_add_51_79_groupi_n_2726 ,csa_tree_add_51_79_groupi_n_1237);
  or csa_tree_add_51_79_groupi_g43054(csa_tree_add_51_79_groupi_n_2907 ,csa_tree_add_51_79_groupi_n_2597 ,csa_tree_add_51_79_groupi_n_1088);
  or csa_tree_add_51_79_groupi_g43055(csa_tree_add_51_79_groupi_n_2906 ,csa_tree_add_51_79_groupi_n_2747 ,csa_tree_add_51_79_groupi_n_1291);
  or csa_tree_add_51_79_groupi_g43056(csa_tree_add_51_79_groupi_n_2905 ,csa_tree_add_51_79_groupi_n_2082 ,csa_tree_add_51_79_groupi_n_1327);
  or csa_tree_add_51_79_groupi_g43057(csa_tree_add_51_79_groupi_n_2904 ,csa_tree_add_51_79_groupi_n_2606 ,csa_tree_add_51_79_groupi_n_1390);
  or csa_tree_add_51_79_groupi_g43058(csa_tree_add_51_79_groupi_n_2903 ,csa_tree_add_51_79_groupi_n_2084 ,csa_tree_add_51_79_groupi_n_1378);
  or csa_tree_add_51_79_groupi_g43059(csa_tree_add_51_79_groupi_n_2902 ,csa_tree_add_51_79_groupi_n_2219 ,csa_tree_add_51_79_groupi_n_1219);
  or csa_tree_add_51_79_groupi_g43060(csa_tree_add_51_79_groupi_n_2901 ,csa_tree_add_51_79_groupi_n_2595 ,csa_tree_add_51_79_groupi_n_1255);
  or csa_tree_add_51_79_groupi_g43061(csa_tree_add_51_79_groupi_n_2900 ,csa_tree_add_51_79_groupi_n_2623 ,csa_tree_add_51_79_groupi_n_1288);
  or csa_tree_add_51_79_groupi_g43062(csa_tree_add_51_79_groupi_n_2899 ,csa_tree_add_51_79_groupi_n_2766 ,csa_tree_add_51_79_groupi_n_1087);
  nor csa_tree_add_51_79_groupi_g43063(csa_tree_add_51_79_groupi_n_2898 ,csa_tree_add_51_79_groupi_n_1755 ,csa_tree_add_51_79_groupi_n_2378);
  nor csa_tree_add_51_79_groupi_g43064(csa_tree_add_51_79_groupi_n_2897 ,csa_tree_add_51_79_groupi_n_1732 ,csa_tree_add_51_79_groupi_n_2377);
  nor csa_tree_add_51_79_groupi_g43065(csa_tree_add_51_79_groupi_n_2896 ,csa_tree_add_51_79_groupi_n_1772 ,csa_tree_add_51_79_groupi_n_2376);
  or csa_tree_add_51_79_groupi_g43066(csa_tree_add_51_79_groupi_n_2895 ,csa_tree_add_51_79_groupi_n_2262 ,csa_tree_add_51_79_groupi_n_1249);
  or csa_tree_add_51_79_groupi_g43067(csa_tree_add_51_79_groupi_n_2894 ,csa_tree_add_51_79_groupi_n_2761 ,csa_tree_add_51_79_groupi_n_1264);
  or csa_tree_add_51_79_groupi_g43068(csa_tree_add_51_79_groupi_n_2893 ,csa_tree_add_51_79_groupi_n_2092 ,csa_tree_add_51_79_groupi_n_1225);
  or csa_tree_add_51_79_groupi_g43069(csa_tree_add_51_79_groupi_n_2892 ,csa_tree_add_51_79_groupi_n_2199 ,csa_tree_add_51_79_groupi_n_1261);
  or csa_tree_add_51_79_groupi_g43070(csa_tree_add_51_79_groupi_n_2891 ,csa_tree_add_51_79_groupi_n_2646 ,csa_tree_add_51_79_groupi_n_1324);
  or csa_tree_add_51_79_groupi_g43071(csa_tree_add_51_79_groupi_n_2890 ,csa_tree_add_51_79_groupi_n_2127 ,csa_tree_add_51_79_groupi_n_1360);
  or csa_tree_add_51_79_groupi_g43072(csa_tree_add_51_79_groupi_n_2889 ,csa_tree_add_51_79_groupi_n_2587 ,csa_tree_add_51_79_groupi_n_1252);
  or csa_tree_add_51_79_groupi_g43073(csa_tree_add_51_79_groupi_n_2888 ,csa_tree_add_51_79_groupi_n_2052 ,csa_tree_add_51_79_groupi_n_1375);
  or csa_tree_add_51_79_groupi_g43074(csa_tree_add_51_79_groupi_n_2887 ,csa_tree_add_51_79_groupi_n_2621 ,csa_tree_add_51_79_groupi_n_1092);
  or csa_tree_add_51_79_groupi_g43075(csa_tree_add_51_79_groupi_n_2886 ,csa_tree_add_51_79_groupi_n_2157 ,csa_tree_add_51_79_groupi_n_1090);
  or csa_tree_add_51_79_groupi_g43076(csa_tree_add_51_79_groupi_n_2885 ,csa_tree_add_51_79_groupi_n_2291 ,csa_tree_add_51_79_groupi_n_1102);
  or csa_tree_add_51_79_groupi_g43078(csa_tree_add_51_79_groupi_n_3373 ,csa_tree_add_51_79_groupi_n_2649 ,csa_tree_add_51_79_groupi_n_1091);
  or csa_tree_add_51_79_groupi_g43079(csa_tree_add_51_79_groupi_n_3372 ,csa_tree_add_51_79_groupi_n_2142 ,csa_tree_add_51_79_groupi_n_1114);
  and csa_tree_add_51_79_groupi_g43080(csa_tree_add_51_79_groupi_n_3370 ,csa_tree_add_51_79_groupi_n_2256 ,csa_tree_add_51_79_groupi_n_1983);
  and csa_tree_add_51_79_groupi_g43081(csa_tree_add_51_79_groupi_n_3368 ,csa_tree_add_51_79_groupi_n_2120 ,csa_tree_add_51_79_groupi_n_1987);
  and csa_tree_add_51_79_groupi_g43082(csa_tree_add_51_79_groupi_n_3366 ,csa_tree_add_51_79_groupi_n_2281 ,csa_tree_add_51_79_groupi_n_1977);
  and csa_tree_add_51_79_groupi_g43083(csa_tree_add_51_79_groupi_n_3364 ,csa_tree_add_51_79_groupi_n_2117 ,csa_tree_add_51_79_groupi_n_2445);
  and csa_tree_add_51_79_groupi_g43084(csa_tree_add_51_79_groupi_n_3362 ,csa_tree_add_51_79_groupi_n_2654 ,csa_tree_add_51_79_groupi_n_2479);
  and csa_tree_add_51_79_groupi_g43085(csa_tree_add_51_79_groupi_n_3360 ,csa_tree_add_51_79_groupi_n_2100 ,csa_tree_add_51_79_groupi_n_2453);
  and csa_tree_add_51_79_groupi_g43086(csa_tree_add_51_79_groupi_n_3358 ,csa_tree_add_51_79_groupi_n_2106 ,csa_tree_add_51_79_groupi_n_1998);
  or csa_tree_add_51_79_groupi_g43087(csa_tree_add_51_79_groupi_n_3357 ,csa_tree_add_51_79_groupi_n_2132 ,csa_tree_add_51_79_groupi_n_1106);
  or csa_tree_add_51_79_groupi_g43088(csa_tree_add_51_79_groupi_n_3356 ,csa_tree_add_51_79_groupi_n_2080 ,csa_tree_add_51_79_groupi_n_1101);
  and csa_tree_add_51_79_groupi_g43089(csa_tree_add_51_79_groupi_n_3354 ,csa_tree_add_51_79_groupi_n_2254 ,csa_tree_add_51_79_groupi_n_1979);
  and csa_tree_add_51_79_groupi_g43090(csa_tree_add_51_79_groupi_n_3352 ,csa_tree_add_51_79_groupi_n_2589 ,csa_tree_add_51_79_groupi_n_1996);
  or csa_tree_add_51_79_groupi_g43091(csa_tree_add_51_79_groupi_n_3351 ,csa_tree_add_51_79_groupi_n_2060 ,csa_tree_add_51_79_groupi_n_1089);
  or csa_tree_add_51_79_groupi_g43092(csa_tree_add_51_79_groupi_n_3350 ,csa_tree_add_51_79_groupi_n_2288 ,csa_tree_add_51_79_groupi_n_1094);
  or csa_tree_add_51_79_groupi_g43093(csa_tree_add_51_79_groupi_n_3349 ,csa_tree_add_51_79_groupi_n_2577 ,csa_tree_add_51_79_groupi_n_1115);
  or csa_tree_add_51_79_groupi_g43094(csa_tree_add_51_79_groupi_n_3348 ,csa_tree_add_51_79_groupi_n_2600 ,csa_tree_add_51_79_groupi_n_1095);
  and csa_tree_add_51_79_groupi_g43095(csa_tree_add_51_79_groupi_n_3346 ,csa_tree_add_51_79_groupi_n_2174 ,csa_tree_add_51_79_groupi_n_1259);
  or csa_tree_add_51_79_groupi_g43096(csa_tree_add_51_79_groupi_n_3345 ,csa_tree_add_51_79_groupi_n_2698 ,csa_tree_add_51_79_groupi_n_1105);
  or csa_tree_add_51_79_groupi_g43097(csa_tree_add_51_79_groupi_n_3344 ,csa_tree_add_51_79_groupi_n_2703 ,csa_tree_add_51_79_groupi_n_1109);
  or csa_tree_add_51_79_groupi_g43098(csa_tree_add_51_79_groupi_n_3343 ,csa_tree_add_51_79_groupi_n_2075 ,csa_tree_add_51_79_groupi_n_1100);
  or csa_tree_add_51_79_groupi_g43099(csa_tree_add_51_79_groupi_n_3342 ,csa_tree_add_51_79_groupi_n_2172 ,csa_tree_add_51_79_groupi_n_1110);
  and csa_tree_add_51_79_groupi_g43100(csa_tree_add_51_79_groupi_n_3340 ,csa_tree_add_51_79_groupi_n_2146 ,csa_tree_add_51_79_groupi_n_1991);
  or csa_tree_add_51_79_groupi_g43101(csa_tree_add_51_79_groupi_n_3339 ,csa_tree_add_51_79_groupi_n_2155 ,csa_tree_add_51_79_groupi_n_1093);
  or csa_tree_add_51_79_groupi_g43102(csa_tree_add_51_79_groupi_n_3338 ,csa_tree_add_51_79_groupi_n_2884 ,csa_tree_add_51_79_groupi_n_1107);
  or csa_tree_add_51_79_groupi_g43105(csa_tree_add_51_79_groupi_n_3337 ,csa_tree_add_51_79_groupi_n_2618 ,csa_tree_add_51_79_groupi_n_1113);
  and csa_tree_add_51_79_groupi_g43106(csa_tree_add_51_79_groupi_n_3335 ,csa_tree_add_51_79_groupi_n_2263 ,csa_tree_add_51_79_groupi_n_1981);
  and csa_tree_add_51_79_groupi_g43107(csa_tree_add_51_79_groupi_n_3334 ,csa_tree_add_51_79_groupi_n_1844 ,csa_tree_add_51_79_groupi_n_1450);
  or csa_tree_add_51_79_groupi_g43108(csa_tree_add_51_79_groupi_n_3333 ,csa_tree_add_51_79_groupi_n_807 ,csa_tree_add_51_79_groupi_n_748);
  or csa_tree_add_51_79_groupi_g43109(csa_tree_add_51_79_groupi_n_3332 ,csa_tree_add_51_79_groupi_n_848 ,csa_tree_add_51_79_groupi_n_682);
  or csa_tree_add_51_79_groupi_g43110(csa_tree_add_51_79_groupi_n_3331 ,csa_tree_add_51_79_groupi_n_846 ,csa_tree_add_51_79_groupi_n_2539);
  and csa_tree_add_51_79_groupi_g43111(csa_tree_add_51_79_groupi_n_3330 ,csa_tree_add_51_79_groupi_n_1964 ,csa_tree_add_51_79_groupi_n_1450);
  or csa_tree_add_51_79_groupi_g43112(csa_tree_add_51_79_groupi_n_3329 ,csa_tree_add_51_79_groupi_n_842 ,csa_tree_add_51_79_groupi_n_1297);
  or csa_tree_add_51_79_groupi_g43113(csa_tree_add_51_79_groupi_n_3328 ,csa_tree_add_51_79_groupi_n_840 ,csa_tree_add_51_79_groupi_n_658);
  and csa_tree_add_51_79_groupi_g43114(csa_tree_add_51_79_groupi_n_3327 ,csa_tree_add_51_79_groupi_n_1927 ,csa_tree_add_51_79_groupi_n_1462);
  or csa_tree_add_51_79_groupi_g43115(csa_tree_add_51_79_groupi_n_3326 ,csa_tree_add_51_79_groupi_n_807 ,csa_tree_add_51_79_groupi_n_697);
  or csa_tree_add_51_79_groupi_g43116(csa_tree_add_51_79_groupi_n_3325 ,csa_tree_add_51_79_groupi_n_807 ,csa_tree_add_51_79_groupi_n_1309);
  or csa_tree_add_51_79_groupi_g43117(csa_tree_add_51_79_groupi_n_3324 ,csa_tree_add_51_79_groupi_n_838 ,csa_tree_add_51_79_groupi_n_700);
  or csa_tree_add_51_79_groupi_g43118(csa_tree_add_51_79_groupi_n_3323 ,csa_tree_add_51_79_groupi_n_570 ,csa_tree_add_51_79_groupi_n_1387);
  or csa_tree_add_51_79_groupi_g43119(csa_tree_add_51_79_groupi_n_3322 ,csa_tree_add_51_79_groupi_n_582 ,csa_tree_add_51_79_groupi_n_712);
  or csa_tree_add_51_79_groupi_g43120(csa_tree_add_51_79_groupi_n_3321 ,csa_tree_add_51_79_groupi_n_567 ,csa_tree_add_51_79_groupi_n_1270);
  or csa_tree_add_51_79_groupi_g43121(csa_tree_add_51_79_groupi_n_3320 ,csa_tree_add_51_79_groupi_n_1932 ,csa_tree_add_51_79_groupi_n_1457);
  or csa_tree_add_51_79_groupi_g43122(csa_tree_add_51_79_groupi_n_3319 ,csa_tree_add_51_79_groupi_n_838 ,csa_tree_add_51_79_groupi_n_1357);
  or csa_tree_add_51_79_groupi_g43123(csa_tree_add_51_79_groupi_n_3318 ,csa_tree_add_51_79_groupi_n_848 ,csa_tree_add_51_79_groupi_n_1471);
  and csa_tree_add_51_79_groupi_g43124(csa_tree_add_51_79_groupi_n_3317 ,csa_tree_add_51_79_groupi_n_1867 ,csa_tree_add_51_79_groupi_n_727);
  or csa_tree_add_51_79_groupi_g43125(csa_tree_add_51_79_groupi_n_3316 ,csa_tree_add_51_79_groupi_n_846 ,csa_tree_add_51_79_groupi_n_724);
  or csa_tree_add_51_79_groupi_g43126(csa_tree_add_51_79_groupi_n_3315 ,csa_tree_add_51_79_groupi_n_807 ,csa_tree_add_51_79_groupi_n_1432);
  or csa_tree_add_51_79_groupi_g43127(csa_tree_add_51_79_groupi_n_3314 ,csa_tree_add_51_79_groupi_n_848 ,csa_tree_add_51_79_groupi_n_1351);
  or csa_tree_add_51_79_groupi_g43128(csa_tree_add_51_79_groupi_n_3313 ,csa_tree_add_51_79_groupi_n_568 ,csa_tree_add_51_79_groupi_n_673);
  or csa_tree_add_51_79_groupi_g43129(csa_tree_add_51_79_groupi_n_3312 ,csa_tree_add_51_79_groupi_n_846 ,csa_tree_add_51_79_groupi_n_1279);
  or csa_tree_add_51_79_groupi_g43130(csa_tree_add_51_79_groupi_n_3311 ,csa_tree_add_51_79_groupi_n_807 ,csa_tree_add_51_79_groupi_n_1460);
  or csa_tree_add_51_79_groupi_g43131(csa_tree_add_51_79_groupi_n_3310 ,csa_tree_add_51_79_groupi_n_576 ,csa_tree_add_51_79_groupi_n_1448);
  or csa_tree_add_51_79_groupi_g43132(csa_tree_add_51_79_groupi_n_3308 ,csa_tree_add_51_79_groupi_n_1912 ,csa_tree_add_51_79_groupi_n_2514);
  or csa_tree_add_51_79_groupi_g43133(csa_tree_add_51_79_groupi_n_3307 ,csa_tree_add_51_79_groupi_n_798 ,csa_tree_add_51_79_groupi_n_676);
  or csa_tree_add_51_79_groupi_g43134(csa_tree_add_51_79_groupi_n_3305 ,csa_tree_add_51_79_groupi_n_1830 ,csa_tree_add_51_79_groupi_n_2534);
  or csa_tree_add_51_79_groupi_g43135(csa_tree_add_51_79_groupi_n_3303 ,csa_tree_add_51_79_groupi_n_1902 ,csa_tree_add_51_79_groupi_n_1471);
  or csa_tree_add_51_79_groupi_g43136(csa_tree_add_51_79_groupi_n_3301 ,csa_tree_add_51_79_groupi_n_1847 ,csa_tree_add_51_79_groupi_n_1122);
  or csa_tree_add_51_79_groupi_g43137(csa_tree_add_51_79_groupi_n_3299 ,csa_tree_add_51_79_groupi_n_1950 ,csa_tree_add_51_79_groupi_n_2525);
  or csa_tree_add_51_79_groupi_g43138(csa_tree_add_51_79_groupi_n_3298 ,csa_tree_add_51_79_groupi_n_844 ,csa_tree_add_51_79_groupi_n_1467);
  and csa_tree_add_51_79_groupi_g43139(csa_tree_add_51_79_groupi_n_3297 ,csa_tree_add_51_79_groupi_n_1957 ,csa_tree_add_51_79_groupi_n_2524);
  or csa_tree_add_51_79_groupi_g43140(csa_tree_add_51_79_groupi_n_3295 ,csa_tree_add_51_79_groupi_n_1874 ,csa_tree_add_51_79_groupi_n_1467);
  or csa_tree_add_51_79_groupi_g43141(csa_tree_add_51_79_groupi_n_3294 ,csa_tree_add_51_79_groupi_n_852 ,csa_tree_add_51_79_groupi_n_736);
  or csa_tree_add_51_79_groupi_g43142(csa_tree_add_51_79_groupi_n_3293 ,csa_tree_add_51_79_groupi_n_561 ,csa_tree_add_51_79_groupi_n_2534);
  or csa_tree_add_51_79_groupi_g43143(csa_tree_add_51_79_groupi_n_3291 ,csa_tree_add_51_79_groupi_n_1924 ,csa_tree_add_51_79_groupi_n_2534);
  and csa_tree_add_51_79_groupi_g43144(csa_tree_add_51_79_groupi_n_3290 ,csa_tree_add_51_79_groupi_n_1926 ,csa_tree_add_51_79_groupi_n_2537);
  or csa_tree_add_51_79_groupi_g43145(csa_tree_add_51_79_groupi_n_3289 ,csa_tree_add_51_79_groupi_n_836 ,csa_tree_add_51_79_groupi_n_1372);
  and csa_tree_add_51_79_groupi_g43146(csa_tree_add_51_79_groupi_n_3288 ,csa_tree_add_51_79_groupi_n_1892 ,csa_tree_add_51_79_groupi_n_1456);
  or csa_tree_add_51_79_groupi_g43147(csa_tree_add_51_79_groupi_n_3287 ,csa_tree_add_51_79_groupi_n_810 ,csa_tree_add_51_79_groupi_n_1435);
  or csa_tree_add_51_79_groupi_g43148(csa_tree_add_51_79_groupi_n_3285 ,csa_tree_add_51_79_groupi_n_1911 ,csa_tree_add_51_79_groupi_n_1122);
  or csa_tree_add_51_79_groupi_g43149(csa_tree_add_51_79_groupi_n_3283 ,csa_tree_add_51_79_groupi_n_1949 ,csa_tree_add_51_79_groupi_n_1457);
  xnor csa_tree_add_51_79_groupi_g43150(csa_tree_add_51_79_groupi_n_3282 ,csa_tree_add_51_79_groupi_n_1785 ,csa_tree_add_51_79_groupi_n_1779);
  and csa_tree_add_51_79_groupi_g43151(csa_tree_add_51_79_groupi_n_3281 ,csa_tree_add_51_79_groupi_n_1944 ,csa_tree_add_51_79_groupi_n_2530);
  and csa_tree_add_51_79_groupi_g43152(csa_tree_add_51_79_groupi_n_3280 ,csa_tree_add_51_79_groupi_n_1923 ,csa_tree_add_51_79_groupi_n_1124);
  or csa_tree_add_51_79_groupi_g43153(csa_tree_add_51_79_groupi_n_3278 ,csa_tree_add_51_79_groupi_n_1836 ,csa_tree_add_51_79_groupi_n_1454);
  or csa_tree_add_51_79_groupi_g43154(csa_tree_add_51_79_groupi_n_3277 ,csa_tree_add_51_79_groupi_n_573 ,csa_tree_add_51_79_groupi_n_1267);
  or csa_tree_add_51_79_groupi_g43155(csa_tree_add_51_79_groupi_n_3275 ,csa_tree_add_51_79_groupi_n_1938 ,csa_tree_add_51_79_groupi_n_1448);
  or csa_tree_add_51_79_groupi_g43156(csa_tree_add_51_79_groupi_n_3274 ,csa_tree_add_51_79_groupi_n_850 ,csa_tree_add_51_79_groupi_n_1285);
  or csa_tree_add_51_79_groupi_g43157(csa_tree_add_51_79_groupi_n_3273 ,csa_tree_add_51_79_groupi_n_1832 ,csa_tree_add_51_79_groupi_n_1457);
  or csa_tree_add_51_79_groupi_g43158(csa_tree_add_51_79_groupi_n_3271 ,csa_tree_add_51_79_groupi_n_1884 ,csa_tree_add_51_79_groupi_n_1460);
  or csa_tree_add_51_79_groupi_g43159(csa_tree_add_51_79_groupi_n_3270 ,csa_tree_add_51_79_groupi_n_844 ,csa_tree_add_51_79_groupi_n_685);
  and csa_tree_add_51_79_groupi_g43160(csa_tree_add_51_79_groupi_n_3269 ,csa_tree_add_51_79_groupi_n_1850 ,csa_tree_add_51_79_groupi_n_2530);
  or csa_tree_add_51_79_groupi_g43161(csa_tree_add_51_79_groupi_n_3268 ,csa_tree_add_51_79_groupi_n_1826 ,csa_tree_add_51_79_groupi_n_2534);
  or csa_tree_add_51_79_groupi_g43162(csa_tree_add_51_79_groupi_n_3267 ,csa_tree_add_51_79_groupi_n_798 ,csa_tree_add_51_79_groupi_n_1291);
  and csa_tree_add_51_79_groupi_g43163(csa_tree_add_51_79_groupi_n_3266 ,csa_tree_add_51_79_groupi_n_1877 ,csa_tree_add_51_79_groupi_n_1459);
  or csa_tree_add_51_79_groupi_g43164(csa_tree_add_51_79_groupi_n_3265 ,csa_tree_add_51_79_groupi_n_798 ,csa_tree_add_51_79_groupi_n_730);
  and csa_tree_add_51_79_groupi_g43165(csa_tree_add_51_79_groupi_n_3264 ,csa_tree_add_51_79_groupi_n_1870 ,csa_tree_add_51_79_groupi_n_2538);
  and csa_tree_add_51_79_groupi_g43166(csa_tree_add_51_79_groupi_n_3263 ,csa_tree_add_51_79_groupi_n_1947 ,csa_tree_add_51_79_groupi_n_670);
  or csa_tree_add_51_79_groupi_g43167(csa_tree_add_51_79_groupi_n_3262 ,csa_tree_add_51_79_groupi_n_579 ,csa_tree_add_51_79_groupi_n_1423);
  or csa_tree_add_51_79_groupi_g43168(csa_tree_add_51_79_groupi_n_3261 ,csa_tree_add_51_79_groupi_n_810 ,csa_tree_add_51_79_groupi_n_751);
  or csa_tree_add_51_79_groupi_g43169(csa_tree_add_51_79_groupi_n_3259 ,csa_tree_add_51_79_groupi_n_1959 ,csa_tree_add_51_79_groupi_n_1471);
  or csa_tree_add_51_79_groupi_g43170(csa_tree_add_51_79_groupi_n_3258 ,csa_tree_add_51_79_groupi_n_844 ,csa_tree_add_51_79_groupi_n_739);
  or csa_tree_add_51_79_groupi_g43171(csa_tree_add_51_79_groupi_n_3257 ,csa_tree_add_51_79_groupi_n_840 ,csa_tree_add_51_79_groupi_n_1378);
  or csa_tree_add_51_79_groupi_g43172(csa_tree_add_51_79_groupi_n_3256 ,csa_tree_add_51_79_groupi_n_1931 ,csa_tree_add_51_79_groupi_n_2519);
  or csa_tree_add_51_79_groupi_g43173(csa_tree_add_51_79_groupi_n_3254 ,csa_tree_add_51_79_groupi_n_1871 ,csa_tree_add_51_79_groupi_n_2516);
  or csa_tree_add_51_79_groupi_g43174(csa_tree_add_51_79_groupi_n_3253 ,csa_tree_add_51_79_groupi_n_574 ,csa_tree_add_51_79_groupi_n_1303);
  or csa_tree_add_51_79_groupi_g43175(csa_tree_add_51_79_groupi_n_3251 ,csa_tree_add_51_79_groupi_n_1901 ,csa_tree_add_51_79_groupi_n_1084);
  and csa_tree_add_51_79_groupi_g43176(csa_tree_add_51_79_groupi_n_3250 ,csa_tree_add_51_79_groupi_n_1825 ,csa_tree_add_51_79_groupi_n_1456);
  or csa_tree_add_51_79_groupi_g43177(csa_tree_add_51_79_groupi_n_3248 ,csa_tree_add_51_79_groupi_n_1898 ,csa_tree_add_51_79_groupi_n_1460);
  and csa_tree_add_51_79_groupi_g43178(csa_tree_add_51_79_groupi_n_3247 ,csa_tree_add_51_79_groupi_n_1961 ,csa_tree_add_51_79_groupi_n_1450);
  and csa_tree_add_51_79_groupi_g43179(csa_tree_add_51_79_groupi_n_3246 ,csa_tree_add_51_79_groupi_n_1855 ,csa_tree_add_51_79_groupi_n_1456);
  and csa_tree_add_51_79_groupi_g43180(csa_tree_add_51_79_groupi_n_3245 ,csa_tree_add_51_79_groupi_n_1948 ,csa_tree_add_51_79_groupi_n_718);
  and csa_tree_add_51_79_groupi_g43181(csa_tree_add_51_79_groupi_n_3244 ,csa_tree_add_51_79_groupi_n_1916 ,csa_tree_add_51_79_groupi_n_1450);
  and csa_tree_add_51_79_groupi_g43182(csa_tree_add_51_79_groupi_n_3243 ,csa_tree_add_51_79_groupi_n_1909 ,csa_tree_add_51_79_groupi_n_727);
  and csa_tree_add_51_79_groupi_g43183(csa_tree_add_51_79_groupi_n_3242 ,csa_tree_add_51_79_groupi_n_1900 ,csa_tree_add_51_79_groupi_n_1462);
  or csa_tree_add_51_79_groupi_g43184(csa_tree_add_51_79_groupi_n_3240 ,csa_tree_add_51_79_groupi_n_1833 ,csa_tree_add_51_79_groupi_n_1471);
  or csa_tree_add_51_79_groupi_g43185(csa_tree_add_51_79_groupi_n_3239 ,csa_tree_add_51_79_groupi_n_1860 ,csa_tree_add_51_79_groupi_n_2534);
  or csa_tree_add_51_79_groupi_g43186(csa_tree_add_51_79_groupi_n_3237 ,csa_tree_add_51_79_groupi_n_1910 ,csa_tree_add_51_79_groupi_n_1467);
  and csa_tree_add_51_79_groupi_g43187(csa_tree_add_51_79_groupi_n_3236 ,csa_tree_add_51_79_groupi_n_1919 ,csa_tree_add_51_79_groupi_n_1124);
  or csa_tree_add_51_79_groupi_g43188(csa_tree_add_51_79_groupi_n_3234 ,csa_tree_add_51_79_groupi_n_1907 ,csa_tree_add_51_79_groupi_n_1122);
  and csa_tree_add_51_79_groupi_g43189(csa_tree_add_51_79_groupi_n_3233 ,csa_tree_add_51_79_groupi_n_1954 ,csa_tree_add_51_79_groupi_n_1456);
  or csa_tree_add_51_79_groupi_g43190(csa_tree_add_51_79_groupi_n_3231 ,csa_tree_add_51_79_groupi_n_1866 ,csa_tree_add_51_79_groupi_n_1467);
  or csa_tree_add_51_79_groupi_g43191(csa_tree_add_51_79_groupi_n_3230 ,csa_tree_add_51_79_groupi_n_564 ,csa_tree_add_51_79_groupi_n_1327);
  or csa_tree_add_51_79_groupi_g43192(csa_tree_add_51_79_groupi_n_3228 ,csa_tree_add_51_79_groupi_n_1928 ,csa_tree_add_51_79_groupi_n_2534);
  or csa_tree_add_51_79_groupi_g43193(csa_tree_add_51_79_groupi_n_3226 ,csa_tree_add_51_79_groupi_n_1872 ,csa_tree_add_51_79_groupi_n_1467);
  or csa_tree_add_51_79_groupi_g43194(csa_tree_add_51_79_groupi_n_3225 ,csa_tree_add_51_79_groupi_n_842 ,csa_tree_add_51_79_groupi_n_1321);
  or csa_tree_add_51_79_groupi_g43195(csa_tree_add_51_79_groupi_n_3224 ,csa_tree_add_51_79_groupi_n_810 ,csa_tree_add_51_79_groupi_n_1078);
  or csa_tree_add_51_79_groupi_g43196(csa_tree_add_51_79_groupi_n_3223 ,csa_tree_add_51_79_groupi_n_850 ,csa_tree_add_51_79_groupi_n_1381);
  or csa_tree_add_51_79_groupi_g43197(csa_tree_add_51_79_groupi_n_3222 ,csa_tree_add_51_79_groupi_n_810 ,csa_tree_add_51_79_groupi_n_1426);
  or csa_tree_add_51_79_groupi_g43198(csa_tree_add_51_79_groupi_n_3221 ,csa_tree_add_51_79_groupi_n_850 ,csa_tree_add_51_79_groupi_n_1339);
  or csa_tree_add_51_79_groupi_g43199(csa_tree_add_51_79_groupi_n_3220 ,csa_tree_add_51_79_groupi_n_585 ,csa_tree_add_51_79_groupi_n_1414);
  or csa_tree_add_51_79_groupi_g43200(csa_tree_add_51_79_groupi_n_3219 ,csa_tree_add_51_79_groupi_n_798 ,csa_tree_add_51_79_groupi_n_706);
  or csa_tree_add_51_79_groupi_g43201(csa_tree_add_51_79_groupi_n_3218 ,csa_tree_add_51_79_groupi_n_842 ,csa_tree_add_51_79_groupi_n_1363);
  or csa_tree_add_51_79_groupi_g43202(csa_tree_add_51_79_groupi_n_3217 ,csa_tree_add_51_79_groupi_n_810 ,csa_tree_add_51_79_groupi_n_1315);
  and csa_tree_add_51_79_groupi_g43203(csa_tree_add_51_79_groupi_n_3216 ,csa_tree_add_51_79_groupi_n_1890 ,csa_tree_add_51_79_groupi_n_1450);
  or csa_tree_add_51_79_groupi_g43204(csa_tree_add_51_79_groupi_n_3214 ,csa_tree_add_51_79_groupi_n_1887 ,csa_tree_add_51_79_groupi_n_1471);
  or csa_tree_add_51_79_groupi_g43205(csa_tree_add_51_79_groupi_n_3212 ,csa_tree_add_51_79_groupi_n_1952 ,csa_tree_add_51_79_groupi_n_2523);
  or csa_tree_add_51_79_groupi_g43206(csa_tree_add_51_79_groupi_n_3211 ,csa_tree_add_51_79_groupi_n_571 ,csa_tree_add_51_79_groupi_n_694);
  and csa_tree_add_51_79_groupi_g43207(csa_tree_add_51_79_groupi_n_3210 ,csa_tree_add_51_79_groupi_n_1888 ,csa_tree_add_51_79_groupi_n_670);
  or csa_tree_add_51_79_groupi_g43208(csa_tree_add_51_79_groupi_n_3209 ,csa_tree_add_51_79_groupi_n_838 ,csa_tree_add_51_79_groupi_n_1122);
  or csa_tree_add_51_79_groupi_g43209(csa_tree_add_51_79_groupi_n_3208 ,csa_tree_add_51_79_groupi_n_852 ,csa_tree_add_51_79_groupi_n_1441);
  or csa_tree_add_51_79_groupi_g43210(csa_tree_add_51_79_groupi_n_3207 ,csa_tree_add_51_79_groupi_n_798 ,csa_tree_add_51_79_groupi_n_1457);
  or csa_tree_add_51_79_groupi_g43211(csa_tree_add_51_79_groupi_n_3206 ,csa_tree_add_51_79_groupi_n_840 ,csa_tree_add_51_79_groupi_n_1333);
  or csa_tree_add_51_79_groupi_g43212(csa_tree_add_51_79_groupi_n_3205 ,csa_tree_add_51_79_groupi_n_836 ,csa_tree_add_51_79_groupi_n_1345);
  and csa_tree_add_51_79_groupi_g43213(csa_tree_add_51_79_groupi_n_3204 ,csa_tree_add_51_79_groupi_n_1848 ,csa_tree_add_51_79_groupi_n_727);
  or csa_tree_add_51_79_groupi_g43214(csa_tree_add_51_79_groupi_n_3203 ,csa_tree_add_51_79_groupi_n_852 ,csa_tree_add_51_79_groupi_n_1408);
  or csa_tree_add_51_79_groupi_g43215(csa_tree_add_51_79_groupi_n_3202 ,csa_tree_add_51_79_groupi_n_562 ,csa_tree_add_51_79_groupi_n_709);
  or csa_tree_add_51_79_groupi_g43216(csa_tree_add_51_79_groupi_n_3201 ,csa_tree_add_51_79_groupi_n_836 ,csa_tree_add_51_79_groupi_n_1080);
  or csa_tree_add_51_79_groupi_g43217(csa_tree_add_51_79_groupi_n_3200 ,csa_tree_add_51_79_groupi_n_583 ,csa_tree_add_51_79_groupi_n_1399);
  or csa_tree_add_51_79_groupi_g43218(csa_tree_add_51_79_groupi_n_3199 ,csa_tree_add_51_79_groupi_n_565 ,csa_tree_add_51_79_groupi_n_1082);
  or csa_tree_add_51_79_groupi_g43219(csa_tree_add_51_79_groupi_n_3198 ,csa_tree_add_51_79_groupi_n_580 ,csa_tree_add_51_79_groupi_n_1454);
  or csa_tree_add_51_79_groupi_g43220(csa_tree_add_51_79_groupi_n_3196 ,csa_tree_add_51_79_groupi_n_1895 ,csa_tree_add_51_79_groupi_n_1460);
  or csa_tree_add_51_79_groupi_g43221(csa_tree_add_51_79_groupi_n_3195 ,csa_tree_add_51_79_groupi_n_577 ,csa_tree_add_51_79_groupi_n_745);
  or csa_tree_add_51_79_groupi_g43222(csa_tree_add_51_79_groupi_n_3194 ,csa_tree_add_51_79_groupi_n_586 ,csa_tree_add_51_79_groupi_n_1396);
  and csa_tree_add_51_79_groupi_g43223(csa_tree_add_51_79_groupi_n_3193 ,csa_tree_add_51_79_groupi_n_1967 ,csa_tree_add_51_79_groupi_n_2537);
  and csa_tree_add_51_79_groupi_g43224(csa_tree_add_51_79_groupi_n_3192 ,csa_tree_add_51_79_groupi_n_1827 ,csa_tree_add_51_79_groupi_n_2530);
  and csa_tree_add_51_79_groupi_g43225(csa_tree_add_51_79_groupi_n_3191 ,csa_tree_add_51_79_groupi_n_1829 ,csa_tree_add_51_79_groupi_n_1462);
  or csa_tree_add_51_79_groupi_g43226(csa_tree_add_51_79_groupi_n_3190 ,csa_tree_add_51_79_groupi_n_1966 ,csa_tree_add_51_79_groupi_n_1418);
  or csa_tree_add_51_79_groupi_g43227(csa_tree_add_51_79_groupi_n_3189 ,csa_tree_add_51_79_groupi_n_2372 ,csa_tree_add_51_79_groupi_n_1346);
  or csa_tree_add_51_79_groupi_g43228(csa_tree_add_51_79_groupi_n_3188 ,csa_tree_add_51_79_groupi_n_2362 ,csa_tree_add_51_79_groupi_n_1238);
  or csa_tree_add_51_79_groupi_g43229(csa_tree_add_51_79_groupi_n_3187 ,csa_tree_add_51_79_groupi_n_1807 ,csa_tree_add_51_79_groupi_n_1244);
  or csa_tree_add_51_79_groupi_g43230(csa_tree_add_51_79_groupi_n_3186 ,csa_tree_add_51_79_groupi_n_1788 ,csa_tree_add_51_79_groupi_n_1223);
  or csa_tree_add_51_79_groupi_g43231(csa_tree_add_51_79_groupi_n_3185 ,csa_tree_add_51_79_groupi_n_1792 ,csa_tree_add_51_79_groupi_n_1328);
  or csa_tree_add_51_79_groupi_g43232(csa_tree_add_51_79_groupi_n_3184 ,csa_tree_add_51_79_groupi_n_1824 ,csa_tree_add_51_79_groupi_n_1229);
  or csa_tree_add_51_79_groupi_g43233(csa_tree_add_51_79_groupi_n_3183 ,csa_tree_add_51_79_groupi_n_2345 ,csa_tree_add_51_79_groupi_n_1436);
  or csa_tree_add_51_79_groupi_g43234(csa_tree_add_51_79_groupi_n_3182 ,csa_tree_add_51_79_groupi_n_1808 ,csa_tree_add_51_79_groupi_n_1322);
  or csa_tree_add_51_79_groupi_g43235(csa_tree_add_51_79_groupi_n_3181 ,csa_tree_add_51_79_groupi_n_2342 ,csa_tree_add_51_79_groupi_n_1220);
  or csa_tree_add_51_79_groupi_g43236(csa_tree_add_51_79_groupi_n_3180 ,csa_tree_add_51_79_groupi_n_1820 ,csa_tree_add_51_79_groupi_n_1253);
  or csa_tree_add_51_79_groupi_g43237(csa_tree_add_51_79_groupi_n_3179 ,csa_tree_add_51_79_groupi_n_1891 ,csa_tree_add_51_79_groupi_n_1211);
  or csa_tree_add_51_79_groupi_g43238(csa_tree_add_51_79_groupi_n_3178 ,csa_tree_add_51_79_groupi_n_1812 ,csa_tree_add_51_79_groupi_n_1241);
  or csa_tree_add_51_79_groupi_g43239(csa_tree_add_51_79_groupi_n_3177 ,csa_tree_add_51_79_groupi_n_1837 ,csa_tree_add_51_79_groupi_n_1442);
  or csa_tree_add_51_79_groupi_g43240(csa_tree_add_51_79_groupi_n_3176 ,csa_tree_add_51_79_groupi_n_1811 ,csa_tree_add_51_79_groupi_n_1256);
  or csa_tree_add_51_79_groupi_g43241(csa_tree_add_51_79_groupi_n_3175 ,csa_tree_add_51_79_groupi_n_1798 ,csa_tree_add_51_79_groupi_n_1316);
  or csa_tree_add_51_79_groupi_g43242(csa_tree_add_51_79_groupi_n_3174 ,csa_tree_add_51_79_groupi_n_2364 ,csa_tree_add_51_79_groupi_n_1373);
  or csa_tree_add_51_79_groupi_g43243(csa_tree_add_51_79_groupi_n_3173 ,csa_tree_add_51_79_groupi_n_1790 ,csa_tree_add_51_79_groupi_n_1235);
  or csa_tree_add_51_79_groupi_g43244(csa_tree_add_51_79_groupi_n_3172 ,csa_tree_add_51_79_groupi_n_2349 ,csa_tree_add_51_79_groupi_n_1262);
  or csa_tree_add_51_79_groupi_g43245(csa_tree_add_51_79_groupi_n_3171 ,csa_tree_add_51_79_groupi_n_2422 ,csa_tree_add_51_79_groupi_n_1403);
  or csa_tree_add_51_79_groupi_g43246(csa_tree_add_51_79_groupi_n_3170 ,csa_tree_add_51_79_groupi_n_1809 ,csa_tree_add_51_79_groupi_n_1247);
  or csa_tree_add_51_79_groupi_g43247(csa_tree_add_51_79_groupi_n_3169 ,in10[0] ,csa_tree_add_51_79_groupi_n_1537);
  or csa_tree_add_51_79_groupi_g43248(csa_tree_add_51_79_groupi_n_3168 ,in2[0] ,csa_tree_add_51_79_groupi_n_1610);
  or csa_tree_add_51_79_groupi_g43249(csa_tree_add_51_79_groupi_n_3167 ,in18[0] ,csa_tree_add_51_79_groupi_n_1601);
  or csa_tree_add_51_79_groupi_g43250(csa_tree_add_51_79_groupi_n_3166 ,csa_tree_add_51_79_groupi_n_2418 ,csa_tree_add_51_79_groupi_n_1400);
  or csa_tree_add_51_79_groupi_g43251(csa_tree_add_51_79_groupi_n_3165 ,csa_tree_add_51_79_groupi_n_1882 ,csa_tree_add_51_79_groupi_n_1226);
  or csa_tree_add_51_79_groupi_g43252(csa_tree_add_51_79_groupi_n_3164 ,in6[0] ,csa_tree_add_51_79_groupi_n_1617);
  or csa_tree_add_51_79_groupi_g43253(csa_tree_add_51_79_groupi_n_3163 ,csa_tree_add_51_79_groupi_n_1804 ,csa_tree_add_51_79_groupi_n_1298);
  or csa_tree_add_51_79_groupi_g43254(csa_tree_add_51_79_groupi_n_3162 ,in8[0] ,csa_tree_add_51_79_groupi_n_1607);
  or csa_tree_add_51_79_groupi_g43255(csa_tree_add_51_79_groupi_n_3161 ,csa_tree_add_51_79_groupi_n_1805 ,csa_tree_add_51_79_groupi_n_1280);
  or csa_tree_add_51_79_groupi_g43256(csa_tree_add_51_79_groupi_n_3160 ,in16[0] ,csa_tree_add_51_79_groupi_n_1612);
  or csa_tree_add_51_79_groupi_g43257(csa_tree_add_51_79_groupi_n_3159 ,csa_tree_add_51_79_groupi_n_2363 ,csa_tree_add_51_79_groupi_n_1310);
  not csa_tree_add_51_79_groupi_g43258(csa_tree_add_51_79_groupi_n_2795 ,csa_tree_add_51_79_groupi_n_2794);
  not csa_tree_add_51_79_groupi_g43259(csa_tree_add_51_79_groupi_n_2773 ,csa_tree_add_51_79_groupi_n_2772);
  not csa_tree_add_51_79_groupi_g43260(csa_tree_add_51_79_groupi_n_2655 ,csa_tree_add_51_79_groupi_n_2654);
  not csa_tree_add_51_79_groupi_g43261(csa_tree_add_51_79_groupi_n_2590 ,csa_tree_add_51_79_groupi_n_2589);
  not csa_tree_add_51_79_groupi_g43262(csa_tree_add_51_79_groupi_n_2569 ,csa_tree_add_51_79_groupi_n_2568);
  not csa_tree_add_51_79_groupi_g43263(csa_tree_add_51_79_groupi_n_2564 ,csa_tree_add_51_79_groupi_n_2563);
  not csa_tree_add_51_79_groupi_g43264(csa_tree_add_51_79_groupi_n_2560 ,csa_tree_add_51_79_groupi_n_2559);
  not csa_tree_add_51_79_groupi_g43265(csa_tree_add_51_79_groupi_n_2549 ,csa_tree_add_51_79_groupi_n_2548);
  not csa_tree_add_51_79_groupi_g43266(csa_tree_add_51_79_groupi_n_2546 ,csa_tree_add_51_79_groupi_n_2545);
  not csa_tree_add_51_79_groupi_g43267(csa_tree_add_51_79_groupi_n_2542 ,csa_tree_add_51_79_groupi_n_2543);
  not csa_tree_add_51_79_groupi_g43269(csa_tree_add_51_79_groupi_n_2538 ,csa_tree_add_51_79_groupi_n_2539);
  buf csa_tree_add_51_79_groupi_g43270(csa_tree_add_51_79_groupi_n_2537 ,csa_tree_add_51_79_groupi_n_2535);
  not csa_tree_add_51_79_groupi_g43271(csa_tree_add_51_79_groupi_n_2536 ,csa_tree_add_51_79_groupi_n_2535);
  buf csa_tree_add_51_79_groupi_g43272(csa_tree_add_51_79_groupi_n_2534 ,csa_tree_add_51_79_groupi_n_2532);
  not csa_tree_add_51_79_groupi_g43273(csa_tree_add_51_79_groupi_n_2533 ,csa_tree_add_51_79_groupi_n_2532);
  buf csa_tree_add_51_79_groupi_g43276(csa_tree_add_51_79_groupi_n_2530 ,csa_tree_add_51_79_groupi_n_2528);
  not csa_tree_add_51_79_groupi_g43277(csa_tree_add_51_79_groupi_n_2529 ,csa_tree_add_51_79_groupi_n_2528);
  not csa_tree_add_51_79_groupi_g43281(csa_tree_add_51_79_groupi_n_2524 ,csa_tree_add_51_79_groupi_n_2525);
  not csa_tree_add_51_79_groupi_g43282(csa_tree_add_51_79_groupi_n_2522 ,csa_tree_add_51_79_groupi_n_2523);
  not csa_tree_add_51_79_groupi_g43287(csa_tree_add_51_79_groupi_n_2518 ,csa_tree_add_51_79_groupi_n_2519);
  not csa_tree_add_51_79_groupi_g43289(csa_tree_add_51_79_groupi_n_2515 ,csa_tree_add_51_79_groupi_n_2516);
  not csa_tree_add_51_79_groupi_g43290(csa_tree_add_51_79_groupi_n_2513 ,csa_tree_add_51_79_groupi_n_2514);
  not csa_tree_add_51_79_groupi_g43294(csa_tree_add_51_79_groupi_n_2510 ,csa_tree_add_51_79_groupi_n_2508);
  not csa_tree_add_51_79_groupi_g43299(csa_tree_add_51_79_groupi_n_2505 ,csa_tree_add_51_79_groupi_n_2503);
  not csa_tree_add_51_79_groupi_g43304(csa_tree_add_51_79_groupi_n_2500 ,csa_tree_add_51_79_groupi_n_2498);
  not csa_tree_add_51_79_groupi_g43307(csa_tree_add_51_79_groupi_n_2497 ,csa_tree_add_51_79_groupi_n_2495);
  not csa_tree_add_51_79_groupi_g43310(csa_tree_add_51_79_groupi_n_2494 ,csa_tree_add_51_79_groupi_n_2492);
  not csa_tree_add_51_79_groupi_g43313(csa_tree_add_51_79_groupi_n_2491 ,csa_tree_add_51_79_groupi_n_2489);
  not csa_tree_add_51_79_groupi_g43318(csa_tree_add_51_79_groupi_n_2486 ,csa_tree_add_51_79_groupi_n_2484);
  not csa_tree_add_51_79_groupi_g43321(csa_tree_add_51_79_groupi_n_2483 ,csa_tree_add_51_79_groupi_n_2481);
  not csa_tree_add_51_79_groupi_g43326(csa_tree_add_51_79_groupi_n_2478 ,csa_tree_add_51_79_groupi_n_2476);
  not csa_tree_add_51_79_groupi_g43329(csa_tree_add_51_79_groupi_n_2475 ,csa_tree_add_51_79_groupi_n_2473);
  not csa_tree_add_51_79_groupi_g43332(csa_tree_add_51_79_groupi_n_2472 ,csa_tree_add_51_79_groupi_n_2470);
  not csa_tree_add_51_79_groupi_g43335(csa_tree_add_51_79_groupi_n_2469 ,csa_tree_add_51_79_groupi_n_2467);
  not csa_tree_add_51_79_groupi_g43338(csa_tree_add_51_79_groupi_n_2466 ,csa_tree_add_51_79_groupi_n_2464);
  not csa_tree_add_51_79_groupi_g43341(csa_tree_add_51_79_groupi_n_2463 ,csa_tree_add_51_79_groupi_n_2461);
  not csa_tree_add_51_79_groupi_g43344(csa_tree_add_51_79_groupi_n_2460 ,csa_tree_add_51_79_groupi_n_2458);
  not csa_tree_add_51_79_groupi_g43347(csa_tree_add_51_79_groupi_n_2457 ,csa_tree_add_51_79_groupi_n_2455);
  not csa_tree_add_51_79_groupi_g43352(csa_tree_add_51_79_groupi_n_2452 ,csa_tree_add_51_79_groupi_n_2450);
  not csa_tree_add_51_79_groupi_g43355(csa_tree_add_51_79_groupi_n_2449 ,csa_tree_add_51_79_groupi_n_2447);
  not csa_tree_add_51_79_groupi_g43360(csa_tree_add_51_79_groupi_n_2444 ,csa_tree_add_51_79_groupi_n_2442);
  not csa_tree_add_51_79_groupi_g43363(csa_tree_add_51_79_groupi_n_2441 ,csa_tree_add_51_79_groupi_n_2439);
  not csa_tree_add_51_79_groupi_g43366(csa_tree_add_51_79_groupi_n_2438 ,csa_tree_add_51_79_groupi_n_2436);
  and csa_tree_add_51_79_groupi_g43371(csa_tree_add_51_79_groupi_n_2433 ,csa_tree_add_51_79_groupi_n_1126 ,csa_tree_add_51_79_groupi_n_1693);
  nor csa_tree_add_51_79_groupi_g43372(csa_tree_add_51_79_groupi_n_2432 ,in16[1] ,csa_tree_add_51_79_groupi_n_1675);
  and csa_tree_add_51_79_groupi_g43373(csa_tree_add_51_79_groupi_n_2431 ,csa_tree_add_51_79_groupi_n_1138 ,csa_tree_add_51_79_groupi_n_1733);
  and csa_tree_add_51_79_groupi_g43374(csa_tree_add_51_79_groupi_n_2430 ,csa_tree_add_51_79_groupi_n_1144 ,csa_tree_add_51_79_groupi_n_1762);
  and csa_tree_add_51_79_groupi_g43375(csa_tree_add_51_79_groupi_n_2429 ,csa_tree_add_51_79_groupi_n_1077 ,csa_tree_add_51_79_groupi_n_1072);
  and csa_tree_add_51_79_groupi_g43376(csa_tree_add_51_79_groupi_n_2428 ,csa_tree_add_51_79_groupi_n_1534 ,csa_tree_add_51_79_groupi_n_1757);
  and csa_tree_add_51_79_groupi_g43377(csa_tree_add_51_79_groupi_n_2427 ,csa_tree_add_51_79_groupi_n_1536 ,csa_tree_add_51_79_groupi_n_1682);
  and csa_tree_add_51_79_groupi_g43378(csa_tree_add_51_79_groupi_n_2426 ,csa_tree_add_51_79_groupi_n_1549 ,csa_tree_add_51_79_groupi_n_1707);
  and csa_tree_add_51_79_groupi_g43379(csa_tree_add_51_79_groupi_n_2425 ,csa_tree_add_51_79_groupi_n_1605 ,csa_tree_add_51_79_groupi_n_1690);
  and csa_tree_add_51_79_groupi_g43380(csa_tree_add_51_79_groupi_n_2424 ,csa_tree_add_51_79_groupi_n_1616 ,csa_tree_add_51_79_groupi_n_1706);
  and csa_tree_add_51_79_groupi_g43381(csa_tree_add_51_79_groupi_n_2423 ,csa_tree_add_51_79_groupi_n_1531 ,csa_tree_add_51_79_groupi_n_1744);
  xnor csa_tree_add_51_79_groupi_g43382(csa_tree_add_51_79_groupi_n_2422 ,in12[7] ,in12[6]);
  and csa_tree_add_51_79_groupi_g43383(csa_tree_add_51_79_groupi_n_2421 ,csa_tree_add_51_79_groupi_n_1134 ,csa_tree_add_51_79_groupi_n_1708);
  and csa_tree_add_51_79_groupi_g43384(csa_tree_add_51_79_groupi_n_2420 ,csa_tree_add_51_79_groupi_n_1544 ,csa_tree_add_51_79_groupi_n_1709);
  xnor csa_tree_add_51_79_groupi_g43386(csa_tree_add_51_79_groupi_n_2418 ,in14[3] ,in14[2]);
  or csa_tree_add_51_79_groupi_g43387(csa_tree_add_51_79_groupi_n_2417 ,csa_tree_add_51_79_groupi_n_1077 ,csa_tree_add_51_79_groupi_n_1072);
  xnor csa_tree_add_51_79_groupi_g43388(csa_tree_add_51_79_groupi_n_2416 ,in11[0] ,in12[5]);
  and csa_tree_add_51_79_groupi_g43389(csa_tree_add_51_79_groupi_n_2415 ,csa_tree_add_51_79_groupi_n_1073 ,csa_tree_add_51_79_groupi_n_1076);
  and csa_tree_add_51_79_groupi_g43390(csa_tree_add_51_79_groupi_n_2414 ,csa_tree_add_51_79_groupi_n_1146 ,csa_tree_add_51_79_groupi_n_1696);
  and csa_tree_add_51_79_groupi_g43391(csa_tree_add_51_79_groupi_n_2413 ,csa_tree_add_51_79_groupi_n_1618 ,csa_tree_add_51_79_groupi_n_1688);
  and csa_tree_add_51_79_groupi_g43392(csa_tree_add_51_79_groupi_n_2412 ,csa_tree_add_51_79_groupi_n_1615 ,csa_tree_add_51_79_groupi_n_1698);
  and csa_tree_add_51_79_groupi_g43393(csa_tree_add_51_79_groupi_n_2411 ,csa_tree_add_51_79_groupi_n_1140 ,csa_tree_add_51_79_groupi_n_1684);
  and csa_tree_add_51_79_groupi_g43394(csa_tree_add_51_79_groupi_n_2410 ,csa_tree_add_51_79_groupi_n_1551 ,csa_tree_add_51_79_groupi_n_1743);
  and csa_tree_add_51_79_groupi_g43395(csa_tree_add_51_79_groupi_n_2409 ,csa_tree_add_51_79_groupi_n_1128 ,csa_tree_add_51_79_groupi_n_1739);
  and csa_tree_add_51_79_groupi_g43396(csa_tree_add_51_79_groupi_n_2408 ,csa_tree_add_51_79_groupi_n_1620 ,csa_tree_add_51_79_groupi_n_1703);
  nor csa_tree_add_51_79_groupi_g43397(csa_tree_add_51_79_groupi_n_2407 ,in18[1] ,csa_tree_add_51_79_groupi_n_1712);
  and csa_tree_add_51_79_groupi_g43399(csa_tree_add_51_79_groupi_n_2405 ,csa_tree_add_51_79_groupi_n_1538 ,csa_tree_add_51_79_groupi_n_1753);
  and csa_tree_add_51_79_groupi_g43400(csa_tree_add_51_79_groupi_n_2404 ,csa_tree_add_51_79_groupi_n_1132 ,csa_tree_add_51_79_groupi_n_1751);
  xnor csa_tree_add_51_79_groupi_g43401(csa_tree_add_51_79_groupi_n_2403 ,in12[5] ,in12[4]);
  nor csa_tree_add_51_79_groupi_g43402(csa_tree_add_51_79_groupi_n_2402 ,in12[1] ,csa_tree_add_51_79_groupi_n_1764);
  and csa_tree_add_51_79_groupi_g43403(csa_tree_add_51_79_groupi_n_2401 ,csa_tree_add_51_79_groupi_n_1613 ,csa_tree_add_51_79_groupi_n_1716);
  and csa_tree_add_51_79_groupi_g43404(csa_tree_add_51_79_groupi_n_2400 ,csa_tree_add_51_79_groupi_n_1611 ,csa_tree_add_51_79_groupi_n_1745);
  nor csa_tree_add_51_79_groupi_g43406(csa_tree_add_51_79_groupi_n_2398 ,in2[1] ,csa_tree_add_51_79_groupi_n_1728);
  nor csa_tree_add_51_79_groupi_g43407(csa_tree_add_51_79_groupi_n_2397 ,in24[1] ,csa_tree_add_51_79_groupi_n_1718);
  and csa_tree_add_51_79_groupi_g43408(csa_tree_add_51_79_groupi_n_2396 ,csa_tree_add_51_79_groupi_n_1604 ,csa_tree_add_51_79_groupi_n_1736);
  nor csa_tree_add_51_79_groupi_g43409(csa_tree_add_51_79_groupi_n_2395 ,in6[1] ,csa_tree_add_51_79_groupi_n_1756);
  and csa_tree_add_51_79_groupi_g43410(csa_tree_add_51_79_groupi_n_2394 ,csa_tree_add_51_79_groupi_n_1075 ,csa_tree_add_51_79_groupi_n_1074);
  or csa_tree_add_51_79_groupi_g43411(csa_tree_add_51_79_groupi_n_2393 ,csa_tree_add_51_79_groupi_n_1073 ,csa_tree_add_51_79_groupi_n_1076);
  nor csa_tree_add_51_79_groupi_g43412(csa_tree_add_51_79_groupi_n_2392 ,in8[1] ,csa_tree_add_51_79_groupi_n_1741);
  and csa_tree_add_51_79_groupi_g43413(csa_tree_add_51_79_groupi_n_2391 ,csa_tree_add_51_79_groupi_n_1546 ,csa_tree_add_51_79_groupi_n_1769);
  nor csa_tree_add_51_79_groupi_g43414(csa_tree_add_51_79_groupi_n_2390 ,in4[1] ,csa_tree_add_51_79_groupi_n_1702);
  or csa_tree_add_51_79_groupi_g43415(csa_tree_add_51_79_groupi_n_2389 ,csa_tree_add_51_79_groupi_n_1075 ,csa_tree_add_51_79_groupi_n_1074);
  and csa_tree_add_51_79_groupi_g43416(csa_tree_add_51_79_groupi_n_2388 ,csa_tree_add_51_79_groupi_n_1596 ,csa_tree_add_51_79_groupi_n_1749);
  nor csa_tree_add_51_79_groupi_g43417(csa_tree_add_51_79_groupi_n_2387 ,in14[1] ,csa_tree_add_51_79_groupi_n_1748);
  and csa_tree_add_51_79_groupi_g43418(csa_tree_add_51_79_groupi_n_2386 ,csa_tree_add_51_79_groupi_n_1130 ,csa_tree_add_51_79_groupi_n_1740);
  nor csa_tree_add_51_79_groupi_g43419(csa_tree_add_51_79_groupi_n_2385 ,in10[1] ,csa_tree_add_51_79_groupi_n_1765);
  and csa_tree_add_51_79_groupi_g43420(csa_tree_add_51_79_groupi_n_2384 ,csa_tree_add_51_79_groupi_n_1142 ,csa_tree_add_51_79_groupi_n_1711);
  and csa_tree_add_51_79_groupi_g43421(csa_tree_add_51_79_groupi_n_2383 ,csa_tree_add_51_79_groupi_n_1597 ,csa_tree_add_51_79_groupi_n_1726);
  and csa_tree_add_51_79_groupi_g43422(csa_tree_add_51_79_groupi_n_2382 ,csa_tree_add_51_79_groupi_n_1600 ,csa_tree_add_51_79_groupi_n_1761);
  and csa_tree_add_51_79_groupi_g43423(csa_tree_add_51_79_groupi_n_2381 ,csa_tree_add_51_79_groupi_n_1136 ,csa_tree_add_51_79_groupi_n_1686);
  and csa_tree_add_51_79_groupi_g43424(csa_tree_add_51_79_groupi_n_2380 ,csa_tree_add_51_79_groupi_n_1541 ,csa_tree_add_51_79_groupi_n_1713);
  and csa_tree_add_51_79_groupi_g43425(csa_tree_add_51_79_groupi_n_2379 ,csa_tree_add_51_79_groupi_n_1548 ,csa_tree_add_51_79_groupi_n_1771);
  and csa_tree_add_51_79_groupi_g43426(csa_tree_add_51_79_groupi_n_2378 ,csa_tree_add_51_79_groupi_n_1595 ,csa_tree_add_51_79_groupi_n_1734);
  and csa_tree_add_51_79_groupi_g43427(csa_tree_add_51_79_groupi_n_2377 ,csa_tree_add_51_79_groupi_n_1598 ,csa_tree_add_51_79_groupi_n_1695);
  and csa_tree_add_51_79_groupi_g43428(csa_tree_add_51_79_groupi_n_2376 ,csa_tree_add_51_79_groupi_n_1619 ,csa_tree_add_51_79_groupi_n_1685);
  and csa_tree_add_51_79_groupi_g43429(csa_tree_add_51_79_groupi_n_2375 ,csa_tree_add_51_79_groupi_n_1608 ,csa_tree_add_51_79_groupi_n_1763);
  nor csa_tree_add_51_79_groupi_g43430(csa_tree_add_51_79_groupi_n_2374 ,in22[1] ,csa_tree_add_51_79_groupi_n_1773);
  nor csa_tree_add_51_79_groupi_g43431(csa_tree_add_51_79_groupi_n_2373 ,in20[1] ,csa_tree_add_51_79_groupi_n_1760);
  xnor csa_tree_add_51_79_groupi_g43432(csa_tree_add_51_79_groupi_n_2372 ,in2[3] ,in2[2]);
  xnor csa_tree_add_51_79_groupi_g43433(csa_tree_add_51_79_groupi_n_2371 ,in23[0] ,in24[1]);
  xnor csa_tree_add_51_79_groupi_g43434(csa_tree_add_51_79_groupi_n_2370 ,in7[0] ,in8[7]);
  xnor csa_tree_add_51_79_groupi_g43435(csa_tree_add_51_79_groupi_n_2369 ,in21[0] ,in22[5]);
  xnor csa_tree_add_51_79_groupi_g43436(csa_tree_add_51_79_groupi_n_2368 ,in21[0] ,in22[7]);
  xnor csa_tree_add_51_79_groupi_g43437(csa_tree_add_51_79_groupi_n_2367 ,in19[0] ,in20[3]);
  xnor csa_tree_add_51_79_groupi_g43438(csa_tree_add_51_79_groupi_n_2366 ,in5[0] ,in6[5]);
  xnor csa_tree_add_51_79_groupi_g43439(csa_tree_add_51_79_groupi_n_2365 ,in4[7] ,in4[6]);
  xnor csa_tree_add_51_79_groupi_g43440(csa_tree_add_51_79_groupi_n_2364 ,in16[3] ,in16[2]);
  xnor csa_tree_add_51_79_groupi_g43441(csa_tree_add_51_79_groupi_n_2363 ,in20[7] ,in20[6]);
  xnor csa_tree_add_51_79_groupi_g43442(csa_tree_add_51_79_groupi_n_2362 ,in24[3] ,in24[2]);
  xnor csa_tree_add_51_79_groupi_g43444(csa_tree_add_51_79_groupi_n_2360 ,in2[7] ,in2[6]);
  xnor csa_tree_add_51_79_groupi_g43445(csa_tree_add_51_79_groupi_n_2359 ,in5[0] ,in6[7]);
  xnor csa_tree_add_51_79_groupi_g43446(csa_tree_add_51_79_groupi_n_2358 ,in13[0] ,in14[7]);
  xnor csa_tree_add_51_79_groupi_g43448(csa_tree_add_51_79_groupi_n_2356 ,in1[0] ,in2[5]);
  xnor csa_tree_add_51_79_groupi_g43449(csa_tree_add_51_79_groupi_n_2355 ,in17[0] ,in18[3]);
  xnor csa_tree_add_51_79_groupi_g43450(csa_tree_add_51_79_groupi_n_2354 ,in6[7] ,in6[6]);
  xnor csa_tree_add_51_79_groupi_g43451(csa_tree_add_51_79_groupi_n_2353 ,in23[0] ,in24[7]);
  xnor csa_tree_add_51_79_groupi_g43452(csa_tree_add_51_79_groupi_n_2352 ,in11[0] ,in12[3]);
  xnor csa_tree_add_51_79_groupi_g43454(csa_tree_add_51_79_groupi_n_2350 ,in15[0] ,in16[7]);
  xnor csa_tree_add_51_79_groupi_g43455(csa_tree_add_51_79_groupi_n_2349 ,in4[3] ,in4[2]);
  xnor csa_tree_add_51_79_groupi_g43456(csa_tree_add_51_79_groupi_n_2348 ,in3[0] ,in4[7]);
  xnor csa_tree_add_51_79_groupi_g43457(csa_tree_add_51_79_groupi_n_2347 ,in6[5] ,in6[4]);
  xnor csa_tree_add_51_79_groupi_g43458(csa_tree_add_51_79_groupi_n_2346 ,in5[0] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g43459(csa_tree_add_51_79_groupi_n_2345 ,in22[3] ,in22[2]);
  xnor csa_tree_add_51_79_groupi_g43462(csa_tree_add_51_79_groupi_n_2342 ,in10[7] ,in10[6]);
  xnor csa_tree_add_51_79_groupi_g43464(csa_tree_add_51_79_groupi_n_2340 ,in17[0] ,in18[5]);
  xnor csa_tree_add_51_79_groupi_g43465(csa_tree_add_51_79_groupi_n_2339 ,in12[3] ,in12[2]);
  xnor csa_tree_add_51_79_groupi_g43466(csa_tree_add_51_79_groupi_n_2338 ,in18[5] ,in18[4]);
  xnor csa_tree_add_51_79_groupi_g43468(csa_tree_add_51_79_groupi_n_2336 ,in17[0] ,in18[1]);
  xnor csa_tree_add_51_79_groupi_g43469(csa_tree_add_51_79_groupi_n_2335 ,in1[0] ,in2[7]);
  xnor csa_tree_add_51_79_groupi_g43470(csa_tree_add_51_79_groupi_n_2334 ,in15[0] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g43471(csa_tree_add_51_79_groupi_n_2333 ,in14[7] ,in14[6]);
  xnor csa_tree_add_51_79_groupi_g43472(csa_tree_add_51_79_groupi_n_2332 ,in18[7] ,in18[6]);
  xnor csa_tree_add_51_79_groupi_g43473(csa_tree_add_51_79_groupi_n_2331 ,in24[5] ,in24[4]);
  xnor csa_tree_add_51_79_groupi_g43475(csa_tree_add_51_79_groupi_n_2329 ,in22[7] ,in22[6]);
  xnor csa_tree_add_51_79_groupi_g43476(csa_tree_add_51_79_groupi_n_2328 ,in9[0] ,in10[3]);
  xnor csa_tree_add_51_79_groupi_g43477(csa_tree_add_51_79_groupi_n_2327 ,in23[0] ,in24[5]);
  xnor csa_tree_add_51_79_groupi_g43479(csa_tree_add_51_79_groupi_n_2325 ,in9[0] ,in10[5]);
  xnor csa_tree_add_51_79_groupi_g43480(csa_tree_add_51_79_groupi_n_2324 ,in3[0] ,in4[3]);
  xnor csa_tree_add_51_79_groupi_g43481(csa_tree_add_51_79_groupi_n_2323 ,in20[5] ,in20[4]);
  xnor csa_tree_add_51_79_groupi_g43483(csa_tree_add_51_79_groupi_n_2321 ,in24[7] ,in24[6]);
  xnor csa_tree_add_51_79_groupi_g43484(csa_tree_add_51_79_groupi_n_2320 ,in13[0] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g43485(csa_tree_add_51_79_groupi_n_2884 ,in1[10] ,in2[7]);
  xnor csa_tree_add_51_79_groupi_g43486(csa_tree_add_51_79_groupi_n_2883 ,in11[8] ,in12[1]);
  xnor csa_tree_add_51_79_groupi_g43487(csa_tree_add_51_79_groupi_n_2882 ,in1[10] ,in2[3]);
  xnor csa_tree_add_51_79_groupi_g43488(csa_tree_add_51_79_groupi_n_2881 ,in15[3] ,in16[7]);
  xnor csa_tree_add_51_79_groupi_g43489(csa_tree_add_51_79_groupi_n_2880 ,in17[7] ,in18[1]);
  xnor csa_tree_add_51_79_groupi_g43490(csa_tree_add_51_79_groupi_n_2879 ,in3[1] ,in4[3]);
  xnor csa_tree_add_51_79_groupi_g43491(csa_tree_add_51_79_groupi_n_2878 ,in11[3] ,in12[5]);
  xnor csa_tree_add_51_79_groupi_g43492(csa_tree_add_51_79_groupi_n_2877 ,in21[7] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g43493(csa_tree_add_51_79_groupi_n_2876 ,in21[1] ,in22[7]);
  xnor csa_tree_add_51_79_groupi_g43494(csa_tree_add_51_79_groupi_n_2875 ,in3[6] ,in4[1]);
  xnor csa_tree_add_51_79_groupi_g43495(csa_tree_add_51_79_groupi_n_2874 ,in11[7] ,in12[7]);
  xnor csa_tree_add_51_79_groupi_g43496(csa_tree_add_51_79_groupi_n_2873 ,in17[1] ,in18[5]);
  xnor csa_tree_add_51_79_groupi_g43497(csa_tree_add_51_79_groupi_n_2872 ,in19[3] ,in20[5]);
  xnor csa_tree_add_51_79_groupi_g43498(csa_tree_add_51_79_groupi_n_2871 ,in19[5] ,in20[3]);
  xnor csa_tree_add_51_79_groupi_g43499(csa_tree_add_51_79_groupi_n_2870 ,in17[4] ,in18[1]);
  xnor csa_tree_add_51_79_groupi_g43500(csa_tree_add_51_79_groupi_n_2869 ,in23[9] ,in24[7]);
  xnor csa_tree_add_51_79_groupi_g43501(csa_tree_add_51_79_groupi_n_2868 ,in1[5] ,in2[7]);
  xnor csa_tree_add_51_79_groupi_g43502(csa_tree_add_51_79_groupi_n_2867 ,in1[7] ,in2[5]);
  xnor csa_tree_add_51_79_groupi_g43503(csa_tree_add_51_79_groupi_n_2866 ,in1[9] ,in2[1]);
  xnor csa_tree_add_51_79_groupi_g43504(csa_tree_add_51_79_groupi_n_2865 ,in15[4] ,in16[7]);
  xnor csa_tree_add_51_79_groupi_g43505(csa_tree_add_51_79_groupi_n_2864 ,in19[5] ,in20[5]);
  xnor csa_tree_add_51_79_groupi_g43506(csa_tree_add_51_79_groupi_n_2863 ,in13[3] ,in14[7]);
  xnor csa_tree_add_51_79_groupi_g43507(csa_tree_add_51_79_groupi_n_2862 ,in21[2] ,in22[7]);
  xnor csa_tree_add_51_79_groupi_g43508(csa_tree_add_51_79_groupi_n_2861 ,in17[5] ,in18[3]);
  xnor csa_tree_add_51_79_groupi_g43509(csa_tree_add_51_79_groupi_n_2860 ,in13[5] ,in14[7]);
  xnor csa_tree_add_51_79_groupi_g43510(csa_tree_add_51_79_groupi_n_2859 ,in23[6] ,in24[5]);
  xnor csa_tree_add_51_79_groupi_g43511(csa_tree_add_51_79_groupi_n_2858 ,in19[10] ,in20[1]);
  xnor csa_tree_add_51_79_groupi_g43512(csa_tree_add_51_79_groupi_n_2857 ,in3[4] ,in4[3]);
  xnor csa_tree_add_51_79_groupi_g43513(csa_tree_add_51_79_groupi_n_2856 ,in17[4] ,in18[7]);
  xnor csa_tree_add_51_79_groupi_g43514(csa_tree_add_51_79_groupi_n_2855 ,in11[2] ,in12[3]);
  xnor csa_tree_add_51_79_groupi_g43515(csa_tree_add_51_79_groupi_n_2854 ,in23[8] ,in24[7]);
  xnor csa_tree_add_51_79_groupi_g43516(csa_tree_add_51_79_groupi_n_2853 ,in21[4] ,in22[5]);
  xnor csa_tree_add_51_79_groupi_g43517(csa_tree_add_51_79_groupi_n_2852 ,in3[3] ,in4[1]);
  xnor csa_tree_add_51_79_groupi_g43518(csa_tree_add_51_79_groupi_n_2851 ,in13[2] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g43519(csa_tree_add_51_79_groupi_n_2850 ,in9[8] ,in10[5]);
  xnor csa_tree_add_51_79_groupi_g43520(csa_tree_add_51_79_groupi_n_2849 ,in21[7] ,in22[7]);
  xnor csa_tree_add_51_79_groupi_g43521(csa_tree_add_51_79_groupi_n_2848 ,in5[7] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g43522(csa_tree_add_51_79_groupi_n_2847 ,in13[3] ,in14[3]);
  xnor csa_tree_add_51_79_groupi_g43523(csa_tree_add_51_79_groupi_n_2846 ,in9[5] ,in10[7]);
  xnor csa_tree_add_51_79_groupi_g43524(csa_tree_add_51_79_groupi_n_2845 ,in15[3] ,in16[5]);
  xnor csa_tree_add_51_79_groupi_g43525(csa_tree_add_51_79_groupi_n_2844 ,in15[1] ,in16[7]);
  xnor csa_tree_add_51_79_groupi_g43526(csa_tree_add_51_79_groupi_n_2843 ,in21[3] ,in22[7]);
  xnor csa_tree_add_51_79_groupi_g43527(csa_tree_add_51_79_groupi_n_2842 ,in9[9] ,in10[3]);
  xnor csa_tree_add_51_79_groupi_g43528(csa_tree_add_51_79_groupi_n_2841 ,in5[6] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g43529(csa_tree_add_51_79_groupi_n_2840 ,in7[5] ,in8[3]);
  xnor csa_tree_add_51_79_groupi_g43530(csa_tree_add_51_79_groupi_n_2839 ,in7[3] ,in8[5]);
  xnor csa_tree_add_51_79_groupi_g43531(csa_tree_add_51_79_groupi_n_2838 ,in13[6] ,in14[5]);
  xnor csa_tree_add_51_79_groupi_g43532(csa_tree_add_51_79_groupi_n_2837 ,in23[3] ,in24[5]);
  xnor csa_tree_add_51_79_groupi_g43533(csa_tree_add_51_79_groupi_n_2836 ,in21[9] ,in22[3]);
  xnor csa_tree_add_51_79_groupi_g43534(csa_tree_add_51_79_groupi_n_2835 ,in23[4] ,in24[7]);
  xnor csa_tree_add_51_79_groupi_g43535(csa_tree_add_51_79_groupi_n_2834 ,in21[7] ,in22[3]);
  xnor csa_tree_add_51_79_groupi_g43536(csa_tree_add_51_79_groupi_n_2833 ,in21[5] ,in22[3]);
  xnor csa_tree_add_51_79_groupi_g43537(csa_tree_add_51_79_groupi_n_2832 ,in13[5] ,in14[3]);
  xnor csa_tree_add_51_79_groupi_g43538(csa_tree_add_51_79_groupi_n_2831 ,in9[5] ,in10[1]);
  xnor csa_tree_add_51_79_groupi_g43539(csa_tree_add_51_79_groupi_n_2830 ,in11[5] ,in12[1]);
  xnor csa_tree_add_51_79_groupi_g43540(csa_tree_add_51_79_groupi_n_2829 ,in7[8] ,in8[7]);
  xnor csa_tree_add_51_79_groupi_g43541(csa_tree_add_51_79_groupi_n_2828 ,in17[3] ,in18[5]);
  xnor csa_tree_add_51_79_groupi_g43542(csa_tree_add_51_79_groupi_n_2827 ,in11[1] ,in12[3]);
  xnor csa_tree_add_51_79_groupi_g43543(csa_tree_add_51_79_groupi_n_2826 ,in21[1] ,in22[3]);
  xnor csa_tree_add_51_79_groupi_g43544(csa_tree_add_51_79_groupi_n_2825 ,in13[4] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g43545(csa_tree_add_51_79_groupi_n_2824 ,in19[7] ,in20[1]);
  xnor csa_tree_add_51_79_groupi_g43546(csa_tree_add_51_79_groupi_n_2823 ,in21[7] ,in22[5]);
  xnor csa_tree_add_51_79_groupi_g43547(csa_tree_add_51_79_groupi_n_2822 ,in11[5] ,in12[7]);
  xnor csa_tree_add_51_79_groupi_g43548(csa_tree_add_51_79_groupi_n_2821 ,in15[9] ,in16[7]);
  xnor csa_tree_add_51_79_groupi_g43549(csa_tree_add_51_79_groupi_n_2820 ,in21[5] ,in22[7]);
  xnor csa_tree_add_51_79_groupi_g43550(csa_tree_add_51_79_groupi_n_2819 ,in23[5] ,in24[3]);
  xnor csa_tree_add_51_79_groupi_g43551(csa_tree_add_51_79_groupi_n_2818 ,in21[5] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g43552(csa_tree_add_51_79_groupi_n_2817 ,in3[5] ,in4[5]);
  xnor csa_tree_add_51_79_groupi_g43553(csa_tree_add_51_79_groupi_n_2816 ,in9[1] ,in10[7]);
  xnor csa_tree_add_51_79_groupi_g43554(csa_tree_add_51_79_groupi_n_2815 ,in13[6] ,in14[7]);
  xnor csa_tree_add_51_79_groupi_g43555(csa_tree_add_51_79_groupi_n_2814 ,in13[9] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g43556(csa_tree_add_51_79_groupi_n_2813 ,in21[8] ,in22[7]);
  xnor csa_tree_add_51_79_groupi_g43557(csa_tree_add_51_79_groupi_n_2812 ,in9[2] ,in10[1]);
  xnor csa_tree_add_51_79_groupi_g43558(csa_tree_add_51_79_groupi_n_2811 ,in23[7] ,in24[3]);
  xnor csa_tree_add_51_79_groupi_g43559(csa_tree_add_51_79_groupi_n_2810 ,in19[4] ,in20[1]);
  xnor csa_tree_add_51_79_groupi_g43560(csa_tree_add_51_79_groupi_n_2809 ,in11[5] ,in12[5]);
  xnor csa_tree_add_51_79_groupi_g43561(csa_tree_add_51_79_groupi_n_2808 ,in1[4] ,in2[3]);
  xnor csa_tree_add_51_79_groupi_g43562(csa_tree_add_51_79_groupi_n_2807 ,in19[8] ,in20[1]);
  xnor csa_tree_add_51_79_groupi_g43563(csa_tree_add_51_79_groupi_n_2806 ,in7[7] ,in8[3]);
  xnor csa_tree_add_51_79_groupi_g43564(csa_tree_add_51_79_groupi_n_2805 ,in9[6] ,in10[5]);
  xnor csa_tree_add_51_79_groupi_g43565(csa_tree_add_51_79_groupi_n_2804 ,in11[6] ,in12[3]);
  xnor csa_tree_add_51_79_groupi_g43566(csa_tree_add_51_79_groupi_n_2803 ,in1[5] ,in2[1]);
  xnor csa_tree_add_51_79_groupi_g43567(csa_tree_add_51_79_groupi_n_2802 ,in11[5] ,in12[3]);
  xnor csa_tree_add_51_79_groupi_g43568(csa_tree_add_51_79_groupi_n_2801 ,in15[8] ,in16[7]);
  xnor csa_tree_add_51_79_groupi_g43569(csa_tree_add_51_79_groupi_n_2800 ,in13[4] ,in14[3]);
  xnor csa_tree_add_51_79_groupi_g43570(csa_tree_add_51_79_groupi_n_2799 ,in23[6] ,in24[1]);
  xnor csa_tree_add_51_79_groupi_g43571(csa_tree_add_51_79_groupi_n_2798 ,in3[8] ,in4[5]);
  xnor csa_tree_add_51_79_groupi_g43572(csa_tree_add_51_79_groupi_n_2797 ,in7[9] ,in8[5]);
  xnor csa_tree_add_51_79_groupi_g43573(csa_tree_add_51_79_groupi_n_2796 ,in17[5] ,in18[7]);
  xnor csa_tree_add_51_79_groupi_g43574(csa_tree_add_51_79_groupi_n_2794 ,csa_tree_add_51_79_groupi_n_1136 ,in11[10]);
  xnor csa_tree_add_51_79_groupi_g43575(csa_tree_add_51_79_groupi_n_2793 ,in21[9] ,in22[5]);
  xnor csa_tree_add_51_79_groupi_g43576(csa_tree_add_51_79_groupi_n_2792 ,in5[4] ,in6[7]);
  xnor csa_tree_add_51_79_groupi_g43577(csa_tree_add_51_79_groupi_n_2791 ,in5[5] ,in6[5]);
  xnor csa_tree_add_51_79_groupi_g43578(csa_tree_add_51_79_groupi_n_2790 ,in21[10] ,in22[7]);
  xnor csa_tree_add_51_79_groupi_g43579(csa_tree_add_51_79_groupi_n_2789 ,in19[9] ,in20[7]);
  xnor csa_tree_add_51_79_groupi_g43580(csa_tree_add_51_79_groupi_n_2788 ,in23[7] ,in24[7]);
  xnor csa_tree_add_51_79_groupi_g43581(csa_tree_add_51_79_groupi_n_2787 ,in17[1] ,in18[3]);
  xnor csa_tree_add_51_79_groupi_g43582(csa_tree_add_51_79_groupi_n_2786 ,in15[4] ,in16[3]);
  xnor csa_tree_add_51_79_groupi_g43583(csa_tree_add_51_79_groupi_n_2785 ,in5[4] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g43584(csa_tree_add_51_79_groupi_n_2784 ,in3[8] ,in4[1]);
  xnor csa_tree_add_51_79_groupi_g43585(csa_tree_add_51_79_groupi_n_2783 ,in5[5] ,in6[7]);
  xnor csa_tree_add_51_79_groupi_g43586(csa_tree_add_51_79_groupi_n_2782 ,in1[4] ,in2[5]);
  xnor csa_tree_add_51_79_groupi_g43587(csa_tree_add_51_79_groupi_n_2781 ,in5[8] ,in6[3]);
  xnor csa_tree_add_51_79_groupi_g43588(csa_tree_add_51_79_groupi_n_2780 ,in9[3] ,in10[7]);
  xnor csa_tree_add_51_79_groupi_g43589(csa_tree_add_51_79_groupi_n_2779 ,in19[4] ,in20[5]);
  xnor csa_tree_add_51_79_groupi_g43590(csa_tree_add_51_79_groupi_n_2778 ,in9[6] ,in10[7]);
  xnor csa_tree_add_51_79_groupi_g43591(csa_tree_add_51_79_groupi_n_2777 ,in5[1] ,in6[5]);
  xnor csa_tree_add_51_79_groupi_g43592(csa_tree_add_51_79_groupi_n_2776 ,in15[5] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g43593(csa_tree_add_51_79_groupi_n_2775 ,in5[7] ,in6[7]);
  xnor csa_tree_add_51_79_groupi_g43594(csa_tree_add_51_79_groupi_n_2774 ,in5[9] ,in6[7]);
  xnor csa_tree_add_51_79_groupi_g43595(csa_tree_add_51_79_groupi_n_2772 ,csa_tree_add_51_79_groupi_n_1138 ,in23[10]);
  xnor csa_tree_add_51_79_groupi_g43596(csa_tree_add_51_79_groupi_n_2771 ,in17[6] ,in18[1]);
  xnor csa_tree_add_51_79_groupi_g43597(csa_tree_add_51_79_groupi_n_2770 ,in13[5] ,in14[5]);
  xnor csa_tree_add_51_79_groupi_g43598(csa_tree_add_51_79_groupi_n_2769 ,in11[4] ,in12[3]);
  xnor csa_tree_add_51_79_groupi_g43599(csa_tree_add_51_79_groupi_n_2768 ,in5[3] ,in6[5]);
  xnor csa_tree_add_51_79_groupi_g43600(csa_tree_add_51_79_groupi_n_2767 ,in9[6] ,in10[1]);
  xnor csa_tree_add_51_79_groupi_g43601(csa_tree_add_51_79_groupi_n_2766 ,in17[2] ,in18[5]);
  xnor csa_tree_add_51_79_groupi_g43602(csa_tree_add_51_79_groupi_n_2765 ,in5[7] ,in6[5]);
  xnor csa_tree_add_51_79_groupi_g43603(csa_tree_add_51_79_groupi_n_2764 ,in21[2] ,in22[5]);
  xnor csa_tree_add_51_79_groupi_g43604(csa_tree_add_51_79_groupi_n_2763 ,in19[8] ,in20[5]);
  xnor csa_tree_add_51_79_groupi_g43605(csa_tree_add_51_79_groupi_n_2762 ,in17[10] ,in18[7]);
  xnor csa_tree_add_51_79_groupi_g43606(csa_tree_add_51_79_groupi_n_2761 ,in3[9] ,in4[3]);
  xnor csa_tree_add_51_79_groupi_g43607(csa_tree_add_51_79_groupi_n_2760 ,in5[2] ,in6[3]);
  xnor csa_tree_add_51_79_groupi_g43608(csa_tree_add_51_79_groupi_n_2759 ,in1[10] ,in2[1]);
  xnor csa_tree_add_51_79_groupi_g43609(csa_tree_add_51_79_groupi_n_2758 ,in1[6] ,in2[1]);
  xnor csa_tree_add_51_79_groupi_g43610(csa_tree_add_51_79_groupi_n_2757 ,in5[10] ,in6[7]);
  xnor csa_tree_add_51_79_groupi_g43611(csa_tree_add_51_79_groupi_n_2756 ,in9[8] ,in10[7]);
  xnor csa_tree_add_51_79_groupi_g43612(csa_tree_add_51_79_groupi_n_2755 ,in23[2] ,in24[5]);
  xnor csa_tree_add_51_79_groupi_g43613(csa_tree_add_51_79_groupi_n_2754 ,in15[5] ,in16[7]);
  xnor csa_tree_add_51_79_groupi_g43614(csa_tree_add_51_79_groupi_n_2753 ,in3[5] ,in4[3]);
  xnor csa_tree_add_51_79_groupi_g43615(csa_tree_add_51_79_groupi_n_2752 ,in7[7] ,in8[5]);
  xnor csa_tree_add_51_79_groupi_g43616(csa_tree_add_51_79_groupi_n_2751 ,in7[9] ,in8[7]);
  xnor csa_tree_add_51_79_groupi_g43617(csa_tree_add_51_79_groupi_n_2750 ,in13[2] ,in14[5]);
  xnor csa_tree_add_51_79_groupi_g43618(csa_tree_add_51_79_groupi_n_2749 ,in17[4] ,in18[5]);
  xnor csa_tree_add_51_79_groupi_g43619(csa_tree_add_51_79_groupi_n_2748 ,in21[6] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g43620(csa_tree_add_51_79_groupi_n_2747 ,in23[3] ,in24[7]);
  xnor csa_tree_add_51_79_groupi_g43621(csa_tree_add_51_79_groupi_n_2746 ,in13[1] ,in14[3]);
  xnor csa_tree_add_51_79_groupi_g43622(csa_tree_add_51_79_groupi_n_2745 ,in23[2] ,in24[1]);
  xnor csa_tree_add_51_79_groupi_g43623(csa_tree_add_51_79_groupi_n_2744 ,in17[8] ,in18[5]);
  xnor csa_tree_add_51_79_groupi_g43624(csa_tree_add_51_79_groupi_n_2743 ,in21[9] ,in22[7]);
  xnor csa_tree_add_51_79_groupi_g43625(csa_tree_add_51_79_groupi_n_2742 ,in7[5] ,in8[7]);
  xnor csa_tree_add_51_79_groupi_g43626(csa_tree_add_51_79_groupi_n_2741 ,in19[2] ,in20[3]);
  xnor csa_tree_add_51_79_groupi_g43627(csa_tree_add_51_79_groupi_n_2740 ,in17[7] ,in18[3]);
  xnor csa_tree_add_51_79_groupi_g43628(csa_tree_add_51_79_groupi_n_2739 ,in17[6] ,in18[5]);
  xnor csa_tree_add_51_79_groupi_g43629(csa_tree_add_51_79_groupi_n_2738 ,in3[6] ,in4[7]);
  xnor csa_tree_add_51_79_groupi_g43630(csa_tree_add_51_79_groupi_n_2737 ,in1[2] ,in2[3]);
  xnor csa_tree_add_51_79_groupi_g43631(csa_tree_add_51_79_groupi_n_2736 ,in15[6] ,in16[7]);
  xnor csa_tree_add_51_79_groupi_g43632(csa_tree_add_51_79_groupi_n_2735 ,in13[6] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g43633(csa_tree_add_51_79_groupi_n_2734 ,in19[6] ,in20[1]);
  xnor csa_tree_add_51_79_groupi_g43634(csa_tree_add_51_79_groupi_n_2733 ,in3[2] ,in4[7]);
  xnor csa_tree_add_51_79_groupi_g43635(csa_tree_add_51_79_groupi_n_2732 ,in5[5] ,in6[3]);
  xnor csa_tree_add_51_79_groupi_g43636(csa_tree_add_51_79_groupi_n_2731 ,in1[6] ,in2[5]);
  xnor csa_tree_add_51_79_groupi_g43637(csa_tree_add_51_79_groupi_n_2730 ,in7[7] ,in8[7]);
  xnor csa_tree_add_51_79_groupi_g43638(csa_tree_add_51_79_groupi_n_2729 ,in1[3] ,in2[5]);
  xnor csa_tree_add_51_79_groupi_g43639(csa_tree_add_51_79_groupi_n_2728 ,in9[2] ,in10[3]);
  xnor csa_tree_add_51_79_groupi_g43640(csa_tree_add_51_79_groupi_n_2727 ,in21[3] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g43641(csa_tree_add_51_79_groupi_n_2726 ,in1[5] ,in2[5]);
  xnor csa_tree_add_51_79_groupi_g43642(csa_tree_add_51_79_groupi_n_2725 ,in11[9] ,in12[3]);
  xnor csa_tree_add_51_79_groupi_g43643(csa_tree_add_51_79_groupi_n_2724 ,in21[4] ,in22[3]);
  xnor csa_tree_add_51_79_groupi_g43644(csa_tree_add_51_79_groupi_n_2723 ,in15[9] ,in16[5]);
  xnor csa_tree_add_51_79_groupi_g43645(csa_tree_add_51_79_groupi_n_2722 ,in5[4] ,in6[3]);
  xnor csa_tree_add_51_79_groupi_g43646(csa_tree_add_51_79_groupi_n_2721 ,in1[8] ,in2[5]);
  xnor csa_tree_add_51_79_groupi_g43647(csa_tree_add_51_79_groupi_n_2720 ,in11[1] ,in12[7]);
  xnor csa_tree_add_51_79_groupi_g43648(csa_tree_add_51_79_groupi_n_2719 ,in23[1] ,in24[3]);
  xnor csa_tree_add_51_79_groupi_g43649(csa_tree_add_51_79_groupi_n_2718 ,in23[8] ,in24[5]);
  xnor csa_tree_add_51_79_groupi_g43650(csa_tree_add_51_79_groupi_n_2717 ,in17[5] ,in18[5]);
  xnor csa_tree_add_51_79_groupi_g43651(csa_tree_add_51_79_groupi_n_2716 ,in21[6] ,in22[7]);
  xnor csa_tree_add_51_79_groupi_g43652(csa_tree_add_51_79_groupi_n_2715 ,in5[8] ,in6[7]);
  xnor csa_tree_add_51_79_groupi_g43653(csa_tree_add_51_79_groupi_n_2714 ,in19[9] ,in20[3]);
  xnor csa_tree_add_51_79_groupi_g43654(csa_tree_add_51_79_groupi_n_2713 ,in23[9] ,in24[1]);
  xnor csa_tree_add_51_79_groupi_g43655(csa_tree_add_51_79_groupi_n_2712 ,in7[5] ,in8[5]);
  xnor csa_tree_add_51_79_groupi_g43656(csa_tree_add_51_79_groupi_n_2711 ,in21[8] ,in22[5]);
  xnor csa_tree_add_51_79_groupi_g43657(csa_tree_add_51_79_groupi_n_2710 ,in19[4] ,in20[3]);
  xnor csa_tree_add_51_79_groupi_g43658(csa_tree_add_51_79_groupi_n_2709 ,in3[7] ,in4[3]);
  xnor csa_tree_add_51_79_groupi_g43659(csa_tree_add_51_79_groupi_n_2708 ,in5[2] ,in6[5]);
  xnor csa_tree_add_51_79_groupi_g43660(csa_tree_add_51_79_groupi_n_2707 ,in7[6] ,in8[7]);
  xnor csa_tree_add_51_79_groupi_g43661(csa_tree_add_51_79_groupi_n_2706 ,in15[10] ,in16[5]);
  xnor csa_tree_add_51_79_groupi_g43662(csa_tree_add_51_79_groupi_n_2705 ,in19[2] ,in20[5]);
  xnor csa_tree_add_51_79_groupi_g43663(csa_tree_add_51_79_groupi_n_2704 ,in3[7] ,in4[5]);
  xnor csa_tree_add_51_79_groupi_g43664(csa_tree_add_51_79_groupi_n_2703 ,in13[10] ,in14[5]);
  xnor csa_tree_add_51_79_groupi_g43665(csa_tree_add_51_79_groupi_n_2702 ,in17[6] ,in18[3]);
  xnor csa_tree_add_51_79_groupi_g43666(csa_tree_add_51_79_groupi_n_2701 ,in13[8] ,in14[5]);
  xnor csa_tree_add_51_79_groupi_g43667(csa_tree_add_51_79_groupi_n_2700 ,in5[1] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g43668(csa_tree_add_51_79_groupi_n_2699 ,in19[3] ,in20[7]);
  xnor csa_tree_add_51_79_groupi_g43669(csa_tree_add_51_79_groupi_n_2698 ,in21[10] ,in22[3]);
  xnor csa_tree_add_51_79_groupi_g43670(csa_tree_add_51_79_groupi_n_2697 ,in19[7] ,in20[3]);
  xnor csa_tree_add_51_79_groupi_g43671(csa_tree_add_51_79_groupi_n_2696 ,in17[2] ,in18[1]);
  xnor csa_tree_add_51_79_groupi_g43672(csa_tree_add_51_79_groupi_n_2695 ,in23[3] ,in24[1]);
  xnor csa_tree_add_51_79_groupi_g43673(csa_tree_add_51_79_groupi_n_2694 ,in9[7] ,in10[7]);
  xnor csa_tree_add_51_79_groupi_g43674(csa_tree_add_51_79_groupi_n_2693 ,in3[10] ,in4[7]);
  xnor csa_tree_add_51_79_groupi_g43675(csa_tree_add_51_79_groupi_n_2692 ,in19[8] ,in20[3]);
  xnor csa_tree_add_51_79_groupi_g43676(csa_tree_add_51_79_groupi_n_2691 ,in15[8] ,in16[5]);
  xnor csa_tree_add_51_79_groupi_g43677(csa_tree_add_51_79_groupi_n_2690 ,in13[3] ,in14[5]);
  xnor csa_tree_add_51_79_groupi_g43678(csa_tree_add_51_79_groupi_n_2689 ,in5[3] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g43679(csa_tree_add_51_79_groupi_n_2688 ,in1[2] ,in2[1]);
  xnor csa_tree_add_51_79_groupi_g43680(csa_tree_add_51_79_groupi_n_2687 ,in19[3] ,in20[3]);
  xnor csa_tree_add_51_79_groupi_g43681(csa_tree_add_51_79_groupi_n_2686 ,in9[7] ,in10[1]);
  xnor csa_tree_add_51_79_groupi_g43682(csa_tree_add_51_79_groupi_n_2685 ,in15[1] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g43683(csa_tree_add_51_79_groupi_n_2684 ,in7[1] ,in8[3]);
  xnor csa_tree_add_51_79_groupi_g43684(csa_tree_add_51_79_groupi_n_2683 ,in11[7] ,in12[1]);
  xnor csa_tree_add_51_79_groupi_g43685(csa_tree_add_51_79_groupi_n_2682 ,in3[9] ,in4[7]);
  xnor csa_tree_add_51_79_groupi_g43686(csa_tree_add_51_79_groupi_n_2681 ,in1[8] ,in2[7]);
  xnor csa_tree_add_51_79_groupi_g43687(csa_tree_add_51_79_groupi_n_2680 ,in17[2] ,in18[3]);
  xnor csa_tree_add_51_79_groupi_g43688(csa_tree_add_51_79_groupi_n_2679 ,in9[5] ,in10[5]);
  xnor csa_tree_add_51_79_groupi_g43689(csa_tree_add_51_79_groupi_n_2678 ,in1[7] ,in2[3]);
  xnor csa_tree_add_51_79_groupi_g43690(csa_tree_add_51_79_groupi_n_2677 ,in7[5] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g43691(csa_tree_add_51_79_groupi_n_2676 ,in13[5] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g43692(csa_tree_add_51_79_groupi_n_2675 ,in5[9] ,in6[3]);
  xnor csa_tree_add_51_79_groupi_g43693(csa_tree_add_51_79_groupi_n_2674 ,in11[8] ,in12[3]);
  xnor csa_tree_add_51_79_groupi_g43694(csa_tree_add_51_79_groupi_n_2673 ,in3[3] ,in4[3]);
  xnor csa_tree_add_51_79_groupi_g43695(csa_tree_add_51_79_groupi_n_2672 ,in11[6] ,in12[5]);
  xnor csa_tree_add_51_79_groupi_g43696(csa_tree_add_51_79_groupi_n_2671 ,in17[10] ,in18[1]);
  xnor csa_tree_add_51_79_groupi_g43697(csa_tree_add_51_79_groupi_n_2670 ,in13[1] ,in14[5]);
  xnor csa_tree_add_51_79_groupi_g43698(csa_tree_add_51_79_groupi_n_2669 ,in11[1] ,in12[5]);
  xnor csa_tree_add_51_79_groupi_g43699(csa_tree_add_51_79_groupi_n_2668 ,in17[7] ,in18[7]);
  xnor csa_tree_add_51_79_groupi_g43700(csa_tree_add_51_79_groupi_n_2667 ,in3[5] ,in4[1]);
  xnor csa_tree_add_51_79_groupi_g43701(csa_tree_add_51_79_groupi_n_2666 ,in17[9] ,in18[5]);
  xnor csa_tree_add_51_79_groupi_g43702(csa_tree_add_51_79_groupi_n_2665 ,in9[3] ,in10[3]);
  xnor csa_tree_add_51_79_groupi_g43703(csa_tree_add_51_79_groupi_n_2664 ,in9[3] ,in10[5]);
  xnor csa_tree_add_51_79_groupi_g43704(csa_tree_add_51_79_groupi_n_2663 ,in5[9] ,in6[5]);
  xnor csa_tree_add_51_79_groupi_g43705(csa_tree_add_51_79_groupi_n_2662 ,in15[7] ,in16[5]);
  xnor csa_tree_add_51_79_groupi_g43706(csa_tree_add_51_79_groupi_n_2661 ,in13[8] ,in14[3]);
  xnor csa_tree_add_51_79_groupi_g43707(csa_tree_add_51_79_groupi_n_2660 ,in17[1] ,in18[7]);
  xnor csa_tree_add_51_79_groupi_g43708(csa_tree_add_51_79_groupi_n_2659 ,in21[6] ,in22[5]);
  xnor csa_tree_add_51_79_groupi_g43709(csa_tree_add_51_79_groupi_n_2658 ,in7[6] ,in8[5]);
  xnor csa_tree_add_51_79_groupi_g43710(csa_tree_add_51_79_groupi_n_2657 ,in23[5] ,in24[1]);
  xnor csa_tree_add_51_79_groupi_g43711(csa_tree_add_51_79_groupi_n_2656 ,in3[2] ,in4[1]);
  xnor csa_tree_add_51_79_groupi_g43712(csa_tree_add_51_79_groupi_n_2654 ,csa_tree_add_51_79_groupi_n_1128 ,in7[10]);
  xnor csa_tree_add_51_79_groupi_g43713(csa_tree_add_51_79_groupi_n_2653 ,in11[10] ,in12[1]);
  xnor csa_tree_add_51_79_groupi_g43714(csa_tree_add_51_79_groupi_n_2652 ,in1[9] ,in2[7]);
  xnor csa_tree_add_51_79_groupi_g43715(csa_tree_add_51_79_groupi_n_2651 ,in7[7] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g43716(csa_tree_add_51_79_groupi_n_2650 ,in7[2] ,in8[5]);
  xnor csa_tree_add_51_79_groupi_g43717(csa_tree_add_51_79_groupi_n_2649 ,in15[10] ,in16[7]);
  xnor csa_tree_add_51_79_groupi_g43718(csa_tree_add_51_79_groupi_n_2648 ,in3[7] ,in4[7]);
  xnor csa_tree_add_51_79_groupi_g43719(csa_tree_add_51_79_groupi_n_2647 ,in13[9] ,in14[3]);
  xnor csa_tree_add_51_79_groupi_g43720(csa_tree_add_51_79_groupi_n_2646 ,in21[1] ,in22[5]);
  xnor csa_tree_add_51_79_groupi_g43721(csa_tree_add_51_79_groupi_n_2645 ,in17[3] ,in18[3]);
  xnor csa_tree_add_51_79_groupi_g43722(csa_tree_add_51_79_groupi_n_2644 ,in21[2] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g43723(csa_tree_add_51_79_groupi_n_2643 ,in23[9] ,in24[3]);
  xnor csa_tree_add_51_79_groupi_g43724(csa_tree_add_51_79_groupi_n_2642 ,in23[3] ,in24[3]);
  xnor csa_tree_add_51_79_groupi_g43725(csa_tree_add_51_79_groupi_n_2641 ,in1[1] ,in2[3]);
  xnor csa_tree_add_51_79_groupi_g43726(csa_tree_add_51_79_groupi_n_2640 ,in9[4] ,in10[5]);
  xnor csa_tree_add_51_79_groupi_g43727(csa_tree_add_51_79_groupi_n_2639 ,in7[4] ,in8[7]);
  xnor csa_tree_add_51_79_groupi_g43728(csa_tree_add_51_79_groupi_n_2638 ,in9[7] ,in10[5]);
  xnor csa_tree_add_51_79_groupi_g43729(csa_tree_add_51_79_groupi_n_2637 ,in15[2] ,in16[5]);
  xnor csa_tree_add_51_79_groupi_g43730(csa_tree_add_51_79_groupi_n_2636 ,in17[3] ,in18[1]);
  xnor csa_tree_add_51_79_groupi_g43731(csa_tree_add_51_79_groupi_n_2635 ,in23[10] ,in24[1]);
  xnor csa_tree_add_51_79_groupi_g43732(csa_tree_add_51_79_groupi_n_2634 ,in3[4] ,in4[7]);
  xnor csa_tree_add_51_79_groupi_g43733(csa_tree_add_51_79_groupi_n_2633 ,in1[3] ,in2[3]);
  xnor csa_tree_add_51_79_groupi_g43734(csa_tree_add_51_79_groupi_n_2632 ,in23[1] ,in24[1]);
  xnor csa_tree_add_51_79_groupi_g43735(csa_tree_add_51_79_groupi_n_2631 ,in1[1] ,in2[1]);
  xnor csa_tree_add_51_79_groupi_g43736(csa_tree_add_51_79_groupi_n_2630 ,in15[6] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g43737(csa_tree_add_51_79_groupi_n_2629 ,in11[4] ,in12[5]);
  xnor csa_tree_add_51_79_groupi_g43738(csa_tree_add_51_79_groupi_n_2628 ,in21[3] ,in22[3]);
  xnor csa_tree_add_51_79_groupi_g43739(csa_tree_add_51_79_groupi_n_2627 ,in17[9] ,in18[1]);
  xnor csa_tree_add_51_79_groupi_g43740(csa_tree_add_51_79_groupi_n_2626 ,in3[2] ,in4[5]);
  xnor csa_tree_add_51_79_groupi_g43741(csa_tree_add_51_79_groupi_n_2625 ,in11[3] ,in12[1]);
  xnor csa_tree_add_51_79_groupi_g43742(csa_tree_add_51_79_groupi_n_2624 ,in7[1] ,in8[5]);
  xnor csa_tree_add_51_79_groupi_g43743(csa_tree_add_51_79_groupi_n_2623 ,in23[6] ,in24[7]);
  xnor csa_tree_add_51_79_groupi_g43744(csa_tree_add_51_79_groupi_n_2622 ,in15[9] ,in16[3]);
  xnor csa_tree_add_51_79_groupi_g43745(csa_tree_add_51_79_groupi_n_2621 ,in7[3] ,in8[7]);
  xnor csa_tree_add_51_79_groupi_g43746(csa_tree_add_51_79_groupi_n_2620 ,in5[3] ,in6[3]);
  xnor csa_tree_add_51_79_groupi_g43747(csa_tree_add_51_79_groupi_n_2619 ,in9[4] ,in10[1]);
  xnor csa_tree_add_51_79_groupi_g43748(csa_tree_add_51_79_groupi_n_2618 ,in23[10] ,in24[7]);
  xnor csa_tree_add_51_79_groupi_g43749(csa_tree_add_51_79_groupi_n_2617 ,in13[10] ,in14[7]);
  xnor csa_tree_add_51_79_groupi_g43750(csa_tree_add_51_79_groupi_n_2616 ,in3[1] ,in4[5]);
  xnor csa_tree_add_51_79_groupi_g43751(csa_tree_add_51_79_groupi_n_2615 ,in15[2] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g43752(csa_tree_add_51_79_groupi_n_2614 ,in15[3] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g43753(csa_tree_add_51_79_groupi_n_2613 ,in7[9] ,in8[3]);
  xnor csa_tree_add_51_79_groupi_g43754(csa_tree_add_51_79_groupi_n_2612 ,in11[7] ,in12[3]);
  xnor csa_tree_add_51_79_groupi_g43755(csa_tree_add_51_79_groupi_n_2611 ,in7[10] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g43756(csa_tree_add_51_79_groupi_n_2610 ,in9[8] ,in10[1]);
  xnor csa_tree_add_51_79_groupi_g43757(csa_tree_add_51_79_groupi_n_2609 ,in5[3] ,in6[7]);
  xnor csa_tree_add_51_79_groupi_g43758(csa_tree_add_51_79_groupi_n_2608 ,in9[9] ,in10[5]);
  xnor csa_tree_add_51_79_groupi_g43759(csa_tree_add_51_79_groupi_n_2607 ,in11[10] ,in12[5]);
  xnor csa_tree_add_51_79_groupi_g43760(csa_tree_add_51_79_groupi_n_2606 ,in1[7] ,in2[7]);
  xnor csa_tree_add_51_79_groupi_g43761(csa_tree_add_51_79_groupi_n_2605 ,in13[6] ,in14[3]);
  xnor csa_tree_add_51_79_groupi_g43762(csa_tree_add_51_79_groupi_n_2604 ,in17[3] ,in18[7]);
  xnor csa_tree_add_51_79_groupi_g43763(csa_tree_add_51_79_groupi_n_2603 ,in3[10] ,in4[1]);
  xnor csa_tree_add_51_79_groupi_g43764(csa_tree_add_51_79_groupi_n_2602 ,in5[8] ,in6[5]);
  xnor csa_tree_add_51_79_groupi_g43765(csa_tree_add_51_79_groupi_n_2601 ,in13[10] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g43766(csa_tree_add_51_79_groupi_n_2600 ,in19[10] ,in20[7]);
  xnor csa_tree_add_51_79_groupi_g43767(csa_tree_add_51_79_groupi_n_2599 ,in9[5] ,in10[3]);
  xnor csa_tree_add_51_79_groupi_g43768(csa_tree_add_51_79_groupi_n_2598 ,in15[8] ,in16[3]);
  xnor csa_tree_add_51_79_groupi_g43769(csa_tree_add_51_79_groupi_n_2597 ,in11[2] ,in12[5]);
  xnor csa_tree_add_51_79_groupi_g43770(csa_tree_add_51_79_groupi_n_2596 ,in13[9] ,in14[5]);
  xnor csa_tree_add_51_79_groupi_g43771(csa_tree_add_51_79_groupi_n_2595 ,in17[9] ,in18[3]);
  xnor csa_tree_add_51_79_groupi_g43772(csa_tree_add_51_79_groupi_n_2594 ,in7[2] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g43773(csa_tree_add_51_79_groupi_n_2593 ,in15[5] ,in16[3]);
  xnor csa_tree_add_51_79_groupi_g43774(csa_tree_add_51_79_groupi_n_2592 ,in11[4] ,in12[7]);
  xnor csa_tree_add_51_79_groupi_g43775(csa_tree_add_51_79_groupi_n_2591 ,in7[8] ,in8[3]);
  xnor csa_tree_add_51_79_groupi_g43776(csa_tree_add_51_79_groupi_n_2589 ,csa_tree_add_51_79_groupi_n_1144 ,in3[10]);
  xnor csa_tree_add_51_79_groupi_g43777(csa_tree_add_51_79_groupi_n_2588 ,in15[4] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g43778(csa_tree_add_51_79_groupi_n_2587 ,in23[5] ,in24[5]);
  xnor csa_tree_add_51_79_groupi_g43779(csa_tree_add_51_79_groupi_n_2586 ,in7[1] ,in8[7]);
  xnor csa_tree_add_51_79_groupi_g43780(csa_tree_add_51_79_groupi_n_2585 ,in13[2] ,in14[3]);
  xnor csa_tree_add_51_79_groupi_g43781(csa_tree_add_51_79_groupi_n_2584 ,in1[4] ,in2[1]);
  xnor csa_tree_add_51_79_groupi_g43782(csa_tree_add_51_79_groupi_n_2583 ,in19[7] ,in20[7]);
  xnor csa_tree_add_51_79_groupi_g43783(csa_tree_add_51_79_groupi_n_2582 ,in15[2] ,in16[3]);
  xnor csa_tree_add_51_79_groupi_g43784(csa_tree_add_51_79_groupi_n_2581 ,in17[8] ,in18[3]);
  xnor csa_tree_add_51_79_groupi_g43785(csa_tree_add_51_79_groupi_n_2580 ,in17[1] ,in18[1]);
  xnor csa_tree_add_51_79_groupi_g43786(csa_tree_add_51_79_groupi_n_2579 ,in13[8] ,in14[7]);
  xnor csa_tree_add_51_79_groupi_g43787(csa_tree_add_51_79_groupi_n_2578 ,in19[1] ,in20[1]);
  xnor csa_tree_add_51_79_groupi_g43788(csa_tree_add_51_79_groupi_n_2577 ,in9[10] ,in10[3]);
  xnor csa_tree_add_51_79_groupi_g43789(csa_tree_add_51_79_groupi_n_2576 ,in13[3] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g43790(csa_tree_add_51_79_groupi_n_2575 ,in5[10] ,in6[5]);
  xnor csa_tree_add_51_79_groupi_g43791(csa_tree_add_51_79_groupi_n_2574 ,in11[4] ,in12[1]);
  xnor csa_tree_add_51_79_groupi_g43792(csa_tree_add_51_79_groupi_n_2573 ,in23[2] ,in24[3]);
  xnor csa_tree_add_51_79_groupi_g43793(csa_tree_add_51_79_groupi_n_2572 ,in21[8] ,in22[3]);
  or csa_tree_add_51_79_groupi_g43794(csa_tree_add_51_79_groupi_n_2571 ,csa_tree_add_51_79_groupi_n_1617 ,csa_tree_add_51_79_groupi_n_1720);
  or csa_tree_add_51_79_groupi_g43795(csa_tree_add_51_79_groupi_n_2570 ,csa_tree_add_51_79_groupi_n_1550 ,csa_tree_add_51_79_groupi_n_1775);
  or csa_tree_add_51_79_groupi_g43796(csa_tree_add_51_79_groupi_n_2568 ,csa_tree_add_51_79_groupi_n_1542 ,csa_tree_add_51_79_groupi_n_1784);
  and csa_tree_add_51_79_groupi_g43797(csa_tree_add_51_79_groupi_n_2567 ,csa_tree_add_51_79_groupi_n_838 ,csa_tree_add_51_79_groupi_n_1664);
  or csa_tree_add_51_79_groupi_g43798(csa_tree_add_51_79_groupi_n_2566 ,in3[0] ,csa_tree_add_51_79_groupi_n_1671);
  or csa_tree_add_51_79_groupi_g43799(csa_tree_add_51_79_groupi_n_2565 ,in19[0] ,csa_tree_add_51_79_groupi_n_1672);
  or csa_tree_add_51_79_groupi_g43800(csa_tree_add_51_79_groupi_n_2563 ,csa_tree_add_51_79_groupi_n_1539 ,csa_tree_add_51_79_groupi_n_1721);
  or csa_tree_add_51_79_groupi_g43801(csa_tree_add_51_79_groupi_n_2562 ,csa_tree_add_51_79_groupi_n_1601 ,csa_tree_add_51_79_groupi_n_1722);
  or csa_tree_add_51_79_groupi_g43802(csa_tree_add_51_79_groupi_n_2561 ,csa_tree_add_51_79_groupi_n_1540 ,csa_tree_add_51_79_groupi_n_1786);
  and csa_tree_add_51_79_groupi_g43803(csa_tree_add_51_79_groupi_n_2559 ,csa_tree_add_51_79_groupi_n_840 ,csa_tree_add_51_79_groupi_n_1663);
  or csa_tree_add_51_79_groupi_g43804(csa_tree_add_51_79_groupi_n_2558 ,csa_tree_add_51_79_groupi_n_1537 ,csa_tree_add_51_79_groupi_n_1777);
  or csa_tree_add_51_79_groupi_g43805(csa_tree_add_51_79_groupi_n_2557 ,csa_tree_add_51_79_groupi_n_1610 ,csa_tree_add_51_79_groupi_n_1782);
  or csa_tree_add_51_79_groupi_g43806(csa_tree_add_51_79_groupi_n_2556 ,csa_tree_add_51_79_groupi_n_1606 ,csa_tree_add_51_79_groupi_n_1778);
  or csa_tree_add_51_79_groupi_g43807(csa_tree_add_51_79_groupi_n_2555 ,csa_tree_add_51_79_groupi_n_1785 ,csa_tree_add_51_79_groupi_n_1779);
  or csa_tree_add_51_79_groupi_g43808(csa_tree_add_51_79_groupi_n_2554 ,csa_tree_add_51_79_groupi_n_1612 ,csa_tree_add_51_79_groupi_n_1774);
  or csa_tree_add_51_79_groupi_g43809(csa_tree_add_51_79_groupi_n_2553 ,csa_tree_add_51_79_groupi_n_1599 ,csa_tree_add_51_79_groupi_n_1776);
  or csa_tree_add_51_79_groupi_g43810(csa_tree_add_51_79_groupi_n_2552 ,csa_tree_add_51_79_groupi_n_1607 ,csa_tree_add_51_79_groupi_n_1780);
  or csa_tree_add_51_79_groupi_g43811(csa_tree_add_51_79_groupi_n_2551 ,in23[0] ,csa_tree_add_51_79_groupi_n_1667);
  and csa_tree_add_51_79_groupi_g43812(csa_tree_add_51_79_groupi_n_2550 ,csa_tree_add_51_79_groupi_n_836 ,csa_tree_add_51_79_groupi_n_1674);
  and csa_tree_add_51_79_groupi_g43813(csa_tree_add_51_79_groupi_n_2548 ,csa_tree_add_51_79_groupi_n_850 ,csa_tree_add_51_79_groupi_n_1665);
  and csa_tree_add_51_79_groupi_g43814(csa_tree_add_51_79_groupi_n_2547 ,csa_tree_add_51_79_groupi_n_846 ,csa_tree_add_51_79_groupi_n_1666);
  and csa_tree_add_51_79_groupi_g43815(csa_tree_add_51_79_groupi_n_2545 ,csa_tree_add_51_79_groupi_n_848 ,csa_tree_add_51_79_groupi_n_1670);
  and csa_tree_add_51_79_groupi_g43816(csa_tree_add_51_79_groupi_n_2544 ,csa_tree_add_51_79_groupi_n_852 ,csa_tree_add_51_79_groupi_n_1669);
  and csa_tree_add_51_79_groupi_g43817(csa_tree_add_51_79_groupi_n_2543 ,csa_tree_add_51_79_groupi_n_842 ,csa_tree_add_51_79_groupi_n_1673);
  and csa_tree_add_51_79_groupi_g43818(csa_tree_add_51_79_groupi_n_2541 ,csa_tree_add_51_79_groupi_n_844 ,csa_tree_add_51_79_groupi_n_1668);
  xnor csa_tree_add_51_79_groupi_g43819(csa_tree_add_51_79_groupi_n_2539 ,in10[10] ,in10[9]);
  xnor csa_tree_add_51_79_groupi_g43820(csa_tree_add_51_79_groupi_n_2535 ,csa_tree_add_51_79_groupi_n_1624 ,in2[10]);
  xnor csa_tree_add_51_79_groupi_g43821(csa_tree_add_51_79_groupi_n_2532 ,in12[10] ,in12[9]);
  xnor csa_tree_add_51_79_groupi_g43822(csa_tree_add_51_79_groupi_n_2531 ,in6[10] ,in6[9]);
  xnor csa_tree_add_51_79_groupi_g43823(csa_tree_add_51_79_groupi_n_2528 ,csa_tree_add_51_79_groupi_n_1555 ,in8[10]);
  xnor csa_tree_add_51_79_groupi_g43824(csa_tree_add_51_79_groupi_n_2527 ,in4[10] ,in4[9]);
  xnor csa_tree_add_51_79_groupi_g43825(csa_tree_add_51_79_groupi_n_2525 ,in22[10] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g43826(csa_tree_add_51_79_groupi_n_2523 ,in16[10] ,in16[9]);
  xnor csa_tree_add_51_79_groupi_g43827(csa_tree_add_51_79_groupi_n_2521 ,in24[10] ,in24[9]);
  xnor csa_tree_add_51_79_groupi_g43828(csa_tree_add_51_79_groupi_n_2519 ,in20[10] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g43829(csa_tree_add_51_79_groupi_n_2516 ,in14[10] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g43830(csa_tree_add_51_79_groupi_n_2514 ,in18[10] ,in18[9]);
  xor csa_tree_add_51_79_groupi_g43831(csa_tree_add_51_79_groupi_n_2511 ,in12[2] ,in12[1]);
  xnor csa_tree_add_51_79_groupi_g43832(csa_tree_add_51_79_groupi_n_2508 ,csa_tree_add_51_79_groupi_n_1620 ,in4[6]);
  xnor csa_tree_add_51_79_groupi_g43833(csa_tree_add_51_79_groupi_n_2506 ,csa_tree_add_51_79_groupi_n_1544 ,in6[8]);
  xnor csa_tree_add_51_79_groupi_g43834(csa_tree_add_51_79_groupi_n_2503 ,csa_tree_add_51_79_groupi_n_1552 ,in12[4]);
  xnor csa_tree_add_51_79_groupi_g43835(csa_tree_add_51_79_groupi_n_2501 ,csa_tree_add_51_79_groupi_n_1146 ,in10[8]);
  xnor csa_tree_add_51_79_groupi_g43836(csa_tree_add_51_79_groupi_n_2498 ,csa_tree_add_51_79_groupi_n_1140 ,in20[4]);
  xnor csa_tree_add_51_79_groupi_g43837(csa_tree_add_51_79_groupi_n_2495 ,csa_tree_add_51_79_groupi_n_1604 ,in20[8]);
  xor csa_tree_add_51_79_groupi_g43838(csa_tree_add_51_79_groupi_n_2492 ,in14[2] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g43839(csa_tree_add_51_79_groupi_n_2489 ,csa_tree_add_51_79_groupi_n_1130 ,in6[4]);
  xnor csa_tree_add_51_79_groupi_g43840(csa_tree_add_51_79_groupi_n_2487 ,csa_tree_add_51_79_groupi_n_1596 ,in12[8]);
  xor csa_tree_add_51_79_groupi_g43841(csa_tree_add_51_79_groupi_n_2484 ,in22[2] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g43842(csa_tree_add_51_79_groupi_n_2481 ,csa_tree_add_51_79_groupi_n_1132 ,in2[6]);
  xor csa_tree_add_51_79_groupi_g43843(csa_tree_add_51_79_groupi_n_2479 ,in8[2] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g43844(csa_tree_add_51_79_groupi_n_2476 ,csa_tree_add_51_79_groupi_n_1615 ,in10[4]);
  xor csa_tree_add_51_79_groupi_g43845(csa_tree_add_51_79_groupi_n_2473 ,in16[2] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g43846(csa_tree_add_51_79_groupi_n_2470 ,csa_tree_add_51_79_groupi_n_1548 ,in14[8]);
  xnor csa_tree_add_51_79_groupi_g43847(csa_tree_add_51_79_groupi_n_2467 ,csa_tree_add_51_79_groupi_n_1608 ,in18[6]);
  xnor csa_tree_add_51_79_groupi_g43848(csa_tree_add_51_79_groupi_n_2464 ,csa_tree_add_51_79_groupi_n_1611 ,in6[6]);
  xor csa_tree_add_51_79_groupi_g43849(csa_tree_add_51_79_groupi_n_2461 ,in2[2] ,in2[1]);
  xnor csa_tree_add_51_79_groupi_g43850(csa_tree_add_51_79_groupi_n_2458 ,csa_tree_add_51_79_groupi_n_1549 ,in14[6]);
  xnor csa_tree_add_51_79_groupi_g43851(csa_tree_add_51_79_groupi_n_2455 ,csa_tree_add_51_79_groupi_n_1531 ,in22[6]);
  xor csa_tree_add_51_79_groupi_g43852(csa_tree_add_51_79_groupi_n_2453 ,in6[2] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g43853(csa_tree_add_51_79_groupi_n_2450 ,csa_tree_add_51_79_groupi_n_1597 ,in16[4]);
  xnor csa_tree_add_51_79_groupi_g43854(csa_tree_add_51_79_groupi_n_2447 ,csa_tree_add_51_79_groupi_n_1541 ,in22[4]);
  xnor csa_tree_add_51_79_groupi_g43855(csa_tree_add_51_79_groupi_n_2445 ,csa_tree_add_51_79_groupi_n_1616 ,in10[6]);
  xnor csa_tree_add_51_79_groupi_g43856(csa_tree_add_51_79_groupi_n_2442 ,csa_tree_add_51_79_groupi_n_1551 ,in18[8]);
  xnor csa_tree_add_51_79_groupi_g43857(csa_tree_add_51_79_groupi_n_2439 ,csa_tree_add_51_79_groupi_n_1534 ,in20[6]);
  xnor csa_tree_add_51_79_groupi_g43858(csa_tree_add_51_79_groupi_n_2436 ,csa_tree_add_51_79_groupi_n_1614 ,in4[4]);
  xnor csa_tree_add_51_79_groupi_g43859(csa_tree_add_51_79_groupi_n_2434 ,csa_tree_add_51_79_groupi_n_1613 ,in2[8]);
  not csa_tree_add_51_79_groupi_g43860(csa_tree_add_51_79_groupi_n_2282 ,csa_tree_add_51_79_groupi_n_2281);
  not csa_tree_add_51_79_groupi_g43861(csa_tree_add_51_79_groupi_n_2264 ,csa_tree_add_51_79_groupi_n_2263);
  not csa_tree_add_51_79_groupi_g43862(csa_tree_add_51_79_groupi_n_2257 ,csa_tree_add_51_79_groupi_n_2256);
  not csa_tree_add_51_79_groupi_g43863(csa_tree_add_51_79_groupi_n_2255 ,csa_tree_add_51_79_groupi_n_2254);
  not csa_tree_add_51_79_groupi_g43864(csa_tree_add_51_79_groupi_n_2229 ,csa_tree_add_51_79_groupi_n_2228);
  not csa_tree_add_51_79_groupi_g43865(csa_tree_add_51_79_groupi_n_2202 ,csa_tree_add_51_79_groupi_n_2201);
  not csa_tree_add_51_79_groupi_g43866(csa_tree_add_51_79_groupi_n_2175 ,csa_tree_add_51_79_groupi_n_2174);
  not csa_tree_add_51_79_groupi_g43867(csa_tree_add_51_79_groupi_n_2167 ,csa_tree_add_51_79_groupi_n_2166);
  not csa_tree_add_51_79_groupi_g43868(csa_tree_add_51_79_groupi_n_2147 ,csa_tree_add_51_79_groupi_n_2146);
  not csa_tree_add_51_79_groupi_g43869(csa_tree_add_51_79_groupi_n_2121 ,csa_tree_add_51_79_groupi_n_2120);
  not csa_tree_add_51_79_groupi_g43870(csa_tree_add_51_79_groupi_n_2118 ,csa_tree_add_51_79_groupi_n_2117);
  not csa_tree_add_51_79_groupi_g43871(csa_tree_add_51_79_groupi_n_2107 ,csa_tree_add_51_79_groupi_n_2106);
  not csa_tree_add_51_79_groupi_g43872(csa_tree_add_51_79_groupi_n_2101 ,csa_tree_add_51_79_groupi_n_2100);
  not csa_tree_add_51_79_groupi_g43873(csa_tree_add_51_79_groupi_n_2024 ,csa_tree_add_51_79_groupi_n_2023);
  not csa_tree_add_51_79_groupi_g43874(csa_tree_add_51_79_groupi_n_2014 ,csa_tree_add_51_79_groupi_n_2012);
  not csa_tree_add_51_79_groupi_g43877(csa_tree_add_51_79_groupi_n_2011 ,csa_tree_add_51_79_groupi_n_2009);
  not csa_tree_add_51_79_groupi_g43880(csa_tree_add_51_79_groupi_n_2008 ,csa_tree_add_51_79_groupi_n_2006);
  not csa_tree_add_51_79_groupi_g43883(csa_tree_add_51_79_groupi_n_2005 ,csa_tree_add_51_79_groupi_n_2003);
  not csa_tree_add_51_79_groupi_g43886(csa_tree_add_51_79_groupi_n_2002 ,csa_tree_add_51_79_groupi_n_2000);
  not csa_tree_add_51_79_groupi_g43893(csa_tree_add_51_79_groupi_n_1995 ,csa_tree_add_51_79_groupi_n_1993);
  not csa_tree_add_51_79_groupi_g43912(csa_tree_add_51_79_groupi_n_1976 ,csa_tree_add_51_79_groupi_n_1974);
  not csa_tree_add_51_79_groupi_g43915(csa_tree_add_51_79_groupi_n_1973 ,csa_tree_add_51_79_groupi_n_1971);
  not csa_tree_add_51_79_groupi_g43918(csa_tree_add_51_79_groupi_n_1970 ,csa_tree_add_51_79_groupi_n_1968);
  xor csa_tree_add_51_79_groupi_g43921(csa_tree_add_51_79_groupi_n_1967 ,in1[10] ,in2[10]);
  xnor csa_tree_add_51_79_groupi_g43922(csa_tree_add_51_79_groupi_n_1966 ,in16[7] ,in16[6]);
  xnor csa_tree_add_51_79_groupi_g43923(csa_tree_add_51_79_groupi_n_1965 ,in19[0] ,in20[5]);
  xor csa_tree_add_51_79_groupi_g43924(csa_tree_add_51_79_groupi_n_1964 ,in17[3] ,in18[10]);
  xor csa_tree_add_51_79_groupi_g43925(csa_tree_add_51_79_groupi_n_1963 ,in23[1] ,in24[10]);
  xor csa_tree_add_51_79_groupi_g43926(csa_tree_add_51_79_groupi_n_1962 ,in21[2] ,in22[10]);
  xor csa_tree_add_51_79_groupi_g43927(csa_tree_add_51_79_groupi_n_1961 ,in17[10] ,in18[10]);
  xor csa_tree_add_51_79_groupi_g43928(csa_tree_add_51_79_groupi_n_1960 ,in19[2] ,in20[10]);
  xnor csa_tree_add_51_79_groupi_g43929(csa_tree_add_51_79_groupi_n_1959 ,in1[3] ,in2[10]);
  xnor csa_tree_add_51_79_groupi_g43930(csa_tree_add_51_79_groupi_n_1958 ,in1[0] ,in2[3]);
  xor csa_tree_add_51_79_groupi_g43931(csa_tree_add_51_79_groupi_n_1957 ,in21[3] ,in22[10]);
  xnor csa_tree_add_51_79_groupi_g43932(csa_tree_add_51_79_groupi_n_1956 ,in15[0] ,in16[3]);
  xor csa_tree_add_51_79_groupi_g43933(csa_tree_add_51_79_groupi_n_1955 ,in13[9] ,in14[10]);
  xor csa_tree_add_51_79_groupi_g43934(csa_tree_add_51_79_groupi_n_1954 ,in15[9] ,in16[10]);
  xnor csa_tree_add_51_79_groupi_g43935(csa_tree_add_51_79_groupi_n_1953 ,in21[0] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g43936(csa_tree_add_51_79_groupi_n_1952 ,in15[7] ,in16[10]);
  xor csa_tree_add_51_79_groupi_g43937(csa_tree_add_51_79_groupi_n_1951 ,in13[3] ,in14[10]);
  xnor csa_tree_add_51_79_groupi_g43938(csa_tree_add_51_79_groupi_n_1950 ,in21[7] ,in22[10]);
  xnor csa_tree_add_51_79_groupi_g43939(csa_tree_add_51_79_groupi_n_1949 ,in23[7] ,in24[10]);
  xor csa_tree_add_51_79_groupi_g43940(csa_tree_add_51_79_groupi_n_1948 ,in19[9] ,in20[10]);
  xor csa_tree_add_51_79_groupi_g43941(csa_tree_add_51_79_groupi_n_1947 ,in21[5] ,in22[10]);
  xor csa_tree_add_51_79_groupi_g43942(csa_tree_add_51_79_groupi_n_1946 ,in13[10] ,in14[10]);
  xor csa_tree_add_51_79_groupi_g43943(csa_tree_add_51_79_groupi_n_1945 ,in13[6] ,in14[10]);
  xor csa_tree_add_51_79_groupi_g43944(csa_tree_add_51_79_groupi_n_1944 ,in7[7] ,in8[10]);
  xor csa_tree_add_51_79_groupi_g43945(csa_tree_add_51_79_groupi_n_1943 ,in5[1] ,in6[10]);
  xor csa_tree_add_51_79_groupi_g43946(csa_tree_add_51_79_groupi_n_1942 ,in17[7] ,in18[10]);
  xor csa_tree_add_51_79_groupi_g43947(csa_tree_add_51_79_groupi_n_1941 ,in11[2] ,in12[10]);
  xnor csa_tree_add_51_79_groupi_g43948(csa_tree_add_51_79_groupi_n_1940 ,in7[0] ,in8[5]);
  xor csa_tree_add_51_79_groupi_g43949(csa_tree_add_51_79_groupi_n_1939 ,in1[1] ,in2[10]);
  xnor csa_tree_add_51_79_groupi_g43950(csa_tree_add_51_79_groupi_n_1938 ,in17[6] ,in18[10]);
  xor csa_tree_add_51_79_groupi_g43951(csa_tree_add_51_79_groupi_n_1937 ,in13[5] ,in14[10]);
  xor csa_tree_add_51_79_groupi_g43952(csa_tree_add_51_79_groupi_n_1936 ,in19[8] ,in20[10]);
  xor csa_tree_add_51_79_groupi_g43953(csa_tree_add_51_79_groupi_n_1935 ,in23[2] ,in24[10]);
  xor csa_tree_add_51_79_groupi_g43954(csa_tree_add_51_79_groupi_n_1934 ,in21[1] ,in22[10]);
  xnor csa_tree_add_51_79_groupi_g43955(csa_tree_add_51_79_groupi_n_1933 ,in9[0] ,in10[7]);
  xnor csa_tree_add_51_79_groupi_g43956(csa_tree_add_51_79_groupi_n_1932 ,in23[9] ,in24[10]);
  xnor csa_tree_add_51_79_groupi_g43957(csa_tree_add_51_79_groupi_n_1931 ,in19[6] ,in20[10]);
  xor csa_tree_add_51_79_groupi_g43958(csa_tree_add_51_79_groupi_n_1930 ,in19[4] ,in20[10]);
  xor csa_tree_add_51_79_groupi_g43959(csa_tree_add_51_79_groupi_n_1929 ,in11[4] ,in12[10]);
  xnor csa_tree_add_51_79_groupi_g43960(csa_tree_add_51_79_groupi_n_1928 ,in11[8] ,in12[10]);
  xor csa_tree_add_51_79_groupi_g43961(csa_tree_add_51_79_groupi_n_1927 ,in3[9] ,in4[10]);
  xor csa_tree_add_51_79_groupi_g43962(csa_tree_add_51_79_groupi_n_1926 ,in1[9] ,in2[10]);
  xnor csa_tree_add_51_79_groupi_g43963(csa_tree_add_51_79_groupi_n_1925 ,in13[0] ,in14[3]);
  xnor csa_tree_add_51_79_groupi_g43964(csa_tree_add_51_79_groupi_n_1924 ,in11[7] ,in12[10]);
  xor csa_tree_add_51_79_groupi_g43965(csa_tree_add_51_79_groupi_n_1923 ,in5[5] ,in6[10]);
  xor csa_tree_add_51_79_groupi_g43966(csa_tree_add_51_79_groupi_n_1922 ,in1[4] ,in2[10]);
  xnor csa_tree_add_51_79_groupi_g43967(csa_tree_add_51_79_groupi_n_1921 ,in10[5] ,in10[4]);
  xor csa_tree_add_51_79_groupi_g43968(csa_tree_add_51_79_groupi_n_1920 ,in3[8] ,in4[10]);
  xor csa_tree_add_51_79_groupi_g43969(csa_tree_add_51_79_groupi_n_1919 ,in5[3] ,in6[10]);
  xor csa_tree_add_51_79_groupi_g43970(csa_tree_add_51_79_groupi_n_1918 ,in3[4] ,in4[10]);
  xor csa_tree_add_51_79_groupi_g43972(csa_tree_add_51_79_groupi_n_1916 ,in17[9] ,in18[10]);
  xor csa_tree_add_51_79_groupi_g43973(csa_tree_add_51_79_groupi_n_1915 ,in13[7] ,in14[10]);
  xor csa_tree_add_51_79_groupi_g43974(csa_tree_add_51_79_groupi_n_1914 ,in9[4] ,in10[10]);
  xor csa_tree_add_51_79_groupi_g43975(csa_tree_add_51_79_groupi_n_1913 ,in19[1] ,in20[10]);
  xnor csa_tree_add_51_79_groupi_g43976(csa_tree_add_51_79_groupi_n_1912 ,in17[1] ,in18[10]);
  xnor csa_tree_add_51_79_groupi_g43977(csa_tree_add_51_79_groupi_n_1911 ,in5[2] ,in6[10]);
  xnor csa_tree_add_51_79_groupi_g43978(csa_tree_add_51_79_groupi_n_1910 ,in7[2] ,in8[10]);
  xor csa_tree_add_51_79_groupi_g43979(csa_tree_add_51_79_groupi_n_1909 ,in9[7] ,in10[10]);
  xnor csa_tree_add_51_79_groupi_g43980(csa_tree_add_51_79_groupi_n_1908 ,in19[0] ,in20[7]);
  xnor csa_tree_add_51_79_groupi_g43981(csa_tree_add_51_79_groupi_n_1907 ,in5[8] ,in6[10]);
  xor csa_tree_add_51_79_groupi_g43982(csa_tree_add_51_79_groupi_n_1906 ,in5[10] ,in6[10]);
  xor csa_tree_add_51_79_groupi_g43984(csa_tree_add_51_79_groupi_n_1904 ,in13[8] ,in14[10]);
  xor csa_tree_add_51_79_groupi_g43985(csa_tree_add_51_79_groupi_n_1903 ,in11[3] ,in12[10]);
  xnor csa_tree_add_51_79_groupi_g43986(csa_tree_add_51_79_groupi_n_1902 ,in1[5] ,in2[10]);
  xnor csa_tree_add_51_79_groupi_g43987(csa_tree_add_51_79_groupi_n_1901 ,in9[6] ,in10[10]);
  xor csa_tree_add_51_79_groupi_g43988(csa_tree_add_51_79_groupi_n_1900 ,in3[7] ,in4[10]);
  xnor csa_tree_add_51_79_groupi_g43989(csa_tree_add_51_79_groupi_n_1899 ,in17[0] ,in18[7]);
  xnor csa_tree_add_51_79_groupi_g43990(csa_tree_add_51_79_groupi_n_1898 ,in3[6] ,in4[10]);
  xor csa_tree_add_51_79_groupi_g43991(csa_tree_add_51_79_groupi_n_1897 ,in7[3] ,in8[10]);
  xnor csa_tree_add_51_79_groupi_g43992(csa_tree_add_51_79_groupi_n_1896 ,in21[0] ,in22[3]);
  xnor csa_tree_add_51_79_groupi_g43993(csa_tree_add_51_79_groupi_n_1895 ,in3[3] ,in4[10]);
  xor csa_tree_add_51_79_groupi_g43994(csa_tree_add_51_79_groupi_n_1894 ,in23[8] ,in24[10]);
  xnor csa_tree_add_51_79_groupi_g43995(csa_tree_add_51_79_groupi_n_1893 ,in23[0] ,in24[3]);
  xor csa_tree_add_51_79_groupi_g43996(csa_tree_add_51_79_groupi_n_1892 ,in15[3] ,in16[10]);
  xnor csa_tree_add_51_79_groupi_g43997(csa_tree_add_51_79_groupi_n_1891 ,in20[3] ,in20[2]);
  xor csa_tree_add_51_79_groupi_g43998(csa_tree_add_51_79_groupi_n_1890 ,in17[8] ,in18[10]);
  xor csa_tree_add_51_79_groupi_g43999(csa_tree_add_51_79_groupi_n_1889 ,in17[2] ,in18[10]);
  xor csa_tree_add_51_79_groupi_g44000(csa_tree_add_51_79_groupi_n_1888 ,in21[4] ,in22[10]);
  xnor csa_tree_add_51_79_groupi_g44001(csa_tree_add_51_79_groupi_n_1887 ,in1[8] ,in2[10]);
  xor csa_tree_add_51_79_groupi_g44002(csa_tree_add_51_79_groupi_n_1886 ,in9[1] ,in10[10]);
  xor csa_tree_add_51_79_groupi_g44003(csa_tree_add_51_79_groupi_n_1885 ,in19[7] ,in20[10]);
  xnor csa_tree_add_51_79_groupi_g44004(csa_tree_add_51_79_groupi_n_1884 ,in3[1] ,in4[10]);
  xor csa_tree_add_51_79_groupi_g44005(csa_tree_add_51_79_groupi_n_1883 ,in19[5] ,in20[10]);
  xnor csa_tree_add_51_79_groupi_g44006(csa_tree_add_51_79_groupi_n_1882 ,in8[3] ,in8[2]);
  xnor csa_tree_add_51_79_groupi_g44007(csa_tree_add_51_79_groupi_n_1881 ,in7[0] ,in8[3]);
  xor csa_tree_add_51_79_groupi_g44008(csa_tree_add_51_79_groupi_n_1880 ,in21[10] ,in22[10]);
  xor csa_tree_add_51_79_groupi_g44009(csa_tree_add_51_79_groupi_n_1879 ,in21[6] ,in22[10]);
  xor csa_tree_add_51_79_groupi_g44010(csa_tree_add_51_79_groupi_n_1878 ,in9[10] ,in10[10]);
  xor csa_tree_add_51_79_groupi_g44011(csa_tree_add_51_79_groupi_n_1877 ,in23[5] ,in24[10]);
  xnor csa_tree_add_51_79_groupi_g44012(csa_tree_add_51_79_groupi_n_1876 ,in11[0] ,in12[7]);
  xor csa_tree_add_51_79_groupi_g44013(csa_tree_add_51_79_groupi_n_1875 ,in3[2] ,in4[10]);
  xnor csa_tree_add_51_79_groupi_g44014(csa_tree_add_51_79_groupi_n_1874 ,in7[4] ,in8[10]);
  xor csa_tree_add_51_79_groupi_g44015(csa_tree_add_51_79_groupi_n_1873 ,in5[6] ,in6[10]);
  xnor csa_tree_add_51_79_groupi_g44016(csa_tree_add_51_79_groupi_n_1872 ,in7[6] ,in8[10]);
  xnor csa_tree_add_51_79_groupi_g44017(csa_tree_add_51_79_groupi_n_1871 ,in13[4] ,in14[10]);
  xor csa_tree_add_51_79_groupi_g44018(csa_tree_add_51_79_groupi_n_1870 ,in9[3] ,in10[10]);
  xor csa_tree_add_51_79_groupi_g44019(csa_tree_add_51_79_groupi_n_1869 ,in13[1] ,in14[10]);
  xor csa_tree_add_51_79_groupi_g44020(csa_tree_add_51_79_groupi_n_1868 ,in11[1] ,in12[10]);
  xor csa_tree_add_51_79_groupi_g44021(csa_tree_add_51_79_groupi_n_1867 ,in9[8] ,in10[10]);
  xnor csa_tree_add_51_79_groupi_g44022(csa_tree_add_51_79_groupi_n_1866 ,in7[1] ,in8[10]);
  xor csa_tree_add_51_79_groupi_g44023(csa_tree_add_51_79_groupi_n_1865 ,in13[2] ,in14[10]);
  xor csa_tree_add_51_79_groupi_g44024(csa_tree_add_51_79_groupi_n_1864 ,in9[9] ,in10[10]);
  xnor csa_tree_add_51_79_groupi_g44025(csa_tree_add_51_79_groupi_n_1863 ,in15[0] ,in16[5]);
  xor csa_tree_add_51_79_groupi_g44026(csa_tree_add_51_79_groupi_n_1862 ,in7[5] ,in8[10]);
  xor csa_tree_add_51_79_groupi_g44027(csa_tree_add_51_79_groupi_n_1861 ,in15[8] ,in16[10]);
  xnor csa_tree_add_51_79_groupi_g44028(csa_tree_add_51_79_groupi_n_1860 ,in11[5] ,in12[10]);
  xor csa_tree_add_51_79_groupi_g44029(csa_tree_add_51_79_groupi_n_1859 ,in5[9] ,in6[10]);
  xor csa_tree_add_51_79_groupi_g44030(csa_tree_add_51_79_groupi_n_1858 ,in9[2] ,in10[10]);
  xor csa_tree_add_51_79_groupi_g44031(csa_tree_add_51_79_groupi_n_1857 ,in15[2] ,in16[10]);
  xor csa_tree_add_51_79_groupi_g44032(csa_tree_add_51_79_groupi_n_1856 ,in23[6] ,in24[10]);
  xor csa_tree_add_51_79_groupi_g44033(csa_tree_add_51_79_groupi_n_1855 ,in15[5] ,in16[10]);
  xor csa_tree_add_51_79_groupi_g44034(csa_tree_add_51_79_groupi_n_1854 ,in19[3] ,in20[10]);
  xnor csa_tree_add_51_79_groupi_g44035(csa_tree_add_51_79_groupi_n_1853 ,in10[3] ,in10[2]);
  xor csa_tree_add_51_79_groupi_g44037(csa_tree_add_51_79_groupi_n_1851 ,in21[9] ,in22[10]);
  xor csa_tree_add_51_79_groupi_g44038(csa_tree_add_51_79_groupi_n_1850 ,in7[9] ,in8[10]);
  xor csa_tree_add_51_79_groupi_g44039(csa_tree_add_51_79_groupi_n_1849 ,in15[1] ,in16[10]);
  xor csa_tree_add_51_79_groupi_g44040(csa_tree_add_51_79_groupi_n_1848 ,in9[5] ,in10[10]);
  xnor csa_tree_add_51_79_groupi_g44041(csa_tree_add_51_79_groupi_n_1847 ,in5[4] ,in6[10]);
  xor csa_tree_add_51_79_groupi_g44042(csa_tree_add_51_79_groupi_n_1846 ,in1[7] ,in2[10]);
  xor csa_tree_add_51_79_groupi_g44043(csa_tree_add_51_79_groupi_n_1845 ,in5[7] ,in6[10]);
  xor csa_tree_add_51_79_groupi_g44044(csa_tree_add_51_79_groupi_n_1844 ,in17[5] ,in18[10]);
  xor csa_tree_add_51_79_groupi_g44045(csa_tree_add_51_79_groupi_n_1843 ,in1[2] ,in2[10]);
  xor csa_tree_add_51_79_groupi_g44046(csa_tree_add_51_79_groupi_n_1842 ,in3[5] ,in4[10]);
  xor csa_tree_add_51_79_groupi_g44047(csa_tree_add_51_79_groupi_n_1841 ,in17[4] ,in18[10]);
  xor csa_tree_add_51_79_groupi_g44048(csa_tree_add_51_79_groupi_n_1840 ,in21[8] ,in22[10]);
  xor csa_tree_add_51_79_groupi_g44049(csa_tree_add_51_79_groupi_n_1839 ,in23[4] ,in24[10]);
  xor csa_tree_add_51_79_groupi_g44050(csa_tree_add_51_79_groupi_n_1838 ,in23[3] ,in24[10]);
  xnor csa_tree_add_51_79_groupi_g44051(csa_tree_add_51_79_groupi_n_1837 ,in8[7] ,in8[6]);
  xnor csa_tree_add_51_79_groupi_g44052(csa_tree_add_51_79_groupi_n_1836 ,in15[6] ,in16[10]);
  xor csa_tree_add_51_79_groupi_g44053(csa_tree_add_51_79_groupi_n_1835 ,in7[8] ,in8[10]);
  xor csa_tree_add_51_79_groupi_g44054(csa_tree_add_51_79_groupi_n_1834 ,in19[10] ,in20[10]);
  xnor csa_tree_add_51_79_groupi_g44055(csa_tree_add_51_79_groupi_n_1833 ,in1[6] ,in2[10]);
  xnor csa_tree_add_51_79_groupi_g44056(csa_tree_add_51_79_groupi_n_1832 ,in23[10] ,in24[10]);
  xor csa_tree_add_51_79_groupi_g44057(csa_tree_add_51_79_groupi_n_1831 ,in11[6] ,in12[10]);
  xnor csa_tree_add_51_79_groupi_g44058(csa_tree_add_51_79_groupi_n_1830 ,in11[9] ,in12[10]);
  xor csa_tree_add_51_79_groupi_g44059(csa_tree_add_51_79_groupi_n_1829 ,in3[10] ,in4[10]);
  xor csa_tree_add_51_79_groupi_g44060(csa_tree_add_51_79_groupi_n_1828 ,in15[4] ,in16[10]);
  xor csa_tree_add_51_79_groupi_g44061(csa_tree_add_51_79_groupi_n_1827 ,in7[10] ,in8[10]);
  xnor csa_tree_add_51_79_groupi_g44062(csa_tree_add_51_79_groupi_n_1826 ,in11[10] ,in12[10]);
  xor csa_tree_add_51_79_groupi_g44063(csa_tree_add_51_79_groupi_n_1825 ,in15[10] ,in16[10]);
  xnor csa_tree_add_51_79_groupi_g44064(csa_tree_add_51_79_groupi_n_1824 ,in16[9] ,in16[8]);
  xnor csa_tree_add_51_79_groupi_g44065(csa_tree_add_51_79_groupi_n_1823 ,in9[0] ,in10[9]);
  xnor csa_tree_add_51_79_groupi_g44066(csa_tree_add_51_79_groupi_n_1822 ,in19[0] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g44067(csa_tree_add_51_79_groupi_n_1821 ,in15[0] ,in16[9]);
  xnor csa_tree_add_51_79_groupi_g44068(csa_tree_add_51_79_groupi_n_1820 ,in18[3] ,in18[2]);
  xnor csa_tree_add_51_79_groupi_g44070(csa_tree_add_51_79_groupi_n_1818 ,in1[0] ,in2[9]);
  xnor csa_tree_add_51_79_groupi_g44071(csa_tree_add_51_79_groupi_n_1817 ,in21[0] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g44072(csa_tree_add_51_79_groupi_n_1816 ,in3[0] ,in4[9]);
  xnor csa_tree_add_51_79_groupi_g44073(csa_tree_add_51_79_groupi_n_1815 ,in11[0] ,in12[9]);
  xnor csa_tree_add_51_79_groupi_g44074(csa_tree_add_51_79_groupi_n_1814 ,in17[0] ,in18[9]);
  xnor csa_tree_add_51_79_groupi_g44075(csa_tree_add_51_79_groupi_n_1813 ,in3[0] ,in4[5]);
  xnor csa_tree_add_51_79_groupi_g44076(csa_tree_add_51_79_groupi_n_1812 ,in24[9] ,in24[8]);
  xnor csa_tree_add_51_79_groupi_g44077(csa_tree_add_51_79_groupi_n_1811 ,in4[9] ,in4[8]);
  xnor csa_tree_add_51_79_groupi_g44078(csa_tree_add_51_79_groupi_n_1810 ,in6[9] ,in6[8]);
  xnor csa_tree_add_51_79_groupi_g44079(csa_tree_add_51_79_groupi_n_1809 ,in10[9] ,in10[8]);
  xnor csa_tree_add_51_79_groupi_g44080(csa_tree_add_51_79_groupi_n_1808 ,in22[5] ,in22[4]);
  xnor csa_tree_add_51_79_groupi_g44081(csa_tree_add_51_79_groupi_n_1807 ,in8[5] ,in8[4]);
  xnor csa_tree_add_51_79_groupi_g44082(csa_tree_add_51_79_groupi_n_1806 ,in7[0] ,in8[9]);
  xnor csa_tree_add_51_79_groupi_g44083(csa_tree_add_51_79_groupi_n_1805 ,in22[9] ,in22[8]);
  xnor csa_tree_add_51_79_groupi_g44084(csa_tree_add_51_79_groupi_n_1804 ,in8[9] ,in8[8]);
  xnor csa_tree_add_51_79_groupi_g44085(csa_tree_add_51_79_groupi_n_1803 ,in5[0] ,in6[9]);
  xnor csa_tree_add_51_79_groupi_g44086(csa_tree_add_51_79_groupi_n_1802 ,in12[9] ,in12[8]);
  xnor csa_tree_add_51_79_groupi_g44087(csa_tree_add_51_79_groupi_n_1801 ,in20[9] ,in20[8]);
  xnor csa_tree_add_51_79_groupi_g44088(csa_tree_add_51_79_groupi_n_1800 ,in13[0] ,in14[5]);
  xnor csa_tree_add_51_79_groupi_g44089(csa_tree_add_51_79_groupi_n_1799 ,in23[0] ,in24[9]);
  xnor csa_tree_add_51_79_groupi_g44090(csa_tree_add_51_79_groupi_n_1798 ,in18[9] ,in18[8]);
  xnor csa_tree_add_51_79_groupi_g44091(csa_tree_add_51_79_groupi_n_1797 ,in13[0] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g44092(csa_tree_add_51_79_groupi_n_1796 ,in2[9] ,in2[8]);
  xnor csa_tree_add_51_79_groupi_g44093(csa_tree_add_51_79_groupi_n_1795 ,in14[9] ,in14[8]);
  xnor csa_tree_add_51_79_groupi_g44094(csa_tree_add_51_79_groupi_n_1794 ,in5[0] ,in6[3]);
  xnor csa_tree_add_51_79_groupi_g44095(csa_tree_add_51_79_groupi_n_1793 ,in7[0] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g44096(csa_tree_add_51_79_groupi_n_1792 ,in16[5] ,in16[4]);
  xnor csa_tree_add_51_79_groupi_g44097(csa_tree_add_51_79_groupi_n_1791 ,in4[5] ,in4[4]);
  xnor csa_tree_add_51_79_groupi_g44098(csa_tree_add_51_79_groupi_n_1790 ,in2[5] ,in2[4]);
  xnor csa_tree_add_51_79_groupi_g44099(csa_tree_add_51_79_groupi_n_1789 ,in14[5] ,in14[4]);
  xnor csa_tree_add_51_79_groupi_g44100(csa_tree_add_51_79_groupi_n_1788 ,in6[3] ,in6[2]);
  xnor csa_tree_add_51_79_groupi_g44101(csa_tree_add_51_79_groupi_n_2319 ,in9[8] ,in10[3]);
  xnor csa_tree_add_51_79_groupi_g44102(csa_tree_add_51_79_groupi_n_2318 ,in23[8] ,in24[3]);
  xnor csa_tree_add_51_79_groupi_g44103(csa_tree_add_51_79_groupi_n_2317 ,in13[4] ,in14[5]);
  xnor csa_tree_add_51_79_groupi_g44104(csa_tree_add_51_79_groupi_n_2316 ,in7[8] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g44105(csa_tree_add_51_79_groupi_n_2315 ,in23[8] ,in24[1]);
  xnor csa_tree_add_51_79_groupi_g44106(csa_tree_add_51_79_groupi_n_2314 ,in15[8] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g44107(csa_tree_add_51_79_groupi_n_2313 ,in7[6] ,in8[3]);
  xnor csa_tree_add_51_79_groupi_g44108(csa_tree_add_51_79_groupi_n_2312 ,in15[7] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g44109(csa_tree_add_51_79_groupi_n_2311 ,in1[1] ,in2[5]);
  xnor csa_tree_add_51_79_groupi_g44110(csa_tree_add_51_79_groupi_n_2310 ,in9[7] ,in10[3]);
  xnor csa_tree_add_51_79_groupi_g44111(csa_tree_add_51_79_groupi_n_2309 ,in19[5] ,in20[1]);
  xnor csa_tree_add_51_79_groupi_g44112(csa_tree_add_51_79_groupi_n_2308 ,in13[1] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g44113(csa_tree_add_51_79_groupi_n_2307 ,in1[5] ,in2[3]);
  xnor csa_tree_add_51_79_groupi_g44114(csa_tree_add_51_79_groupi_n_2306 ,in13[2] ,in14[7]);
  xnor csa_tree_add_51_79_groupi_g44115(csa_tree_add_51_79_groupi_n_2305 ,in11[3] ,in12[3]);
  xnor csa_tree_add_51_79_groupi_g44116(csa_tree_add_51_79_groupi_n_2304 ,in23[1] ,in24[5]);
  xnor csa_tree_add_51_79_groupi_g44117(csa_tree_add_51_79_groupi_n_2303 ,in15[6] ,in16[3]);
  xnor csa_tree_add_51_79_groupi_g44118(csa_tree_add_51_79_groupi_n_2302 ,in19[2] ,in20[7]);
  xnor csa_tree_add_51_79_groupi_g44119(csa_tree_add_51_79_groupi_n_2301 ,in3[6] ,in4[3]);
  xnor csa_tree_add_51_79_groupi_g44120(csa_tree_add_51_79_groupi_n_2300 ,in11[1] ,in12[1]);
  xnor csa_tree_add_51_79_groupi_g44121(csa_tree_add_51_79_groupi_n_2299 ,in1[9] ,in2[5]);
  xnor csa_tree_add_51_79_groupi_g44122(csa_tree_add_51_79_groupi_n_2298 ,in23[7] ,in24[1]);
  xnor csa_tree_add_51_79_groupi_g44123(csa_tree_add_51_79_groupi_n_2297 ,in9[3] ,in10[1]);
  xnor csa_tree_add_51_79_groupi_g44124(csa_tree_add_51_79_groupi_n_2296 ,in11[3] ,in12[7]);
  xnor csa_tree_add_51_79_groupi_g44125(csa_tree_add_51_79_groupi_n_2295 ,in15[2] ,in16[7]);
  xnor csa_tree_add_51_79_groupi_g44126(csa_tree_add_51_79_groupi_n_2294 ,in19[6] ,in20[7]);
  xnor csa_tree_add_51_79_groupi_g44127(csa_tree_add_51_79_groupi_n_2293 ,in5[8] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g44128(csa_tree_add_51_79_groupi_n_2292 ,in19[1] ,in20[5]);
  xnor csa_tree_add_51_79_groupi_g44129(csa_tree_add_51_79_groupi_n_2291 ,in17[9] ,in18[7]);
  xnor csa_tree_add_51_79_groupi_g44130(csa_tree_add_51_79_groupi_n_2290 ,in13[7] ,in14[5]);
  xnor csa_tree_add_51_79_groupi_g44131(csa_tree_add_51_79_groupi_n_2289 ,in15[4] ,in16[5]);
  xnor csa_tree_add_51_79_groupi_g44132(csa_tree_add_51_79_groupi_n_2288 ,in3[10] ,in4[5]);
  xnor csa_tree_add_51_79_groupi_g44133(csa_tree_add_51_79_groupi_n_2287 ,in19[5] ,in20[7]);
  xnor csa_tree_add_51_79_groupi_g44134(csa_tree_add_51_79_groupi_n_2286 ,in19[10] ,in20[5]);
  xnor csa_tree_add_51_79_groupi_g44135(csa_tree_add_51_79_groupi_n_2285 ,in17[5] ,in18[1]);
  xnor csa_tree_add_51_79_groupi_g44136(csa_tree_add_51_79_groupi_n_2284 ,in21[3] ,in22[5]);
  xnor csa_tree_add_51_79_groupi_g44137(csa_tree_add_51_79_groupi_n_2283 ,in11[6] ,in12[1]);
  xnor csa_tree_add_51_79_groupi_g44138(csa_tree_add_51_79_groupi_n_2281 ,csa_tree_add_51_79_groupi_n_1134 ,in23[10]);
  xnor csa_tree_add_51_79_groupi_g44139(csa_tree_add_51_79_groupi_n_2280 ,in3[5] ,in4[7]);
  xnor csa_tree_add_51_79_groupi_g44140(csa_tree_add_51_79_groupi_n_2279 ,in3[9] ,in4[5]);
  xnor csa_tree_add_51_79_groupi_g44141(csa_tree_add_51_79_groupi_n_2278 ,in9[1] ,in10[5]);
  xnor csa_tree_add_51_79_groupi_g44142(csa_tree_add_51_79_groupi_n_2277 ,in3[8] ,in4[7]);
  xnor csa_tree_add_51_79_groupi_g44143(csa_tree_add_51_79_groupi_n_2276 ,in15[5] ,in16[5]);
  xnor csa_tree_add_51_79_groupi_g44144(csa_tree_add_51_79_groupi_n_2275 ,in19[6] ,in20[3]);
  xnor csa_tree_add_51_79_groupi_g44145(csa_tree_add_51_79_groupi_n_2274 ,in23[2] ,in24[7]);
  xnor csa_tree_add_51_79_groupi_g44146(csa_tree_add_51_79_groupi_n_2273 ,in9[9] ,in10[9]);
  xnor csa_tree_add_51_79_groupi_g44147(csa_tree_add_51_79_groupi_n_2272 ,in17[1] ,in18[9]);
  xnor csa_tree_add_51_79_groupi_g44148(csa_tree_add_51_79_groupi_n_2271 ,in11[1] ,in12[9]);
  xnor csa_tree_add_51_79_groupi_g44149(csa_tree_add_51_79_groupi_n_2270 ,in15[1] ,in16[9]);
  xnor csa_tree_add_51_79_groupi_g44150(csa_tree_add_51_79_groupi_n_2269 ,in13[3] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g44151(csa_tree_add_51_79_groupi_n_2268 ,in15[8] ,in16[9]);
  xnor csa_tree_add_51_79_groupi_g44152(csa_tree_add_51_79_groupi_n_2267 ,in19[10] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g44153(csa_tree_add_51_79_groupi_n_2266 ,in1[3] ,in2[9]);
  xnor csa_tree_add_51_79_groupi_g44154(csa_tree_add_51_79_groupi_n_2265 ,in17[8] ,in18[9]);
  xnor csa_tree_add_51_79_groupi_g44155(csa_tree_add_51_79_groupi_n_2263 ,csa_tree_add_51_79_groupi_n_1126 ,in7[10]);
  xnor csa_tree_add_51_79_groupi_g44156(csa_tree_add_51_79_groupi_n_2262 ,in9[6] ,in10[9]);
  xnor csa_tree_add_51_79_groupi_g44157(csa_tree_add_51_79_groupi_n_2261 ,in21[4] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g44158(csa_tree_add_51_79_groupi_n_2260 ,in7[9] ,in8[9]);
  xnor csa_tree_add_51_79_groupi_g44159(csa_tree_add_51_79_groupi_n_2259 ,in15[5] ,in16[9]);
  xnor csa_tree_add_51_79_groupi_g44160(csa_tree_add_51_79_groupi_n_2258 ,in13[4] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g44161(csa_tree_add_51_79_groupi_n_2256 ,csa_tree_add_51_79_groupi_n_1627 ,in15[10]);
  xnor csa_tree_add_51_79_groupi_g44162(csa_tree_add_51_79_groupi_n_2254 ,csa_tree_add_51_79_groupi_n_1553 ,in23[10]);
  xnor csa_tree_add_51_79_groupi_g44163(csa_tree_add_51_79_groupi_n_2253 ,in3[6] ,in4[9]);
  xnor csa_tree_add_51_79_groupi_g44164(csa_tree_add_51_79_groupi_n_2252 ,in5[4] ,in6[5]);
  xnor csa_tree_add_51_79_groupi_g44165(csa_tree_add_51_79_groupi_n_2251 ,in17[9] ,in18[9]);
  xnor csa_tree_add_51_79_groupi_g44166(csa_tree_add_51_79_groupi_n_2250 ,in5[6] ,in6[3]);
  xnor csa_tree_add_51_79_groupi_g44167(csa_tree_add_51_79_groupi_n_2249 ,in7[2] ,in8[7]);
  xnor csa_tree_add_51_79_groupi_g44168(csa_tree_add_51_79_groupi_n_2248 ,in1[7] ,in2[9]);
  xnor csa_tree_add_51_79_groupi_g44169(csa_tree_add_51_79_groupi_n_2247 ,in7[4] ,in8[9]);
  xnor csa_tree_add_51_79_groupi_g44170(csa_tree_add_51_79_groupi_n_2246 ,in13[6] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g44171(csa_tree_add_51_79_groupi_n_2245 ,in21[6] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g44172(csa_tree_add_51_79_groupi_n_2244 ,in13[7] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g44173(csa_tree_add_51_79_groupi_n_2243 ,in19[4] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g44174(csa_tree_add_51_79_groupi_n_2242 ,in15[7] ,in16[9]);
  xnor csa_tree_add_51_79_groupi_g44175(csa_tree_add_51_79_groupi_n_2241 ,in13[5] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g44176(csa_tree_add_51_79_groupi_n_2240 ,in5[2] ,in6[7]);
  xnor csa_tree_add_51_79_groupi_g44177(csa_tree_add_51_79_groupi_n_2239 ,in15[6] ,in16[9]);
  xnor csa_tree_add_51_79_groupi_g44178(csa_tree_add_51_79_groupi_n_2238 ,in21[8] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g44179(csa_tree_add_51_79_groupi_n_2237 ,in9[7] ,in10[9]);
  xnor csa_tree_add_51_79_groupi_g44180(csa_tree_add_51_79_groupi_n_2236 ,in17[3] ,in18[9]);
  xnor csa_tree_add_51_79_groupi_g44181(csa_tree_add_51_79_groupi_n_2235 ,in23[9] ,in24[5]);
  xnor csa_tree_add_51_79_groupi_g44182(csa_tree_add_51_79_groupi_n_2234 ,in13[10] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g44183(csa_tree_add_51_79_groupi_n_2233 ,in1[8] ,in2[9]);
  xnor csa_tree_add_51_79_groupi_g44184(csa_tree_add_51_79_groupi_n_2232 ,in7[3] ,in8[9]);
  xnor csa_tree_add_51_79_groupi_g44185(csa_tree_add_51_79_groupi_n_2231 ,in5[7] ,in6[9]);
  xnor csa_tree_add_51_79_groupi_g44186(csa_tree_add_51_79_groupi_n_2230 ,in23[5] ,in24[9]);
  xnor csa_tree_add_51_79_groupi_g44187(csa_tree_add_51_79_groupi_n_2228 ,csa_tree_add_51_79_groupi_n_1625 ,in11[10]);
  xnor csa_tree_add_51_79_groupi_g44188(csa_tree_add_51_79_groupi_n_2227 ,in3[4] ,in4[9]);
  xnor csa_tree_add_51_79_groupi_g44189(csa_tree_add_51_79_groupi_n_2226 ,in3[2] ,in4[3]);
  xnor csa_tree_add_51_79_groupi_g44190(csa_tree_add_51_79_groupi_n_2225 ,in11[9] ,in12[9]);
  xnor csa_tree_add_51_79_groupi_g44191(csa_tree_add_51_79_groupi_n_2224 ,in1[9] ,in2[9]);
  xnor csa_tree_add_51_79_groupi_g44192(csa_tree_add_51_79_groupi_n_2223 ,in7[2] ,in8[3]);
  xnor csa_tree_add_51_79_groupi_g44193(csa_tree_add_51_79_groupi_n_2222 ,in9[2] ,in10[9]);
  xnor csa_tree_add_51_79_groupi_g44194(csa_tree_add_51_79_groupi_n_2221 ,in23[1] ,in24[9]);
  xnor csa_tree_add_51_79_groupi_g44195(csa_tree_add_51_79_groupi_n_2220 ,in17[2] ,in18[9]);
  xnor csa_tree_add_51_79_groupi_g44196(csa_tree_add_51_79_groupi_n_2219 ,in1[1] ,in2[9]);
  xnor csa_tree_add_51_79_groupi_g44197(csa_tree_add_51_79_groupi_n_2218 ,in11[3] ,in12[9]);
  xnor csa_tree_add_51_79_groupi_g44198(csa_tree_add_51_79_groupi_n_2217 ,in3[7] ,in4[9]);
  xnor csa_tree_add_51_79_groupi_g44199(csa_tree_add_51_79_groupi_n_2216 ,in7[5] ,in8[9]);
  xnor csa_tree_add_51_79_groupi_g44200(csa_tree_add_51_79_groupi_n_2215 ,in15[4] ,in16[9]);
  xnor csa_tree_add_51_79_groupi_g44201(csa_tree_add_51_79_groupi_n_2214 ,in19[9] ,in20[1]);
  xnor csa_tree_add_51_79_groupi_g44202(csa_tree_add_51_79_groupi_n_2213 ,in23[2] ,in24[9]);
  xnor csa_tree_add_51_79_groupi_g44203(csa_tree_add_51_79_groupi_n_2212 ,in23[3] ,in24[9]);
  xnor csa_tree_add_51_79_groupi_g44204(csa_tree_add_51_79_groupi_n_2211 ,in3[5] ,in4[9]);
  xnor csa_tree_add_51_79_groupi_g44205(csa_tree_add_51_79_groupi_n_2210 ,in3[9] ,in4[9]);
  xnor csa_tree_add_51_79_groupi_g44206(csa_tree_add_51_79_groupi_n_2209 ,in19[6] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g44207(csa_tree_add_51_79_groupi_n_2208 ,in21[2] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g44208(csa_tree_add_51_79_groupi_n_2207 ,in7[6] ,in8[9]);
  xnor csa_tree_add_51_79_groupi_g44209(csa_tree_add_51_79_groupi_n_2206 ,in23[8] ,in24[9]);
  xnor csa_tree_add_51_79_groupi_g44210(csa_tree_add_51_79_groupi_n_2205 ,in17[5] ,in18[9]);
  xnor csa_tree_add_51_79_groupi_g44211(csa_tree_add_51_79_groupi_n_2204 ,in5[5] ,in6[9]);
  xnor csa_tree_add_51_79_groupi_g44212(csa_tree_add_51_79_groupi_n_2203 ,in11[7] ,in12[9]);
  xnor csa_tree_add_51_79_groupi_g44213(csa_tree_add_51_79_groupi_n_2201 ,csa_tree_add_51_79_groupi_n_1624 ,in1[10]);
  xnor csa_tree_add_51_79_groupi_g44214(csa_tree_add_51_79_groupi_n_2200 ,in21[9] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g44215(csa_tree_add_51_79_groupi_n_2199 ,in5[9] ,in6[9]);
  xnor csa_tree_add_51_79_groupi_g44216(csa_tree_add_51_79_groupi_n_2198 ,in19[6] ,in20[5]);
  xnor csa_tree_add_51_79_groupi_g44217(csa_tree_add_51_79_groupi_n_2197 ,in17[7] ,in18[9]);
  xnor csa_tree_add_51_79_groupi_g44218(csa_tree_add_51_79_groupi_n_2196 ,in5[1] ,in6[9]);
  xnor csa_tree_add_51_79_groupi_g44219(csa_tree_add_51_79_groupi_n_2195 ,in19[7] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g44220(csa_tree_add_51_79_groupi_n_2194 ,in15[3] ,in16[9]);
  xnor csa_tree_add_51_79_groupi_g44221(csa_tree_add_51_79_groupi_n_2193 ,in17[4] ,in18[9]);
  xnor csa_tree_add_51_79_groupi_g44222(csa_tree_add_51_79_groupi_n_2192 ,in3[3] ,in4[7]);
  xnor csa_tree_add_51_79_groupi_g44223(csa_tree_add_51_79_groupi_n_2191 ,in1[5] ,in2[9]);
  xnor csa_tree_add_51_79_groupi_g44224(csa_tree_add_51_79_groupi_n_2190 ,in19[8] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g44225(csa_tree_add_51_79_groupi_n_2189 ,in7[1] ,in8[9]);
  xnor csa_tree_add_51_79_groupi_g44226(csa_tree_add_51_79_groupi_n_2188 ,in9[3] ,in10[9]);
  xnor csa_tree_add_51_79_groupi_g44227(csa_tree_add_51_79_groupi_n_2187 ,in9[1] ,in10[9]);
  xnor csa_tree_add_51_79_groupi_g44228(csa_tree_add_51_79_groupi_n_2186 ,in11[5] ,in12[9]);
  xnor csa_tree_add_51_79_groupi_g44229(csa_tree_add_51_79_groupi_n_2185 ,in19[8] ,in20[7]);
  xnor csa_tree_add_51_79_groupi_g44230(csa_tree_add_51_79_groupi_n_2184 ,in21[7] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g44231(csa_tree_add_51_79_groupi_n_2183 ,in19[2] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g44232(csa_tree_add_51_79_groupi_n_2182 ,in21[3] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g44233(csa_tree_add_51_79_groupi_n_2181 ,in23[6] ,in24[9]);
  xnor csa_tree_add_51_79_groupi_g44234(csa_tree_add_51_79_groupi_n_2180 ,in11[8] ,in12[9]);
  xnor csa_tree_add_51_79_groupi_g44235(csa_tree_add_51_79_groupi_n_2179 ,in21[1] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g44236(csa_tree_add_51_79_groupi_n_2178 ,in23[7] ,in24[9]);
  xnor csa_tree_add_51_79_groupi_g44237(csa_tree_add_51_79_groupi_n_2177 ,in13[1] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g44238(csa_tree_add_51_79_groupi_n_2176 ,in5[2] ,in6[9]);
  xnor csa_tree_add_51_79_groupi_g44239(csa_tree_add_51_79_groupi_n_2174 ,csa_tree_add_51_79_groupi_n_1626 ,in5[10]);
  xnor csa_tree_add_51_79_groupi_g44240(csa_tree_add_51_79_groupi_n_2173 ,in19[9] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g44241(csa_tree_add_51_79_groupi_n_2172 ,in17[10] ,in18[9]);
  xnor csa_tree_add_51_79_groupi_g44242(csa_tree_add_51_79_groupi_n_2171 ,in11[2] ,in12[9]);
  xnor csa_tree_add_51_79_groupi_g44243(csa_tree_add_51_79_groupi_n_2170 ,in11[2] ,in12[1]);
  xnor csa_tree_add_51_79_groupi_g44244(csa_tree_add_51_79_groupi_n_2169 ,in13[8] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g44245(csa_tree_add_51_79_groupi_n_2168 ,in21[10] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g44246(csa_tree_add_51_79_groupi_n_2166 ,csa_tree_add_51_79_groupi_n_1623 ,in9[10]);
  xnor csa_tree_add_51_79_groupi_g44247(csa_tree_add_51_79_groupi_n_2165 ,in3[3] ,in4[9]);
  xnor csa_tree_add_51_79_groupi_g44248(csa_tree_add_51_79_groupi_n_2164 ,in5[4] ,in6[9]);
  xnor csa_tree_add_51_79_groupi_g44249(csa_tree_add_51_79_groupi_n_2163 ,in1[2] ,in2[9]);
  xnor csa_tree_add_51_79_groupi_g44250(csa_tree_add_51_79_groupi_n_2162 ,in7[7] ,in8[9]);
  xnor csa_tree_add_51_79_groupi_g44251(csa_tree_add_51_79_groupi_n_2161 ,in5[3] ,in6[9]);
  xnor csa_tree_add_51_79_groupi_g44252(csa_tree_add_51_79_groupi_n_2160 ,in5[6] ,in6[9]);
  xnor csa_tree_add_51_79_groupi_g44253(csa_tree_add_51_79_groupi_n_2159 ,in3[1] ,in4[9]);
  xnor csa_tree_add_51_79_groupi_g44254(csa_tree_add_51_79_groupi_n_2158 ,in3[8] ,in4[9]);
  xnor csa_tree_add_51_79_groupi_g44255(csa_tree_add_51_79_groupi_n_2157 ,in19[5] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g44256(csa_tree_add_51_79_groupi_n_2156 ,in9[4] ,in10[9]);
  xnor csa_tree_add_51_79_groupi_g44257(csa_tree_add_51_79_groupi_n_2155 ,in21[10] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g44258(csa_tree_add_51_79_groupi_n_2154 ,in9[5] ,in10[9]);
  xnor csa_tree_add_51_79_groupi_g44259(csa_tree_add_51_79_groupi_n_2153 ,in15[2] ,in16[9]);
  xnor csa_tree_add_51_79_groupi_g44260(csa_tree_add_51_79_groupi_n_2152 ,in15[9] ,in16[9]);
  xnor csa_tree_add_51_79_groupi_g44261(csa_tree_add_51_79_groupi_n_2151 ,in13[2] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g44262(csa_tree_add_51_79_groupi_n_2150 ,in23[5] ,in24[7]);
  xnor csa_tree_add_51_79_groupi_g44263(csa_tree_add_51_79_groupi_n_2149 ,in17[6] ,in18[9]);
  xnor csa_tree_add_51_79_groupi_g44264(csa_tree_add_51_79_groupi_n_2148 ,in13[9] ,in14[9]);
  xnor csa_tree_add_51_79_groupi_g44265(csa_tree_add_51_79_groupi_n_2146 ,csa_tree_add_51_79_groupi_n_1557 ,in3[10]);
  xnor csa_tree_add_51_79_groupi_g44266(csa_tree_add_51_79_groupi_n_2145 ,in1[9] ,in2[3]);
  xnor csa_tree_add_51_79_groupi_g44267(csa_tree_add_51_79_groupi_n_2144 ,in11[4] ,in12[9]);
  xnor csa_tree_add_51_79_groupi_g44268(csa_tree_add_51_79_groupi_n_2143 ,in23[4] ,in24[9]);
  xnor csa_tree_add_51_79_groupi_g44269(csa_tree_add_51_79_groupi_n_2142 ,in21[10] ,in22[5]);
  xnor csa_tree_add_51_79_groupi_g44270(csa_tree_add_51_79_groupi_n_2141 ,in11[6] ,in12[7]);
  xnor csa_tree_add_51_79_groupi_g44271(csa_tree_add_51_79_groupi_n_2140 ,in11[8] ,in12[5]);
  xnor csa_tree_add_51_79_groupi_g44272(csa_tree_add_51_79_groupi_n_2139 ,in23[6] ,in24[3]);
  xnor csa_tree_add_51_79_groupi_g44273(csa_tree_add_51_79_groupi_n_2138 ,in19[1] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g44274(csa_tree_add_51_79_groupi_n_2137 ,in1[6] ,in2[9]);
  xnor csa_tree_add_51_79_groupi_g44275(csa_tree_add_51_79_groupi_n_2136 ,in21[2] ,in22[3]);
  xnor csa_tree_add_51_79_groupi_g44276(csa_tree_add_51_79_groupi_n_2135 ,in5[8] ,in6[9]);
  xnor csa_tree_add_51_79_groupi_g44277(csa_tree_add_51_79_groupi_n_2134 ,in1[4] ,in2[9]);
  xnor csa_tree_add_51_79_groupi_g44278(csa_tree_add_51_79_groupi_n_2133 ,in3[2] ,in4[9]);
  xnor csa_tree_add_51_79_groupi_g44279(csa_tree_add_51_79_groupi_n_2132 ,in7[10] ,in8[9]);
  xnor csa_tree_add_51_79_groupi_g44280(csa_tree_add_51_79_groupi_n_2131 ,in21[5] ,in22[9]);
  xnor csa_tree_add_51_79_groupi_g44281(csa_tree_add_51_79_groupi_n_2130 ,in9[8] ,in10[9]);
  xnor csa_tree_add_51_79_groupi_g44282(csa_tree_add_51_79_groupi_n_2129 ,in11[2] ,in12[7]);
  xnor csa_tree_add_51_79_groupi_g44283(csa_tree_add_51_79_groupi_n_2128 ,in19[3] ,in20[9]);
  xnor csa_tree_add_51_79_groupi_g44284(csa_tree_add_51_79_groupi_n_2127 ,in17[2] ,in18[7]);
  xnor csa_tree_add_51_79_groupi_g44285(csa_tree_add_51_79_groupi_n_2126 ,in5[2] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g44286(csa_tree_add_51_79_groupi_n_2125 ,in7[8] ,in8[9]);
  xnor csa_tree_add_51_79_groupi_g44287(csa_tree_add_51_79_groupi_n_2124 ,in23[9] ,in24[9]);
  xnor csa_tree_add_51_79_groupi_g44288(csa_tree_add_51_79_groupi_n_2123 ,in7[2] ,in8[9]);
  xnor csa_tree_add_51_79_groupi_g44289(csa_tree_add_51_79_groupi_n_2122 ,in11[6] ,in12[9]);
  xnor csa_tree_add_51_79_groupi_g44290(csa_tree_add_51_79_groupi_n_2120 ,csa_tree_add_51_79_groupi_n_1142 ,in17[10]);
  xnor csa_tree_add_51_79_groupi_g44291(csa_tree_add_51_79_groupi_n_2119 ,in7[9] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g44292(csa_tree_add_51_79_groupi_n_2117 ,csa_tree_add_51_79_groupi_n_1543 ,in9[10]);
  xnor csa_tree_add_51_79_groupi_g44293(csa_tree_add_51_79_groupi_n_2116 ,in7[8] ,in8[5]);
  xnor csa_tree_add_51_79_groupi_g44294(csa_tree_add_51_79_groupi_n_2115 ,in17[7] ,in18[5]);
  xnor csa_tree_add_51_79_groupi_g44295(csa_tree_add_51_79_groupi_n_2114 ,in7[3] ,in8[3]);
  xnor csa_tree_add_51_79_groupi_g44296(csa_tree_add_51_79_groupi_n_2113 ,in19[3] ,in20[1]);
  xnor csa_tree_add_51_79_groupi_g44297(csa_tree_add_51_79_groupi_n_2112 ,in21[6] ,in22[3]);
  xnor csa_tree_add_51_79_groupi_g44298(csa_tree_add_51_79_groupi_n_2111 ,in5[10] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g44299(csa_tree_add_51_79_groupi_n_2110 ,in19[2] ,in20[1]);
  xnor csa_tree_add_51_79_groupi_g44300(csa_tree_add_51_79_groupi_n_2109 ,in1[8] ,in2[3]);
  xnor csa_tree_add_51_79_groupi_g44301(csa_tree_add_51_79_groupi_n_2108 ,in7[3] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g44302(csa_tree_add_51_79_groupi_n_2106 ,csa_tree_add_51_79_groupi_n_1603 ,in19[10]);
  xnor csa_tree_add_51_79_groupi_g44303(csa_tree_add_51_79_groupi_n_2105 ,in9[4] ,in10[7]);
  xnor csa_tree_add_51_79_groupi_g44304(csa_tree_add_51_79_groupi_n_2104 ,in13[8] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g44305(csa_tree_add_51_79_groupi_n_2103 ,in3[3] ,in4[5]);
  xnor csa_tree_add_51_79_groupi_g44306(csa_tree_add_51_79_groupi_n_2102 ,in9[2] ,in10[7]);
  xnor csa_tree_add_51_79_groupi_g44307(csa_tree_add_51_79_groupi_n_2100 ,csa_tree_add_51_79_groupi_n_1533 ,in5[10]);
  xnor csa_tree_add_51_79_groupi_g44308(csa_tree_add_51_79_groupi_n_2099 ,in1[8] ,in2[1]);
  xnor csa_tree_add_51_79_groupi_g44309(csa_tree_add_51_79_groupi_n_2098 ,in21[8] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g44310(csa_tree_add_51_79_groupi_n_2097 ,in7[10] ,in8[7]);
  xnor csa_tree_add_51_79_groupi_g44311(csa_tree_add_51_79_groupi_n_2096 ,in1[2] ,in2[5]);
  xnor csa_tree_add_51_79_groupi_g44312(csa_tree_add_51_79_groupi_n_2095 ,in17[8] ,in18[1]);
  xnor csa_tree_add_51_79_groupi_g44313(csa_tree_add_51_79_groupi_n_2094 ,in1[1] ,in2[7]);
  xnor csa_tree_add_51_79_groupi_g44314(csa_tree_add_51_79_groupi_n_2093 ,in7[4] ,in8[5]);
  xnor csa_tree_add_51_79_groupi_g44315(csa_tree_add_51_79_groupi_n_2092 ,in5[7] ,in6[3]);
  xnor csa_tree_add_51_79_groupi_g44316(csa_tree_add_51_79_groupi_n_2091 ,in1[3] ,in2[7]);
  xnor csa_tree_add_51_79_groupi_g44317(csa_tree_add_51_79_groupi_n_2090 ,in3[8] ,in4[3]);
  xnor csa_tree_add_51_79_groupi_g44318(csa_tree_add_51_79_groupi_n_2089 ,in15[6] ,in16[5]);
  xnor csa_tree_add_51_79_groupi_g44319(csa_tree_add_51_79_groupi_n_2088 ,in5[1] ,in6[3]);
  xnor csa_tree_add_51_79_groupi_g44320(csa_tree_add_51_79_groupi_n_2087 ,in15[1] ,in16[5]);
  xnor csa_tree_add_51_79_groupi_g44321(csa_tree_add_51_79_groupi_n_2086 ,in5[6] ,in6[7]);
  xnor csa_tree_add_51_79_groupi_g44322(csa_tree_add_51_79_groupi_n_2085 ,in13[7] ,in14[3]);
  xnor csa_tree_add_51_79_groupi_g44323(csa_tree_add_51_79_groupi_n_2084 ,in15[3] ,in16[3]);
  xnor csa_tree_add_51_79_groupi_g44324(csa_tree_add_51_79_groupi_n_2083 ,in7[6] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g44325(csa_tree_add_51_79_groupi_n_2082 ,in21[5] ,in22[5]);
  xnor csa_tree_add_51_79_groupi_g44326(csa_tree_add_51_79_groupi_n_2081 ,in17[8] ,in18[7]);
  xnor csa_tree_add_51_79_groupi_g44327(csa_tree_add_51_79_groupi_n_2080 ,in9[10] ,in10[5]);
  xnor csa_tree_add_51_79_groupi_g44328(csa_tree_add_51_79_groupi_n_2079 ,in7[4] ,in8[3]);
  xnor csa_tree_add_51_79_groupi_g44329(csa_tree_add_51_79_groupi_n_2078 ,in9[6] ,in10[3]);
  xnor csa_tree_add_51_79_groupi_g44330(csa_tree_add_51_79_groupi_n_2077 ,in15[9] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g44331(csa_tree_add_51_79_groupi_n_2076 ,in21[1] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g44332(csa_tree_add_51_79_groupi_n_2075 ,in15[10] ,in16[3]);
  xnor csa_tree_add_51_79_groupi_g44333(csa_tree_add_51_79_groupi_n_2074 ,in9[9] ,in10[7]);
  xnor csa_tree_add_51_79_groupi_g44334(csa_tree_add_51_79_groupi_n_2073 ,in1[7] ,in2[1]);
  xnor csa_tree_add_51_79_groupi_g44335(csa_tree_add_51_79_groupi_n_2072 ,in5[5] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g44336(csa_tree_add_51_79_groupi_n_2071 ,in1[6] ,in2[7]);
  xnor csa_tree_add_51_79_groupi_g44337(csa_tree_add_51_79_groupi_n_2070 ,in11[7] ,in12[5]);
  xnor csa_tree_add_51_79_groupi_g44338(csa_tree_add_51_79_groupi_n_2069 ,in3[1] ,in4[7]);
  xnor csa_tree_add_51_79_groupi_g44339(csa_tree_add_51_79_groupi_n_2068 ,in1[4] ,in2[7]);
  xnor csa_tree_add_51_79_groupi_g44340(csa_tree_add_51_79_groupi_n_2067 ,in11[9] ,in12[5]);
  xnor csa_tree_add_51_79_groupi_g44341(csa_tree_add_51_79_groupi_n_2066 ,in17[4] ,in18[3]);
  xnor csa_tree_add_51_79_groupi_g44342(csa_tree_add_51_79_groupi_n_2065 ,in17[10] ,in18[5]);
  xnor csa_tree_add_51_79_groupi_g44343(csa_tree_add_51_79_groupi_n_2064 ,in19[9] ,in20[5]);
  xnor csa_tree_add_51_79_groupi_g44344(csa_tree_add_51_79_groupi_n_2063 ,in23[4] ,in24[5]);
  xnor csa_tree_add_51_79_groupi_g44345(csa_tree_add_51_79_groupi_n_2062 ,in3[4] ,in4[1]);
  xnor csa_tree_add_51_79_groupi_g44346(csa_tree_add_51_79_groupi_n_2061 ,in11[9] ,in12[1]);
  xnor csa_tree_add_51_79_groupi_g44347(csa_tree_add_51_79_groupi_n_2060 ,in13[10] ,in14[3]);
  xnor csa_tree_add_51_79_groupi_g44348(csa_tree_add_51_79_groupi_n_2059 ,in9[10] ,in10[1]);
  xnor csa_tree_add_51_79_groupi_g44349(csa_tree_add_51_79_groupi_n_2058 ,in5[9] ,in6[1]);
  xnor csa_tree_add_51_79_groupi_g44350(csa_tree_add_51_79_groupi_n_2057 ,in11[8] ,in12[7]);
  xnor csa_tree_add_51_79_groupi_g44351(csa_tree_add_51_79_groupi_n_2056 ,in23[1] ,in24[7]);
  xnor csa_tree_add_51_79_groupi_g44352(csa_tree_add_51_79_groupi_n_2055 ,in13[1] ,in14[7]);
  xnor csa_tree_add_51_79_groupi_g44353(csa_tree_add_51_79_groupi_n_2054 ,in13[9] ,in14[7]);
  xnor csa_tree_add_51_79_groupi_g44354(csa_tree_add_51_79_groupi_n_2053 ,in21[9] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g44355(csa_tree_add_51_79_groupi_n_2052 ,in15[7] ,in16[3]);
  xnor csa_tree_add_51_79_groupi_g44356(csa_tree_add_51_79_groupi_n_2051 ,in23[7] ,in24[5]);
  xnor csa_tree_add_51_79_groupi_g44357(csa_tree_add_51_79_groupi_n_2050 ,in3[4] ,in4[5]);
  xnor csa_tree_add_51_79_groupi_g44358(csa_tree_add_51_79_groupi_n_2049 ,in5[6] ,in6[5]);
  xnor csa_tree_add_51_79_groupi_g44359(csa_tree_add_51_79_groupi_n_2048 ,in1[3] ,in2[1]);
  xnor csa_tree_add_51_79_groupi_g44360(csa_tree_add_51_79_groupi_n_2047 ,in9[9] ,in10[1]);
  xnor csa_tree_add_51_79_groupi_g44361(csa_tree_add_51_79_groupi_n_2046 ,in11[10] ,in12[7]);
  xnor csa_tree_add_51_79_groupi_g44362(csa_tree_add_51_79_groupi_n_2045 ,in11[9] ,in12[7]);
  xnor csa_tree_add_51_79_groupi_g44363(csa_tree_add_51_79_groupi_n_2044 ,in13[4] ,in14[7]);
  xnor csa_tree_add_51_79_groupi_g44364(csa_tree_add_51_79_groupi_n_2043 ,in23[4] ,in24[3]);
  xnor csa_tree_add_51_79_groupi_g44365(csa_tree_add_51_79_groupi_n_2042 ,in21[4] ,in22[7]);
  xnor csa_tree_add_51_79_groupi_g44366(csa_tree_add_51_79_groupi_n_2041 ,in9[1] ,in10[3]);
  xnor csa_tree_add_51_79_groupi_g44367(csa_tree_add_51_79_groupi_n_2040 ,in1[2] ,in2[7]);
  xnor csa_tree_add_51_79_groupi_g44368(csa_tree_add_51_79_groupi_n_2039 ,in5[1] ,in6[7]);
  xnor csa_tree_add_51_79_groupi_g44369(csa_tree_add_51_79_groupi_n_2038 ,in13[7] ,in14[1]);
  xnor csa_tree_add_51_79_groupi_g44370(csa_tree_add_51_79_groupi_n_2037 ,in7[1] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g44371(csa_tree_add_51_79_groupi_n_2036 ,in9[2] ,in10[5]);
  xnor csa_tree_add_51_79_groupi_g44372(csa_tree_add_51_79_groupi_n_2035 ,in3[7] ,in4[1]);
  xnor csa_tree_add_51_79_groupi_g44373(csa_tree_add_51_79_groupi_n_2034 ,in17[6] ,in18[7]);
  xnor csa_tree_add_51_79_groupi_g44374(csa_tree_add_51_79_groupi_n_2033 ,in13[7] ,in14[7]);
  xnor csa_tree_add_51_79_groupi_g44375(csa_tree_add_51_79_groupi_n_2032 ,in19[4] ,in20[7]);
  xnor csa_tree_add_51_79_groupi_g44376(csa_tree_add_51_79_groupi_n_2031 ,in3[6] ,in4[5]);
  xnor csa_tree_add_51_79_groupi_g44377(csa_tree_add_51_79_groupi_n_2030 ,in19[1] ,in20[3]);
  xnor csa_tree_add_51_79_groupi_g44378(csa_tree_add_51_79_groupi_n_2029 ,in9[1] ,in10[1]);
  xnor csa_tree_add_51_79_groupi_g44379(csa_tree_add_51_79_groupi_n_2028 ,in3[1] ,in4[1]);
  xnor csa_tree_add_51_79_groupi_g44380(csa_tree_add_51_79_groupi_n_2027 ,in15[10] ,in16[1]);
  xnor csa_tree_add_51_79_groupi_g44381(csa_tree_add_51_79_groupi_n_2026 ,in19[7] ,in20[5]);
  xnor csa_tree_add_51_79_groupi_g44382(csa_tree_add_51_79_groupi_n_2025 ,in21[4] ,in22[1]);
  xnor csa_tree_add_51_79_groupi_g44383(csa_tree_add_51_79_groupi_n_2023 ,csa_tree_add_51_79_groupi_n_1535 ,in1[10]);
  xnor csa_tree_add_51_79_groupi_g44384(csa_tree_add_51_79_groupi_n_2022 ,in3[9] ,in4[1]);
  xnor csa_tree_add_51_79_groupi_g44385(csa_tree_add_51_79_groupi_n_2021 ,in15[1] ,in16[3]);
  xnor csa_tree_add_51_79_groupi_g44386(csa_tree_add_51_79_groupi_n_2020 ,in19[1] ,in20[7]);
  xnor csa_tree_add_51_79_groupi_g44387(csa_tree_add_51_79_groupi_n_2019 ,in9[4] ,in10[3]);
  xnor csa_tree_add_51_79_groupi_g44388(csa_tree_add_51_79_groupi_n_2018 ,in7[4] ,in8[1]);
  xnor csa_tree_add_51_79_groupi_g44389(csa_tree_add_51_79_groupi_n_2017 ,in15[7] ,in16[7]);
  xnor csa_tree_add_51_79_groupi_g44390(csa_tree_add_51_79_groupi_n_2016 ,in23[4] ,in24[1]);
  xnor csa_tree_add_51_79_groupi_g44391(csa_tree_add_51_79_groupi_n_2015 ,in1[6] ,in2[3]);
  xnor csa_tree_add_51_79_groupi_g44392(csa_tree_add_51_79_groupi_n_2012 ,csa_tree_add_51_79_groupi_n_1619 ,in8[8]);
  xnor csa_tree_add_51_79_groupi_g44393(csa_tree_add_51_79_groupi_n_2009 ,csa_tree_add_51_79_groupi_n_1532 ,in18[4]);
  xnor csa_tree_add_51_79_groupi_g44394(csa_tree_add_51_79_groupi_n_2006 ,csa_tree_add_51_79_groupi_n_1547 ,in24[6]);
  xnor csa_tree_add_51_79_groupi_g44395(csa_tree_add_51_79_groupi_n_2003 ,csa_tree_add_51_79_groupi_n_1595 ,in22[8]);
  xnor csa_tree_add_51_79_groupi_g44396(csa_tree_add_51_79_groupi_n_2000 ,csa_tree_add_51_79_groupi_n_1537 ,in10[2]);
  xnor csa_tree_add_51_79_groupi_g44397(csa_tree_add_51_79_groupi_n_1998 ,csa_tree_add_51_79_groupi_n_1599 ,in20[2]);
  xnor csa_tree_add_51_79_groupi_g44398(csa_tree_add_51_79_groupi_n_1996 ,csa_tree_add_51_79_groupi_n_1606 ,in4[2]);
  xnor csa_tree_add_51_79_groupi_g44399(csa_tree_add_51_79_groupi_n_1993 ,csa_tree_add_51_79_groupi_n_1602 ,in8[6]);
  xnor csa_tree_add_51_79_groupi_g44400(csa_tree_add_51_79_groupi_n_1991 ,csa_tree_add_51_79_groupi_n_1598 ,in4[8]);
  xnor csa_tree_add_51_79_groupi_g44401(csa_tree_add_51_79_groupi_n_1989 ,csa_tree_add_51_79_groupi_n_1618 ,in2[4]);
  xnor csa_tree_add_51_79_groupi_g44402(csa_tree_add_51_79_groupi_n_1987 ,csa_tree_add_51_79_groupi_n_1601 ,in18[2]);
  xnor csa_tree_add_51_79_groupi_g44403(csa_tree_add_51_79_groupi_n_1985 ,csa_tree_add_51_79_groupi_n_1545 ,in24[4]);
  xnor csa_tree_add_51_79_groupi_g44404(csa_tree_add_51_79_groupi_n_1983 ,csa_tree_add_51_79_groupi_n_1546 ,in16[8]);
  xnor csa_tree_add_51_79_groupi_g44405(csa_tree_add_51_79_groupi_n_1981 ,csa_tree_add_51_79_groupi_n_1609 ,in8[4]);
  xnor csa_tree_add_51_79_groupi_g44406(csa_tree_add_51_79_groupi_n_1979 ,csa_tree_add_51_79_groupi_n_1536 ,in24[8]);
  xnor csa_tree_add_51_79_groupi_g44407(csa_tree_add_51_79_groupi_n_1977 ,csa_tree_add_51_79_groupi_n_1542 ,in24[2]);
  xnor csa_tree_add_51_79_groupi_g44408(csa_tree_add_51_79_groupi_n_1974 ,csa_tree_add_51_79_groupi_n_1538 ,in16[6]);
  xnor csa_tree_add_51_79_groupi_g44409(csa_tree_add_51_79_groupi_n_1971 ,csa_tree_add_51_79_groupi_n_1600 ,in14[4]);
  xnor csa_tree_add_51_79_groupi_g44410(csa_tree_add_51_79_groupi_n_1968 ,csa_tree_add_51_79_groupi_n_1605 ,in12[6]);
  not csa_tree_add_51_79_groupi_g44411(csa_tree_add_51_79_groupi_n_1787 ,csa_tree_add_51_79_groupi_n_1786);
  not csa_tree_add_51_79_groupi_g44412(csa_tree_add_51_79_groupi_n_1785 ,csa_tree_add_51_79_groupi_n_1784);
  not csa_tree_add_51_79_groupi_g44413(csa_tree_add_51_79_groupi_n_1783 ,csa_tree_add_51_79_groupi_n_1782);
  not csa_tree_add_51_79_groupi_g44414(csa_tree_add_51_79_groupi_n_1781 ,csa_tree_add_51_79_groupi_n_1780);
  not csa_tree_add_51_79_groupi_g44415(csa_tree_add_51_79_groupi_n_1779 ,csa_tree_add_51_79_groupi_n_1778);
  and csa_tree_add_51_79_groupi_g44420(csa_tree_add_51_79_groupi_n_1773 ,in21[0] ,in22[2]);
  nor csa_tree_add_51_79_groupi_g44421(csa_tree_add_51_79_groupi_n_1772 ,in7[0] ,in8[8]);
  or csa_tree_add_51_79_groupi_g44422(csa_tree_add_51_79_groupi_n_1771 ,csa_tree_add_51_79_groupi_n_836 ,csa_tree_add_51_79_groupi_n_1662);
  nor csa_tree_add_51_79_groupi_g44423(csa_tree_add_51_79_groupi_n_1770 ,in7[0] ,in8[4]);
  or csa_tree_add_51_79_groupi_g44424(csa_tree_add_51_79_groupi_n_1769 ,csa_tree_add_51_79_groupi_n_840 ,csa_tree_add_51_79_groupi_n_1586);
  nor csa_tree_add_51_79_groupi_g44425(csa_tree_add_51_79_groupi_n_1768 ,in7[0] ,in8[2]);
  nor csa_tree_add_51_79_groupi_g44426(csa_tree_add_51_79_groupi_n_1767 ,in21[0] ,in22[2]);
  nor csa_tree_add_51_79_groupi_g44427(csa_tree_add_51_79_groupi_n_1766 ,in1[0] ,in2[8]);
  and csa_tree_add_51_79_groupi_g44428(csa_tree_add_51_79_groupi_n_1765 ,in9[0] ,in10[2]);
  and csa_tree_add_51_79_groupi_g44429(csa_tree_add_51_79_groupi_n_1764 ,in11[0] ,in12[2]);
  or csa_tree_add_51_79_groupi_g44430(csa_tree_add_51_79_groupi_n_1763 ,csa_tree_add_51_79_groupi_n_842 ,csa_tree_add_51_79_groupi_n_1581);
  or csa_tree_add_51_79_groupi_g44431(csa_tree_add_51_79_groupi_n_1762 ,csa_tree_add_51_79_groupi_n_807 ,csa_tree_add_51_79_groupi_n_1655);
  or csa_tree_add_51_79_groupi_g44432(csa_tree_add_51_79_groupi_n_1761 ,csa_tree_add_51_79_groupi_n_836 ,csa_tree_add_51_79_groupi_n_1658);
  and csa_tree_add_51_79_groupi_g44433(csa_tree_add_51_79_groupi_n_1760 ,in19[0] ,in20[2]);
  nor csa_tree_add_51_79_groupi_g44434(csa_tree_add_51_79_groupi_n_1759 ,in7[0] ,in8[6]);
  nor csa_tree_add_51_79_groupi_g44435(csa_tree_add_51_79_groupi_n_1758 ,in21[0] ,in22[4]);
  or csa_tree_add_51_79_groupi_g44436(csa_tree_add_51_79_groupi_n_1757 ,csa_tree_add_51_79_groupi_n_810 ,csa_tree_add_51_79_groupi_n_1594);
  and csa_tree_add_51_79_groupi_g44437(csa_tree_add_51_79_groupi_n_1756 ,in5[0] ,in6[2]);
  nor csa_tree_add_51_79_groupi_g44438(csa_tree_add_51_79_groupi_n_1755 ,in21[0] ,in22[8]);
  nor csa_tree_add_51_79_groupi_g44439(csa_tree_add_51_79_groupi_n_1754 ,in1[0] ,in2[6]);
  or csa_tree_add_51_79_groupi_g44440(csa_tree_add_51_79_groupi_n_1753 ,csa_tree_add_51_79_groupi_n_840 ,csa_tree_add_51_79_groupi_n_1649);
  nor csa_tree_add_51_79_groupi_g44441(csa_tree_add_51_79_groupi_n_1752 ,in19[0] ,in20[2]);
  or csa_tree_add_51_79_groupi_g44442(csa_tree_add_51_79_groupi_n_1751 ,csa_tree_add_51_79_groupi_n_848 ,csa_tree_add_51_79_groupi_n_1588);
  nor csa_tree_add_51_79_groupi_g44443(csa_tree_add_51_79_groupi_n_1750 ,in9[0] ,in10[2]);
  or csa_tree_add_51_79_groupi_g44444(csa_tree_add_51_79_groupi_n_1749 ,csa_tree_add_51_79_groupi_n_852 ,csa_tree_add_51_79_groupi_n_1651);
  and csa_tree_add_51_79_groupi_g44445(csa_tree_add_51_79_groupi_n_1748 ,in13[0] ,in14[2]);
  nor csa_tree_add_51_79_groupi_g44446(csa_tree_add_51_79_groupi_n_1747 ,in9[0] ,in10[8]);
  nor csa_tree_add_51_79_groupi_g44447(csa_tree_add_51_79_groupi_n_1746 ,in17[0] ,in18[8]);
  or csa_tree_add_51_79_groupi_g44448(csa_tree_add_51_79_groupi_n_1745 ,csa_tree_add_51_79_groupi_n_838 ,csa_tree_add_51_79_groupi_n_1657);
  or csa_tree_add_51_79_groupi_g44449(csa_tree_add_51_79_groupi_n_1744 ,csa_tree_add_51_79_groupi_n_850 ,csa_tree_add_51_79_groupi_n_1592);
  or csa_tree_add_51_79_groupi_g44450(csa_tree_add_51_79_groupi_n_1743 ,csa_tree_add_51_79_groupi_n_842 ,csa_tree_add_51_79_groupi_n_1654);
  nor csa_tree_add_51_79_groupi_g44451(csa_tree_add_51_79_groupi_n_1742 ,in11[0] ,in12[4]);
  and csa_tree_add_51_79_groupi_g44452(csa_tree_add_51_79_groupi_n_1741 ,in7[0] ,in8[2]);
  or csa_tree_add_51_79_groupi_g44453(csa_tree_add_51_79_groupi_n_1740 ,csa_tree_add_51_79_groupi_n_838 ,csa_tree_add_51_79_groupi_n_1579);
  or csa_tree_add_51_79_groupi_g44454(csa_tree_add_51_79_groupi_n_1739 ,csa_tree_add_51_79_groupi_n_844 ,csa_tree_add_51_79_groupi_n_1590);
  nor csa_tree_add_51_79_groupi_g44455(csa_tree_add_51_79_groupi_n_1738 ,in17[0] ,in18[6]);
  nor csa_tree_add_51_79_groupi_g44456(csa_tree_add_51_79_groupi_n_1737 ,in5[0] ,in6[8]);
  or csa_tree_add_51_79_groupi_g44457(csa_tree_add_51_79_groupi_n_1736 ,csa_tree_add_51_79_groupi_n_810 ,csa_tree_add_51_79_groupi_n_1652);
  nor csa_tree_add_51_79_groupi_g44458(csa_tree_add_51_79_groupi_n_1735 ,in15[0] ,in16[8]);
  or csa_tree_add_51_79_groupi_g44459(csa_tree_add_51_79_groupi_n_1734 ,csa_tree_add_51_79_groupi_n_850 ,csa_tree_add_51_79_groupi_n_1645);
  or csa_tree_add_51_79_groupi_g44460(csa_tree_add_51_79_groupi_n_1733 ,csa_tree_add_51_79_groupi_n_798 ,csa_tree_add_51_79_groupi_n_1661);
  nor csa_tree_add_51_79_groupi_g44461(csa_tree_add_51_79_groupi_n_1732 ,in3[0] ,in4[8]);
  nor csa_tree_add_51_79_groupi_g44462(csa_tree_add_51_79_groupi_n_1731 ,in1[0] ,in2[2]);
  nor csa_tree_add_51_79_groupi_g44463(csa_tree_add_51_79_groupi_n_1730 ,in15[0] ,in16[2]);
  nor csa_tree_add_51_79_groupi_g44464(csa_tree_add_51_79_groupi_n_1729 ,in15[0] ,in16[6]);
  and csa_tree_add_51_79_groupi_g44465(csa_tree_add_51_79_groupi_n_1728 ,in1[0] ,in2[2]);
  nor csa_tree_add_51_79_groupi_g44466(csa_tree_add_51_79_groupi_n_1727 ,in13[0] ,in14[8]);
  or csa_tree_add_51_79_groupi_g44467(csa_tree_add_51_79_groupi_n_1726 ,csa_tree_add_51_79_groupi_n_580 ,csa_tree_add_51_79_groupi_n_1653);
  nor csa_tree_add_51_79_groupi_g44468(csa_tree_add_51_79_groupi_n_1725 ,in19[0] ,in20[4]);
  nor csa_tree_add_51_79_groupi_g44469(csa_tree_add_51_79_groupi_n_1724 ,in15[0] ,in16[4]);
  nor csa_tree_add_51_79_groupi_g44470(csa_tree_add_51_79_groupi_n_1723 ,in5[0] ,in6[6]);
  and csa_tree_add_51_79_groupi_g44471(csa_tree_add_51_79_groupi_n_1786 ,in11[0] ,in12[0]);
  and csa_tree_add_51_79_groupi_g44472(csa_tree_add_51_79_groupi_n_1784 ,in23[0] ,in24[0]);
  and csa_tree_add_51_79_groupi_g44473(csa_tree_add_51_79_groupi_n_1782 ,in1[0] ,in2[0]);
  and csa_tree_add_51_79_groupi_g44474(csa_tree_add_51_79_groupi_n_1780 ,in7[0] ,in8[0]);
  and csa_tree_add_51_79_groupi_g44475(csa_tree_add_51_79_groupi_n_1778 ,in3[0] ,in4[0]);
  and csa_tree_add_51_79_groupi_g44476(csa_tree_add_51_79_groupi_n_1777 ,in9[0] ,in10[0]);
  and csa_tree_add_51_79_groupi_g44477(csa_tree_add_51_79_groupi_n_1776 ,in19[0] ,in20[0]);
  and csa_tree_add_51_79_groupi_g44478(csa_tree_add_51_79_groupi_n_1775 ,in13[0] ,in14[0]);
  and csa_tree_add_51_79_groupi_g44479(csa_tree_add_51_79_groupi_n_1774 ,in15[0] ,in16[0]);
  nor csa_tree_add_51_79_groupi_g44483(csa_tree_add_51_79_groupi_n_1719 ,in23[0] ,in24[8]);
  and csa_tree_add_51_79_groupi_g44484(csa_tree_add_51_79_groupi_n_1718 ,in23[0] ,in24[2]);
  nor csa_tree_add_51_79_groupi_g44485(csa_tree_add_51_79_groupi_n_1717 ,in5[0] ,in6[4]);
  or csa_tree_add_51_79_groupi_g44486(csa_tree_add_51_79_groupi_n_1716 ,csa_tree_add_51_79_groupi_n_848 ,csa_tree_add_51_79_groupi_n_1585);
  nor csa_tree_add_51_79_groupi_g44487(csa_tree_add_51_79_groupi_n_1715 ,in19[0] ,in20[8]);
  nor csa_tree_add_51_79_groupi_g44488(csa_tree_add_51_79_groupi_n_1714 ,in17[0] ,in18[4]);
  or csa_tree_add_51_79_groupi_g44489(csa_tree_add_51_79_groupi_n_1713 ,csa_tree_add_51_79_groupi_n_565 ,csa_tree_add_51_79_groupi_n_1646);
  and csa_tree_add_51_79_groupi_g44490(csa_tree_add_51_79_groupi_n_1712 ,in17[0] ,in18[2]);
  or csa_tree_add_51_79_groupi_g44491(csa_tree_add_51_79_groupi_n_1711 ,csa_tree_add_51_79_groupi_n_577 ,csa_tree_add_51_79_groupi_n_1656);
  nor csa_tree_add_51_79_groupi_g44492(csa_tree_add_51_79_groupi_n_1710 ,in11[0] ,in12[8]);
  or csa_tree_add_51_79_groupi_g44493(csa_tree_add_51_79_groupi_n_1709 ,csa_tree_add_51_79_groupi_n_583 ,csa_tree_add_51_79_groupi_n_1648);
  or csa_tree_add_51_79_groupi_g44494(csa_tree_add_51_79_groupi_n_1708 ,csa_tree_add_51_79_groupi_n_798 ,csa_tree_add_51_79_groupi_n_1593);
  or csa_tree_add_51_79_groupi_g44495(csa_tree_add_51_79_groupi_n_1707 ,csa_tree_add_51_79_groupi_n_586 ,csa_tree_add_51_79_groupi_n_1587);
  or csa_tree_add_51_79_groupi_g44496(csa_tree_add_51_79_groupi_n_1706 ,csa_tree_add_51_79_groupi_n_846 ,csa_tree_add_51_79_groupi_n_1650);
  nor csa_tree_add_51_79_groupi_g44497(csa_tree_add_51_79_groupi_n_1705 ,in11[0] ,in12[2]);
  nor csa_tree_add_51_79_groupi_g44498(csa_tree_add_51_79_groupi_n_1704 ,in23[0] ,in24[4]);
  or csa_tree_add_51_79_groupi_g44499(csa_tree_add_51_79_groupi_n_1703 ,csa_tree_add_51_79_groupi_n_807 ,csa_tree_add_51_79_groupi_n_1589);
  and csa_tree_add_51_79_groupi_g44500(csa_tree_add_51_79_groupi_n_1702 ,in3[0] ,in4[2]);
  nor csa_tree_add_51_79_groupi_g44501(csa_tree_add_51_79_groupi_n_1701 ,in5[0] ,in6[2]);
  nor csa_tree_add_51_79_groupi_g44502(csa_tree_add_51_79_groupi_n_1700 ,in19[0] ,in20[6]);
  nor csa_tree_add_51_79_groupi_g44503(csa_tree_add_51_79_groupi_n_1699 ,in13[0] ,in14[4]);
  or csa_tree_add_51_79_groupi_g44504(csa_tree_add_51_79_groupi_n_1698 ,csa_tree_add_51_79_groupi_n_846 ,csa_tree_add_51_79_groupi_n_1659);
  nor csa_tree_add_51_79_groupi_g44505(csa_tree_add_51_79_groupi_n_1697 ,in9[0] ,in10[6]);
  or csa_tree_add_51_79_groupi_g44506(csa_tree_add_51_79_groupi_n_1696 ,csa_tree_add_51_79_groupi_n_571 ,csa_tree_add_51_79_groupi_n_1647);
  or csa_tree_add_51_79_groupi_g44507(csa_tree_add_51_79_groupi_n_1695 ,csa_tree_add_51_79_groupi_n_807 ,csa_tree_add_51_79_groupi_n_1577);
  nor csa_tree_add_51_79_groupi_g44508(csa_tree_add_51_79_groupi_n_1694 ,in23[0] ,in24[2]);
  or csa_tree_add_51_79_groupi_g44509(csa_tree_add_51_79_groupi_n_1693 ,csa_tree_add_51_79_groupi_n_844 ,csa_tree_add_51_79_groupi_n_1582);
  nor csa_tree_add_51_79_groupi_g44510(csa_tree_add_51_79_groupi_n_1692 ,in1[0] ,in2[4]);
  nor csa_tree_add_51_79_groupi_g44511(csa_tree_add_51_79_groupi_n_1691 ,in21[0] ,in22[6]);
  or csa_tree_add_51_79_groupi_g44512(csa_tree_add_51_79_groupi_n_1690 ,csa_tree_add_51_79_groupi_n_852 ,csa_tree_add_51_79_groupi_n_1591);
  nor csa_tree_add_51_79_groupi_g44513(csa_tree_add_51_79_groupi_n_1689 ,in3[0] ,in4[2]);
  or csa_tree_add_51_79_groupi_g44514(csa_tree_add_51_79_groupi_n_1688 ,csa_tree_add_51_79_groupi_n_568 ,csa_tree_add_51_79_groupi_n_1583);
  nor csa_tree_add_51_79_groupi_g44515(csa_tree_add_51_79_groupi_n_1687 ,in9[0] ,in10[4]);
  or csa_tree_add_51_79_groupi_g44516(csa_tree_add_51_79_groupi_n_1686 ,csa_tree_add_51_79_groupi_n_562 ,csa_tree_add_51_79_groupi_n_1660);
  or csa_tree_add_51_79_groupi_g44517(csa_tree_add_51_79_groupi_n_1685 ,csa_tree_add_51_79_groupi_n_574 ,csa_tree_add_51_79_groupi_n_1580);
  or csa_tree_add_51_79_groupi_g44518(csa_tree_add_51_79_groupi_n_1684 ,csa_tree_add_51_79_groupi_n_810 ,csa_tree_add_51_79_groupi_n_1578);
  nor csa_tree_add_51_79_groupi_g44519(csa_tree_add_51_79_groupi_n_1683 ,in13[0] ,in14[2]);
  or csa_tree_add_51_79_groupi_g44520(csa_tree_add_51_79_groupi_n_1682 ,csa_tree_add_51_79_groupi_n_798 ,csa_tree_add_51_79_groupi_n_1584);
  nor csa_tree_add_51_79_groupi_g44521(csa_tree_add_51_79_groupi_n_1681 ,in11[0] ,in12[6]);
  nor csa_tree_add_51_79_groupi_g44522(csa_tree_add_51_79_groupi_n_1680 ,in3[0] ,in4[4]);
  nor csa_tree_add_51_79_groupi_g44523(csa_tree_add_51_79_groupi_n_1679 ,in3[0] ,in4[6]);
  nor csa_tree_add_51_79_groupi_g44524(csa_tree_add_51_79_groupi_n_1678 ,in13[0] ,in14[6]);
  nor csa_tree_add_51_79_groupi_g44525(csa_tree_add_51_79_groupi_n_1677 ,in23[0] ,in24[6]);
  nor csa_tree_add_51_79_groupi_g44526(csa_tree_add_51_79_groupi_n_1676 ,in17[0] ,in18[2]);
  and csa_tree_add_51_79_groupi_g44527(csa_tree_add_51_79_groupi_n_1675 ,in15[0] ,in16[2]);
  nor csa_tree_add_51_79_groupi_g44528(csa_tree_add_51_79_groupi_n_1674 ,csa_tree_add_51_79_groupi_n_1636 ,in14[9]);
  nor csa_tree_add_51_79_groupi_g44529(csa_tree_add_51_79_groupi_n_1673 ,csa_tree_add_51_79_groupi_n_1640 ,in18[9]);
  or csa_tree_add_51_79_groupi_g44530(csa_tree_add_51_79_groupi_n_1672 ,csa_tree_add_51_79_groupi_n_1639 ,in20[9]);
  or csa_tree_add_51_79_groupi_g44531(csa_tree_add_51_79_groupi_n_1671 ,csa_tree_add_51_79_groupi_n_1568 ,in4[9]);
  nor csa_tree_add_51_79_groupi_g44532(csa_tree_add_51_79_groupi_n_1670 ,csa_tree_add_51_79_groupi_n_1638 ,in2[9]);
  nor csa_tree_add_51_79_groupi_g44533(csa_tree_add_51_79_groupi_n_1669 ,csa_tree_add_51_79_groupi_n_1565 ,in12[9]);
  nor csa_tree_add_51_79_groupi_g44534(csa_tree_add_51_79_groupi_n_1668 ,csa_tree_add_51_79_groupi_n_1567 ,in8[9]);
  or csa_tree_add_51_79_groupi_g44535(csa_tree_add_51_79_groupi_n_1667 ,csa_tree_add_51_79_groupi_n_1633 ,in24[9]);
  nor csa_tree_add_51_79_groupi_g44536(csa_tree_add_51_79_groupi_n_1666 ,csa_tree_add_51_79_groupi_n_1634 ,in10[9]);
  nor csa_tree_add_51_79_groupi_g44537(csa_tree_add_51_79_groupi_n_1665 ,csa_tree_add_51_79_groupi_n_1637 ,in22[9]);
  nor csa_tree_add_51_79_groupi_g44538(csa_tree_add_51_79_groupi_n_1664 ,csa_tree_add_51_79_groupi_n_1566 ,in6[9]);
  nor csa_tree_add_51_79_groupi_g44539(csa_tree_add_51_79_groupi_n_1663 ,csa_tree_add_51_79_groupi_n_1635 ,in16[9]);
  and csa_tree_add_51_79_groupi_g44540(csa_tree_add_51_79_groupi_n_1722 ,in17[0] ,in18[0]);
  and csa_tree_add_51_79_groupi_g44541(csa_tree_add_51_79_groupi_n_1721 ,in21[0] ,in22[0]);
  and csa_tree_add_51_79_groupi_g44542(csa_tree_add_51_79_groupi_n_1720 ,in5[0] ,in6[0]);
  not csa_tree_add_51_79_groupi_g44543(csa_tree_add_51_79_groupi_n_1662 ,in14[8]);
  not csa_tree_add_51_79_groupi_g44544(csa_tree_add_51_79_groupi_n_1661 ,in24[6]);
  not csa_tree_add_51_79_groupi_g44545(csa_tree_add_51_79_groupi_n_1660 ,in12[4]);
  not csa_tree_add_51_79_groupi_g44546(csa_tree_add_51_79_groupi_n_1659 ,in10[4]);
  not csa_tree_add_51_79_groupi_g44547(csa_tree_add_51_79_groupi_n_1658 ,in14[4]);
  not csa_tree_add_51_79_groupi_g44548(csa_tree_add_51_79_groupi_n_1657 ,in6[6]);
  not csa_tree_add_51_79_groupi_g44549(csa_tree_add_51_79_groupi_n_1656 ,in18[4]);
  not csa_tree_add_51_79_groupi_g44550(csa_tree_add_51_79_groupi_n_1655 ,in4[4]);
  not csa_tree_add_51_79_groupi_g44551(csa_tree_add_51_79_groupi_n_1654 ,in18[8]);
  not csa_tree_add_51_79_groupi_g44552(csa_tree_add_51_79_groupi_n_1653 ,in16[4]);
  not csa_tree_add_51_79_groupi_g44553(csa_tree_add_51_79_groupi_n_1652 ,in20[8]);
  not csa_tree_add_51_79_groupi_g44554(csa_tree_add_51_79_groupi_n_1651 ,in12[8]);
  not csa_tree_add_51_79_groupi_g44555(csa_tree_add_51_79_groupi_n_1650 ,in10[6]);
  not csa_tree_add_51_79_groupi_g44556(csa_tree_add_51_79_groupi_n_1649 ,in16[6]);
  not csa_tree_add_51_79_groupi_g44557(csa_tree_add_51_79_groupi_n_1648 ,in6[8]);
  not csa_tree_add_51_79_groupi_g44558(csa_tree_add_51_79_groupi_n_1647 ,in10[8]);
  not csa_tree_add_51_79_groupi_g44559(csa_tree_add_51_79_groupi_n_1646 ,in22[4]);
  not csa_tree_add_51_79_groupi_g44560(csa_tree_add_51_79_groupi_n_1645 ,in22[8]);
  not csa_tree_add_51_79_groupi_g44561(csa_tree_add_51_79_groupi_n_1644 ,in10[0]);
  not csa_tree_add_51_79_groupi_g44562(csa_tree_add_51_79_groupi_n_1643 ,in8[0]);
  not csa_tree_add_51_79_groupi_g44563(csa_tree_add_51_79_groupi_n_1642 ,in12[0]);
  not csa_tree_add_51_79_groupi_g44564(csa_tree_add_51_79_groupi_n_1641 ,in20[0]);
  not csa_tree_add_51_79_groupi_g44565(csa_tree_add_51_79_groupi_n_1640 ,in18[10]);
  not csa_tree_add_51_79_groupi_g44566(csa_tree_add_51_79_groupi_n_1639 ,in20[10]);
  not csa_tree_add_51_79_groupi_g44567(csa_tree_add_51_79_groupi_n_1638 ,in2[10]);
  not csa_tree_add_51_79_groupi_g44568(csa_tree_add_51_79_groupi_n_1637 ,in22[10]);
  not csa_tree_add_51_79_groupi_g44569(csa_tree_add_51_79_groupi_n_1636 ,in14[10]);
  not csa_tree_add_51_79_groupi_g44570(csa_tree_add_51_79_groupi_n_1635 ,in16[10]);
  not csa_tree_add_51_79_groupi_g44571(csa_tree_add_51_79_groupi_n_1634 ,in10[10]);
  not csa_tree_add_51_79_groupi_g44572(csa_tree_add_51_79_groupi_n_1633 ,in24[10]);
  not csa_tree_add_51_79_groupi_g44573(csa_tree_add_51_79_groupi_n_1632 ,in23[0]);
  not csa_tree_add_51_79_groupi_g44574(csa_tree_add_51_79_groupi_n_1631 ,in11[0]);
  not csa_tree_add_51_79_groupi_g44575(csa_tree_add_51_79_groupi_n_1630 ,in21[0]);
  not csa_tree_add_51_79_groupi_g44576(csa_tree_add_51_79_groupi_n_1629 ,in1[0]);
  not csa_tree_add_51_79_groupi_g44577(csa_tree_add_51_79_groupi_n_1628 ,in9[0]);
  not csa_tree_add_51_79_groupi_g44578(csa_tree_add_51_79_groupi_n_1627 ,in16[9]);
  not csa_tree_add_51_79_groupi_g44579(csa_tree_add_51_79_groupi_n_1626 ,in6[9]);
  not csa_tree_add_51_79_groupi_g44580(csa_tree_add_51_79_groupi_n_1625 ,in12[9]);
  not csa_tree_add_51_79_groupi_g44581(csa_tree_add_51_79_groupi_n_1624 ,in2[9]);
  not csa_tree_add_51_79_groupi_g44582(csa_tree_add_51_79_groupi_n_1623 ,in10[9]);
  not csa_tree_add_51_79_groupi_g44583(csa_tree_add_51_79_groupi_n_1622 ,in14[9]);
  not csa_tree_add_51_79_groupi_g44584(csa_tree_add_51_79_groupi_n_1621 ,in18[9]);
  not csa_tree_add_51_79_groupi_g44585(csa_tree_add_51_79_groupi_n_1620 ,in4[5]);
  not csa_tree_add_51_79_groupi_g44586(csa_tree_add_51_79_groupi_n_1619 ,in8[7]);
  not csa_tree_add_51_79_groupi_g44587(csa_tree_add_51_79_groupi_n_1618 ,in2[3]);
  not csa_tree_add_51_79_groupi_g44588(csa_tree_add_51_79_groupi_n_1617 ,in6[1]);
  not csa_tree_add_51_79_groupi_g44589(csa_tree_add_51_79_groupi_n_1616 ,in10[5]);
  not csa_tree_add_51_79_groupi_g44590(csa_tree_add_51_79_groupi_n_1615 ,in10[3]);
  not csa_tree_add_51_79_groupi_g44591(csa_tree_add_51_79_groupi_n_1614 ,in4[3]);
  not csa_tree_add_51_79_groupi_g44592(csa_tree_add_51_79_groupi_n_1613 ,in2[7]);
  not csa_tree_add_51_79_groupi_g44593(csa_tree_add_51_79_groupi_n_1612 ,in16[1]);
  not csa_tree_add_51_79_groupi_g44594(csa_tree_add_51_79_groupi_n_1611 ,in6[5]);
  not csa_tree_add_51_79_groupi_g44595(csa_tree_add_51_79_groupi_n_1610 ,in2[1]);
  not csa_tree_add_51_79_groupi_g44596(csa_tree_add_51_79_groupi_n_1609 ,in8[3]);
  not csa_tree_add_51_79_groupi_g44597(csa_tree_add_51_79_groupi_n_1608 ,in18[5]);
  not csa_tree_add_51_79_groupi_g44598(csa_tree_add_51_79_groupi_n_1607 ,in8[1]);
  not csa_tree_add_51_79_groupi_g44599(csa_tree_add_51_79_groupi_n_1606 ,in4[1]);
  not csa_tree_add_51_79_groupi_g44600(csa_tree_add_51_79_groupi_n_1605 ,in12[5]);
  not csa_tree_add_51_79_groupi_g44601(csa_tree_add_51_79_groupi_n_1604 ,in20[7]);
  not csa_tree_add_51_79_groupi_g44602(csa_tree_add_51_79_groupi_n_1603 ,in20[3]);
  not csa_tree_add_51_79_groupi_g44603(csa_tree_add_51_79_groupi_n_1602 ,in8[5]);
  not csa_tree_add_51_79_groupi_g44604(csa_tree_add_51_79_groupi_n_1601 ,in18[1]);
  not csa_tree_add_51_79_groupi_g44605(csa_tree_add_51_79_groupi_n_1600 ,in14[3]);
  not csa_tree_add_51_79_groupi_g44606(csa_tree_add_51_79_groupi_n_1599 ,in20[1]);
  not csa_tree_add_51_79_groupi_g44607(csa_tree_add_51_79_groupi_n_1598 ,in4[7]);
  not csa_tree_add_51_79_groupi_g44608(csa_tree_add_51_79_groupi_n_1597 ,in16[3]);
  not csa_tree_add_51_79_groupi_g44609(csa_tree_add_51_79_groupi_n_1596 ,in12[7]);
  not csa_tree_add_51_79_groupi_g44610(csa_tree_add_51_79_groupi_n_1595 ,in22[7]);
  not csa_tree_add_51_79_groupi_g44611(csa_tree_add_51_79_groupi_n_1594 ,in20[6]);
  not csa_tree_add_51_79_groupi_g44612(csa_tree_add_51_79_groupi_n_1593 ,in24[4]);
  not csa_tree_add_51_79_groupi_g44613(csa_tree_add_51_79_groupi_n_1592 ,in22[6]);
  not csa_tree_add_51_79_groupi_g44614(csa_tree_add_51_79_groupi_n_1591 ,in12[6]);
  not csa_tree_add_51_79_groupi_g44615(csa_tree_add_51_79_groupi_n_1590 ,in8[4]);
  not csa_tree_add_51_79_groupi_g44616(csa_tree_add_51_79_groupi_n_1589 ,in4[6]);
  not csa_tree_add_51_79_groupi_g44617(csa_tree_add_51_79_groupi_n_1588 ,in2[6]);
  not csa_tree_add_51_79_groupi_g44618(csa_tree_add_51_79_groupi_n_1587 ,in14[6]);
  not csa_tree_add_51_79_groupi_g44619(csa_tree_add_51_79_groupi_n_1586 ,in16[8]);
  not csa_tree_add_51_79_groupi_g44620(csa_tree_add_51_79_groupi_n_1585 ,in2[8]);
  not csa_tree_add_51_79_groupi_g44621(csa_tree_add_51_79_groupi_n_1584 ,in24[8]);
  not csa_tree_add_51_79_groupi_g44622(csa_tree_add_51_79_groupi_n_1583 ,in2[4]);
  not csa_tree_add_51_79_groupi_g44623(csa_tree_add_51_79_groupi_n_1582 ,in8[6]);
  not csa_tree_add_51_79_groupi_g44624(csa_tree_add_51_79_groupi_n_1581 ,in18[6]);
  not csa_tree_add_51_79_groupi_g44625(csa_tree_add_51_79_groupi_n_1580 ,in8[8]);
  not csa_tree_add_51_79_groupi_g44626(csa_tree_add_51_79_groupi_n_1579 ,in6[4]);
  not csa_tree_add_51_79_groupi_g44627(csa_tree_add_51_79_groupi_n_1578 ,in20[4]);
  not csa_tree_add_51_79_groupi_g44628(csa_tree_add_51_79_groupi_n_1577 ,in4[8]);
  not csa_tree_add_51_79_groupi_g44629(csa_tree_add_51_79_groupi_n_1576 ,in18[0]);
  not csa_tree_add_51_79_groupi_g44630(csa_tree_add_51_79_groupi_n_1575 ,in22[0]);
  not csa_tree_add_51_79_groupi_g44631(csa_tree_add_51_79_groupi_n_1574 ,in16[0]);
  not csa_tree_add_51_79_groupi_g44632(csa_tree_add_51_79_groupi_n_1573 ,in24[0]);
  not csa_tree_add_51_79_groupi_g44633(csa_tree_add_51_79_groupi_n_1572 ,in2[0]);
  not csa_tree_add_51_79_groupi_g44634(csa_tree_add_51_79_groupi_n_1571 ,in6[0]);
  not csa_tree_add_51_79_groupi_g44635(csa_tree_add_51_79_groupi_n_1570 ,in4[0]);
  not csa_tree_add_51_79_groupi_g44636(csa_tree_add_51_79_groupi_n_1569 ,in14[0]);
  not csa_tree_add_51_79_groupi_g44637(csa_tree_add_51_79_groupi_n_1568 ,in4[10]);
  not csa_tree_add_51_79_groupi_g44638(csa_tree_add_51_79_groupi_n_1567 ,in8[10]);
  not csa_tree_add_51_79_groupi_g44639(csa_tree_add_51_79_groupi_n_1566 ,in6[10]);
  not csa_tree_add_51_79_groupi_g44640(csa_tree_add_51_79_groupi_n_1565 ,in12[10]);
  not csa_tree_add_51_79_groupi_g44641(csa_tree_add_51_79_groupi_n_1564 ,in7[0]);
  not csa_tree_add_51_79_groupi_g44642(csa_tree_add_51_79_groupi_n_1563 ,in17[0]);
  not csa_tree_add_51_79_groupi_g44643(csa_tree_add_51_79_groupi_n_1562 ,in13[0]);
  not csa_tree_add_51_79_groupi_g44644(csa_tree_add_51_79_groupi_n_1561 ,in3[0]);
  not csa_tree_add_51_79_groupi_g44645(csa_tree_add_51_79_groupi_n_1560 ,in15[0]);
  not csa_tree_add_51_79_groupi_g44646(csa_tree_add_51_79_groupi_n_1559 ,in19[0]);
  not csa_tree_add_51_79_groupi_g44647(csa_tree_add_51_79_groupi_n_1558 ,in5[0]);
  not csa_tree_add_51_79_groupi_g44648(csa_tree_add_51_79_groupi_n_1557 ,in4[9]);
  not csa_tree_add_51_79_groupi_g44649(csa_tree_add_51_79_groupi_n_1556 ,in22[9]);
  not csa_tree_add_51_79_groupi_g44650(csa_tree_add_51_79_groupi_n_1555 ,in8[9]);
  not csa_tree_add_51_79_groupi_g44651(csa_tree_add_51_79_groupi_n_1554 ,in20[9]);
  not csa_tree_add_51_79_groupi_g44652(csa_tree_add_51_79_groupi_n_1553 ,in24[9]);
  not csa_tree_add_51_79_groupi_g44653(csa_tree_add_51_79_groupi_n_1552 ,in12[3]);
  not csa_tree_add_51_79_groupi_g44654(csa_tree_add_51_79_groupi_n_1551 ,in18[7]);
  not csa_tree_add_51_79_groupi_g44655(csa_tree_add_51_79_groupi_n_1550 ,in14[1]);
  not csa_tree_add_51_79_groupi_g44656(csa_tree_add_51_79_groupi_n_1549 ,in14[5]);
  not csa_tree_add_51_79_groupi_g44657(csa_tree_add_51_79_groupi_n_1548 ,in14[7]);
  not csa_tree_add_51_79_groupi_g44658(csa_tree_add_51_79_groupi_n_1547 ,in24[5]);
  not csa_tree_add_51_79_groupi_g44659(csa_tree_add_51_79_groupi_n_1546 ,in16[7]);
  not csa_tree_add_51_79_groupi_g44660(csa_tree_add_51_79_groupi_n_1545 ,in24[3]);
  not csa_tree_add_51_79_groupi_g44661(csa_tree_add_51_79_groupi_n_1544 ,in6[7]);
  not csa_tree_add_51_79_groupi_g44662(csa_tree_add_51_79_groupi_n_1543 ,in10[7]);
  not csa_tree_add_51_79_groupi_g44663(csa_tree_add_51_79_groupi_n_1542 ,in24[1]);
  not csa_tree_add_51_79_groupi_g44664(csa_tree_add_51_79_groupi_n_1541 ,in22[3]);
  not csa_tree_add_51_79_groupi_g44665(csa_tree_add_51_79_groupi_n_1540 ,in12[1]);
  not csa_tree_add_51_79_groupi_g44666(csa_tree_add_51_79_groupi_n_1539 ,in22[1]);
  not csa_tree_add_51_79_groupi_g44667(csa_tree_add_51_79_groupi_n_1538 ,in16[5]);
  not csa_tree_add_51_79_groupi_g44668(csa_tree_add_51_79_groupi_n_1537 ,in10[1]);
  not csa_tree_add_51_79_groupi_g44669(csa_tree_add_51_79_groupi_n_1536 ,in24[7]);
  not csa_tree_add_51_79_groupi_g44670(csa_tree_add_51_79_groupi_n_1535 ,in2[5]);
  not csa_tree_add_51_79_groupi_g44671(csa_tree_add_51_79_groupi_n_1534 ,in20[5]);
  not csa_tree_add_51_79_groupi_g44672(csa_tree_add_51_79_groupi_n_1533 ,in6[3]);
  not csa_tree_add_51_79_groupi_g44673(csa_tree_add_51_79_groupi_n_1532 ,in18[3]);
  not csa_tree_add_51_79_groupi_g44674(csa_tree_add_51_79_groupi_n_1531 ,in22[5]);
  not csa_tree_add_51_79_groupi_drc_bufs45199(csa_tree_add_51_79_groupi_n_1471 ,csa_tree_add_51_79_groupi_n_1470);
  not csa_tree_add_51_79_groupi_drc_bufs45200(csa_tree_add_51_79_groupi_n_1470 ,csa_tree_add_51_79_groupi_n_2536);
  not csa_tree_add_51_79_groupi_drc_bufs45203(csa_tree_add_51_79_groupi_n_1469 ,csa_tree_add_51_79_groupi_n_1468);
  not csa_tree_add_51_79_groupi_drc_bufs45204(csa_tree_add_51_79_groupi_n_1468 ,csa_tree_add_51_79_groupi_n_2533);
  not csa_tree_add_51_79_groupi_drc_bufs45207(csa_tree_add_51_79_groupi_n_1467 ,csa_tree_add_51_79_groupi_n_1466);
  not csa_tree_add_51_79_groupi_drc_bufs45208(csa_tree_add_51_79_groupi_n_1466 ,csa_tree_add_51_79_groupi_n_2529);
  not csa_tree_add_51_79_groupi_drc_bufs45226(csa_tree_add_51_79_groupi_n_1462 ,csa_tree_add_51_79_groupi_n_1460);
  not csa_tree_add_51_79_groupi_drc_bufs45228(csa_tree_add_51_79_groupi_n_1460 ,csa_tree_add_51_79_groupi_n_1524);
  not csa_tree_add_51_79_groupi_drc_bufs45230(csa_tree_add_51_79_groupi_n_1459 ,csa_tree_add_51_79_groupi_n_1457);
  not csa_tree_add_51_79_groupi_drc_bufs45232(csa_tree_add_51_79_groupi_n_1457 ,csa_tree_add_51_79_groupi_n_1521);
  not csa_tree_add_51_79_groupi_drc_bufs45234(csa_tree_add_51_79_groupi_n_1456 ,csa_tree_add_51_79_groupi_n_1454);
  not csa_tree_add_51_79_groupi_drc_bufs45236(csa_tree_add_51_79_groupi_n_1454 ,csa_tree_add_51_79_groupi_n_2522);
  not csa_tree_add_51_79_groupi_drc_bufs45242(csa_tree_add_51_79_groupi_n_1450 ,csa_tree_add_51_79_groupi_n_1448);
  not csa_tree_add_51_79_groupi_drc_bufs45244(csa_tree_add_51_79_groupi_n_1448 ,csa_tree_add_51_79_groupi_n_2513);
  not csa_tree_add_51_79_groupi_drc_bufs45250(csa_tree_add_51_79_groupi_n_1444 ,csa_tree_add_51_79_groupi_n_1442);
  not csa_tree_add_51_79_groupi_drc_bufs45252(csa_tree_add_51_79_groupi_n_1442 ,csa_tree_add_51_79_groupi_n_1995);
  not csa_tree_add_51_79_groupi_drc_bufs45254(csa_tree_add_51_79_groupi_n_1441 ,csa_tree_add_51_79_groupi_n_1439);
  not csa_tree_add_51_79_groupi_drc_bufs45256(csa_tree_add_51_79_groupi_n_1439 ,csa_tree_add_51_79_groupi_n_1393);
  not csa_tree_add_51_79_groupi_drc_bufs45258(csa_tree_add_51_79_groupi_n_1438 ,csa_tree_add_51_79_groupi_n_1436);
  not csa_tree_add_51_79_groupi_drc_bufs45260(csa_tree_add_51_79_groupi_n_1436 ,csa_tree_add_51_79_groupi_n_2486);
  not csa_tree_add_51_79_groupi_drc_bufs45262(csa_tree_add_51_79_groupi_n_1435 ,csa_tree_add_51_79_groupi_n_1433);
  not csa_tree_add_51_79_groupi_drc_bufs45264(csa_tree_add_51_79_groupi_n_1433 ,csa_tree_add_51_79_groupi_n_1429);
  not csa_tree_add_51_79_groupi_drc_bufs45266(csa_tree_add_51_79_groupi_n_1432 ,csa_tree_add_51_79_groupi_n_1430);
  not csa_tree_add_51_79_groupi_drc_bufs45268(csa_tree_add_51_79_groupi_n_1430 ,csa_tree_add_51_79_groupi_n_1273);
  not csa_tree_add_51_79_groupi_drc_bufs45270(csa_tree_add_51_79_groupi_n_1429 ,csa_tree_add_51_79_groupi_n_1427);
  not csa_tree_add_51_79_groupi_drc_bufs45272(csa_tree_add_51_79_groupi_n_1427 ,csa_tree_add_51_79_groupi_n_2500);
  not csa_tree_add_51_79_groupi_drc_bufs45274(csa_tree_add_51_79_groupi_n_1426 ,csa_tree_add_51_79_groupi_n_1424);
  not csa_tree_add_51_79_groupi_drc_bufs45276(csa_tree_add_51_79_groupi_n_1424 ,csa_tree_add_51_79_groupi_n_1417);
  not csa_tree_add_51_79_groupi_drc_bufs45278(csa_tree_add_51_79_groupi_n_1423 ,csa_tree_add_51_79_groupi_n_1421);
  not csa_tree_add_51_79_groupi_drc_bufs45280(csa_tree_add_51_79_groupi_n_1421 ,csa_tree_add_51_79_groupi_n_1420);
  not csa_tree_add_51_79_groupi_drc_bufs45282(csa_tree_add_51_79_groupi_n_1420 ,csa_tree_add_51_79_groupi_n_1418);
  not csa_tree_add_51_79_groupi_drc_bufs45284(csa_tree_add_51_79_groupi_n_1418 ,csa_tree_add_51_79_groupi_n_1976);
  not csa_tree_add_51_79_groupi_drc_bufs45286(csa_tree_add_51_79_groupi_n_1417 ,csa_tree_add_51_79_groupi_n_1415);
  not csa_tree_add_51_79_groupi_drc_bufs45288(csa_tree_add_51_79_groupi_n_1415 ,csa_tree_add_51_79_groupi_n_2497);
  not csa_tree_add_51_79_groupi_drc_bufs45290(csa_tree_add_51_79_groupi_n_1414 ,csa_tree_add_51_79_groupi_n_1412);
  not csa_tree_add_51_79_groupi_drc_bufs45292(csa_tree_add_51_79_groupi_n_1412 ,csa_tree_add_51_79_groupi_n_1402);
  not csa_tree_add_51_79_groupi_drc_bufs45294(csa_tree_add_51_79_groupi_n_1411 ,csa_tree_add_51_79_groupi_n_1409);
  not csa_tree_add_51_79_groupi_drc_bufs45296(csa_tree_add_51_79_groupi_n_1409 ,csa_tree_add_51_79_groupi_n_1973);
  not csa_tree_add_51_79_groupi_drc_bufs45298(csa_tree_add_51_79_groupi_n_1408 ,csa_tree_add_51_79_groupi_n_1406);
  not csa_tree_add_51_79_groupi_drc_bufs45300(csa_tree_add_51_79_groupi_n_1406 ,csa_tree_add_51_79_groupi_n_1405);
  not csa_tree_add_51_79_groupi_drc_bufs45302(csa_tree_add_51_79_groupi_n_1405 ,csa_tree_add_51_79_groupi_n_1403);
  not csa_tree_add_51_79_groupi_drc_bufs45304(csa_tree_add_51_79_groupi_n_1403 ,csa_tree_add_51_79_groupi_n_1970);
  not csa_tree_add_51_79_groupi_drc_bufs45306(csa_tree_add_51_79_groupi_n_1402 ,csa_tree_add_51_79_groupi_n_1400);
  not csa_tree_add_51_79_groupi_drc_bufs45308(csa_tree_add_51_79_groupi_n_1400 ,csa_tree_add_51_79_groupi_n_2494);
  not csa_tree_add_51_79_groupi_drc_bufs45310(csa_tree_add_51_79_groupi_n_1399 ,csa_tree_add_51_79_groupi_n_1397);
  not csa_tree_add_51_79_groupi_drc_bufs45312(csa_tree_add_51_79_groupi_n_1397 ,csa_tree_add_51_79_groupi_n_1366);
  not csa_tree_add_51_79_groupi_drc_bufs45314(csa_tree_add_51_79_groupi_n_1396 ,csa_tree_add_51_79_groupi_n_1394);
  not csa_tree_add_51_79_groupi_drc_bufs45316(csa_tree_add_51_79_groupi_n_1394 ,csa_tree_add_51_79_groupi_n_1411);
  not csa_tree_add_51_79_groupi_drc_bufs45318(csa_tree_add_51_79_groupi_n_1393 ,csa_tree_add_51_79_groupi_n_1391);
  not csa_tree_add_51_79_groupi_drc_bufs45320(csa_tree_add_51_79_groupi_n_1391 ,csa_tree_add_51_79_groupi_n_2505);
  not csa_tree_add_51_79_groupi_drc_bufs45322(csa_tree_add_51_79_groupi_n_1390 ,csa_tree_add_51_79_groupi_n_1388);
  not csa_tree_add_51_79_groupi_drc_bufs45324(csa_tree_add_51_79_groupi_n_1388 ,csa_tree_add_51_79_groupi_n_2483);
  not csa_tree_add_51_79_groupi_drc_bufs45326(csa_tree_add_51_79_groupi_n_1387 ,csa_tree_add_51_79_groupi_n_1385);
  not csa_tree_add_51_79_groupi_drc_bufs45328(csa_tree_add_51_79_groupi_n_1385 ,csa_tree_add_51_79_groupi_n_1384);
  not csa_tree_add_51_79_groupi_drc_bufs45330(csa_tree_add_51_79_groupi_n_1384 ,csa_tree_add_51_79_groupi_n_1382);
  not csa_tree_add_51_79_groupi_drc_bufs45332(csa_tree_add_51_79_groupi_n_1382 ,csa_tree_add_51_79_groupi_n_2478);
  not csa_tree_add_51_79_groupi_drc_bufs45334(csa_tree_add_51_79_groupi_n_1381 ,csa_tree_add_51_79_groupi_n_1379);
  not csa_tree_add_51_79_groupi_drc_bufs45336(csa_tree_add_51_79_groupi_n_1379 ,csa_tree_add_51_79_groupi_n_1438);
  not csa_tree_add_51_79_groupi_drc_bufs45338(csa_tree_add_51_79_groupi_n_1378 ,csa_tree_add_51_79_groupi_n_1376);
  not csa_tree_add_51_79_groupi_drc_bufs45340(csa_tree_add_51_79_groupi_n_1376 ,csa_tree_add_51_79_groupi_n_1375);
  not csa_tree_add_51_79_groupi_drc_bufs45342(csa_tree_add_51_79_groupi_n_1375 ,csa_tree_add_51_79_groupi_n_1373);
  not csa_tree_add_51_79_groupi_drc_bufs45344(csa_tree_add_51_79_groupi_n_1373 ,csa_tree_add_51_79_groupi_n_2475);
  not csa_tree_add_51_79_groupi_drc_bufs45346(csa_tree_add_51_79_groupi_n_1372 ,csa_tree_add_51_79_groupi_n_1370);
  not csa_tree_add_51_79_groupi_drc_bufs45348(csa_tree_add_51_79_groupi_n_1370 ,csa_tree_add_51_79_groupi_n_1369);
  not csa_tree_add_51_79_groupi_drc_bufs45350(csa_tree_add_51_79_groupi_n_1369 ,csa_tree_add_51_79_groupi_n_1367);
  not csa_tree_add_51_79_groupi_drc_bufs45352(csa_tree_add_51_79_groupi_n_1367 ,csa_tree_add_51_79_groupi_n_2472);
  not csa_tree_add_51_79_groupi_drc_bufs45354(csa_tree_add_51_79_groupi_n_1366 ,csa_tree_add_51_79_groupi_n_1364);
  not csa_tree_add_51_79_groupi_drc_bufs45356(csa_tree_add_51_79_groupi_n_1364 ,csa_tree_add_51_79_groupi_n_2491);
  not csa_tree_add_51_79_groupi_drc_bufs45358(csa_tree_add_51_79_groupi_n_1363 ,csa_tree_add_51_79_groupi_n_1361);
  not csa_tree_add_51_79_groupi_drc_bufs45360(csa_tree_add_51_79_groupi_n_1361 ,csa_tree_add_51_79_groupi_n_1360);
  not csa_tree_add_51_79_groupi_drc_bufs45362(csa_tree_add_51_79_groupi_n_1360 ,csa_tree_add_51_79_groupi_n_1358);
  not csa_tree_add_51_79_groupi_drc_bufs45364(csa_tree_add_51_79_groupi_n_1358 ,csa_tree_add_51_79_groupi_n_2469);
  not csa_tree_add_51_79_groupi_drc_bufs45366(csa_tree_add_51_79_groupi_n_1357 ,csa_tree_add_51_79_groupi_n_1355);
  not csa_tree_add_51_79_groupi_drc_bufs45368(csa_tree_add_51_79_groupi_n_1355 ,csa_tree_add_51_79_groupi_n_1354);
  not csa_tree_add_51_79_groupi_drc_bufs45370(csa_tree_add_51_79_groupi_n_1354 ,csa_tree_add_51_79_groupi_n_1352);
  not csa_tree_add_51_79_groupi_drc_bufs45372(csa_tree_add_51_79_groupi_n_1352 ,csa_tree_add_51_79_groupi_n_2466);
  not csa_tree_add_51_79_groupi_drc_bufs45374(csa_tree_add_51_79_groupi_n_1351 ,csa_tree_add_51_79_groupi_n_1349);
  not csa_tree_add_51_79_groupi_drc_bufs45376(csa_tree_add_51_79_groupi_n_1349 ,csa_tree_add_51_79_groupi_n_1348);
  not csa_tree_add_51_79_groupi_drc_bufs45378(csa_tree_add_51_79_groupi_n_1348 ,csa_tree_add_51_79_groupi_n_1346);
  not csa_tree_add_51_79_groupi_drc_bufs45380(csa_tree_add_51_79_groupi_n_1346 ,csa_tree_add_51_79_groupi_n_2463);
  not csa_tree_add_51_79_groupi_drc_bufs45382(csa_tree_add_51_79_groupi_n_1345 ,csa_tree_add_51_79_groupi_n_1343);
  not csa_tree_add_51_79_groupi_drc_bufs45384(csa_tree_add_51_79_groupi_n_1343 ,csa_tree_add_51_79_groupi_n_1342);
  not csa_tree_add_51_79_groupi_drc_bufs45386(csa_tree_add_51_79_groupi_n_1342 ,csa_tree_add_51_79_groupi_n_1340);
  not csa_tree_add_51_79_groupi_drc_bufs45388(csa_tree_add_51_79_groupi_n_1340 ,csa_tree_add_51_79_groupi_n_2460);
  not csa_tree_add_51_79_groupi_drc_bufs45390(csa_tree_add_51_79_groupi_n_1339 ,csa_tree_add_51_79_groupi_n_1337);
  not csa_tree_add_51_79_groupi_drc_bufs45392(csa_tree_add_51_79_groupi_n_1337 ,csa_tree_add_51_79_groupi_n_1336);
  not csa_tree_add_51_79_groupi_drc_bufs45394(csa_tree_add_51_79_groupi_n_1336 ,csa_tree_add_51_79_groupi_n_1334);
  not csa_tree_add_51_79_groupi_drc_bufs45396(csa_tree_add_51_79_groupi_n_1334 ,csa_tree_add_51_79_groupi_n_2457);
  not csa_tree_add_51_79_groupi_drc_bufs45398(csa_tree_add_51_79_groupi_n_1333 ,csa_tree_add_51_79_groupi_n_1331);
  not csa_tree_add_51_79_groupi_drc_bufs45400(csa_tree_add_51_79_groupi_n_1331 ,csa_tree_add_51_79_groupi_n_1330);
  not csa_tree_add_51_79_groupi_drc_bufs45402(csa_tree_add_51_79_groupi_n_1330 ,csa_tree_add_51_79_groupi_n_1328);
  not csa_tree_add_51_79_groupi_drc_bufs45404(csa_tree_add_51_79_groupi_n_1328 ,csa_tree_add_51_79_groupi_n_2452);
  not csa_tree_add_51_79_groupi_drc_bufs45406(csa_tree_add_51_79_groupi_n_1327 ,csa_tree_add_51_79_groupi_n_1325);
  not csa_tree_add_51_79_groupi_drc_bufs45408(csa_tree_add_51_79_groupi_n_1325 ,csa_tree_add_51_79_groupi_n_1324);
  not csa_tree_add_51_79_groupi_drc_bufs45410(csa_tree_add_51_79_groupi_n_1324 ,csa_tree_add_51_79_groupi_n_1322);
  not csa_tree_add_51_79_groupi_drc_bufs45412(csa_tree_add_51_79_groupi_n_1322 ,csa_tree_add_51_79_groupi_n_2449);
  not csa_tree_add_51_79_groupi_drc_bufs45414(csa_tree_add_51_79_groupi_n_1321 ,csa_tree_add_51_79_groupi_n_1319);
  not csa_tree_add_51_79_groupi_drc_bufs45416(csa_tree_add_51_79_groupi_n_1319 ,csa_tree_add_51_79_groupi_n_1318);
  not csa_tree_add_51_79_groupi_drc_bufs45418(csa_tree_add_51_79_groupi_n_1318 ,csa_tree_add_51_79_groupi_n_1316);
  not csa_tree_add_51_79_groupi_drc_bufs45420(csa_tree_add_51_79_groupi_n_1316 ,csa_tree_add_51_79_groupi_n_2444);
  not csa_tree_add_51_79_groupi_drc_bufs45422(csa_tree_add_51_79_groupi_n_1315 ,csa_tree_add_51_79_groupi_n_1313);
  not csa_tree_add_51_79_groupi_drc_bufs45424(csa_tree_add_51_79_groupi_n_1313 ,csa_tree_add_51_79_groupi_n_1312);
  not csa_tree_add_51_79_groupi_drc_bufs45426(csa_tree_add_51_79_groupi_n_1312 ,csa_tree_add_51_79_groupi_n_1310);
  not csa_tree_add_51_79_groupi_drc_bufs45428(csa_tree_add_51_79_groupi_n_1310 ,csa_tree_add_51_79_groupi_n_2441);
  not csa_tree_add_51_79_groupi_drc_bufs45430(csa_tree_add_51_79_groupi_n_1309 ,csa_tree_add_51_79_groupi_n_1307);
  not csa_tree_add_51_79_groupi_drc_bufs45432(csa_tree_add_51_79_groupi_n_1307 ,csa_tree_add_51_79_groupi_n_1306);
  not csa_tree_add_51_79_groupi_drc_bufs45434(csa_tree_add_51_79_groupi_n_1306 ,csa_tree_add_51_79_groupi_n_1304);
  not csa_tree_add_51_79_groupi_drc_bufs45436(csa_tree_add_51_79_groupi_n_1304 ,csa_tree_add_51_79_groupi_n_2438);
  not csa_tree_add_51_79_groupi_drc_bufs45438(csa_tree_add_51_79_groupi_n_1303 ,csa_tree_add_51_79_groupi_n_1301);
  not csa_tree_add_51_79_groupi_drc_bufs45440(csa_tree_add_51_79_groupi_n_1301 ,csa_tree_add_51_79_groupi_n_1300);
  not csa_tree_add_51_79_groupi_drc_bufs45442(csa_tree_add_51_79_groupi_n_1300 ,csa_tree_add_51_79_groupi_n_1298);
  not csa_tree_add_51_79_groupi_drc_bufs45444(csa_tree_add_51_79_groupi_n_1298 ,csa_tree_add_51_79_groupi_n_2014);
  not csa_tree_add_51_79_groupi_drc_bufs45446(csa_tree_add_51_79_groupi_n_1297 ,csa_tree_add_51_79_groupi_n_1295);
  not csa_tree_add_51_79_groupi_drc_bufs45448(csa_tree_add_51_79_groupi_n_1295 ,csa_tree_add_51_79_groupi_n_1294);
  not csa_tree_add_51_79_groupi_drc_bufs45450(csa_tree_add_51_79_groupi_n_1294 ,csa_tree_add_51_79_groupi_n_1292);
  not csa_tree_add_51_79_groupi_drc_bufs45452(csa_tree_add_51_79_groupi_n_1292 ,csa_tree_add_51_79_groupi_n_2011);
  not csa_tree_add_51_79_groupi_drc_bufs45454(csa_tree_add_51_79_groupi_n_1291 ,csa_tree_add_51_79_groupi_n_1289);
  not csa_tree_add_51_79_groupi_drc_bufs45456(csa_tree_add_51_79_groupi_n_1289 ,csa_tree_add_51_79_groupi_n_1288);
  not csa_tree_add_51_79_groupi_drc_bufs45458(csa_tree_add_51_79_groupi_n_1288 ,csa_tree_add_51_79_groupi_n_1286);
  not csa_tree_add_51_79_groupi_drc_bufs45460(csa_tree_add_51_79_groupi_n_1286 ,csa_tree_add_51_79_groupi_n_2008);
  not csa_tree_add_51_79_groupi_drc_bufs45462(csa_tree_add_51_79_groupi_n_1285 ,csa_tree_add_51_79_groupi_n_1283);
  not csa_tree_add_51_79_groupi_drc_bufs45464(csa_tree_add_51_79_groupi_n_1283 ,csa_tree_add_51_79_groupi_n_1282);
  not csa_tree_add_51_79_groupi_drc_bufs45466(csa_tree_add_51_79_groupi_n_1282 ,csa_tree_add_51_79_groupi_n_1280);
  not csa_tree_add_51_79_groupi_drc_bufs45468(csa_tree_add_51_79_groupi_n_1280 ,csa_tree_add_51_79_groupi_n_2005);
  not csa_tree_add_51_79_groupi_drc_bufs45470(csa_tree_add_51_79_groupi_n_1279 ,csa_tree_add_51_79_groupi_n_1277);
  not csa_tree_add_51_79_groupi_drc_bufs45472(csa_tree_add_51_79_groupi_n_1277 ,csa_tree_add_51_79_groupi_n_1276);
  not csa_tree_add_51_79_groupi_drc_bufs45474(csa_tree_add_51_79_groupi_n_1276 ,csa_tree_add_51_79_groupi_n_1274);
  not csa_tree_add_51_79_groupi_drc_bufs45476(csa_tree_add_51_79_groupi_n_1274 ,csa_tree_add_51_79_groupi_n_2002);
  not csa_tree_add_51_79_groupi_drc_bufs45478(csa_tree_add_51_79_groupi_n_1273 ,csa_tree_add_51_79_groupi_n_1271);
  not csa_tree_add_51_79_groupi_drc_bufs45480(csa_tree_add_51_79_groupi_n_1271 ,csa_tree_add_51_79_groupi_n_2510);
  not csa_tree_add_51_79_groupi_drc_bufs45482(csa_tree_add_51_79_groupi_n_1270 ,csa_tree_add_51_79_groupi_n_1268);
  not csa_tree_add_51_79_groupi_drc_bufs45484(csa_tree_add_51_79_groupi_n_1268 ,csa_tree_add_51_79_groupi_n_1390);
  not csa_tree_add_51_79_groupi_drc_bufs45486(csa_tree_add_51_79_groupi_n_1267 ,csa_tree_add_51_79_groupi_n_1265);
  not csa_tree_add_51_79_groupi_drc_bufs45488(csa_tree_add_51_79_groupi_n_1265 ,csa_tree_add_51_79_groupi_n_1444);
  not csa_tree_add_51_79_groupi_drc_bufs45490(csa_tree_add_51_79_groupi_n_1264 ,csa_tree_add_51_79_groupi_n_1262);
  not csa_tree_add_51_79_groupi_drc_bufs45492(csa_tree_add_51_79_groupi_n_1262 ,csa_tree_add_51_79_groupi_n_1484);
  not csa_tree_add_51_79_groupi_drc_bufs45494(csa_tree_add_51_79_groupi_n_1261 ,csa_tree_add_51_79_groupi_n_1259);
  not csa_tree_add_51_79_groupi_drc_bufs45496(csa_tree_add_51_79_groupi_n_1259 ,csa_tree_add_51_79_groupi_n_1517);
  not csa_tree_add_51_79_groupi_drc_bufs45498(csa_tree_add_51_79_groupi_n_1258 ,csa_tree_add_51_79_groupi_n_1256);
  not csa_tree_add_51_79_groupi_drc_bufs45500(csa_tree_add_51_79_groupi_n_1256 ,csa_tree_add_51_79_groupi_n_1482);
  not csa_tree_add_51_79_groupi_drc_bufs45502(csa_tree_add_51_79_groupi_n_1255 ,csa_tree_add_51_79_groupi_n_1253);
  not csa_tree_add_51_79_groupi_drc_bufs45504(csa_tree_add_51_79_groupi_n_1253 ,csa_tree_add_51_79_groupi_n_1480);
  not csa_tree_add_51_79_groupi_drc_bufs45506(csa_tree_add_51_79_groupi_n_1252 ,csa_tree_add_51_79_groupi_n_1250);
  not csa_tree_add_51_79_groupi_drc_bufs45508(csa_tree_add_51_79_groupi_n_1250 ,csa_tree_add_51_79_groupi_n_1479);
  not csa_tree_add_51_79_groupi_drc_bufs45510(csa_tree_add_51_79_groupi_n_1249 ,csa_tree_add_51_79_groupi_n_1247);
  not csa_tree_add_51_79_groupi_drc_bufs45512(csa_tree_add_51_79_groupi_n_1247 ,csa_tree_add_51_79_groupi_n_1515);
  not csa_tree_add_51_79_groupi_drc_bufs45514(csa_tree_add_51_79_groupi_n_1246 ,csa_tree_add_51_79_groupi_n_1244);
  not csa_tree_add_51_79_groupi_drc_bufs45516(csa_tree_add_51_79_groupi_n_1244 ,csa_tree_add_51_79_groupi_n_1477);
  not csa_tree_add_51_79_groupi_drc_bufs45518(csa_tree_add_51_79_groupi_n_1243 ,csa_tree_add_51_79_groupi_n_1241);
  not csa_tree_add_51_79_groupi_drc_bufs45520(csa_tree_add_51_79_groupi_n_1241 ,csa_tree_add_51_79_groupi_n_1476);
  not csa_tree_add_51_79_groupi_drc_bufs45522(csa_tree_add_51_79_groupi_n_1240 ,csa_tree_add_51_79_groupi_n_1238);
  not csa_tree_add_51_79_groupi_drc_bufs45524(csa_tree_add_51_79_groupi_n_1238 ,csa_tree_add_51_79_groupi_n_1475);
  not csa_tree_add_51_79_groupi_drc_bufs45526(csa_tree_add_51_79_groupi_n_1237 ,csa_tree_add_51_79_groupi_n_1235);
  not csa_tree_add_51_79_groupi_drc_bufs45528(csa_tree_add_51_79_groupi_n_1235 ,csa_tree_add_51_79_groupi_n_1481);
  not csa_tree_add_51_79_groupi_drc_bufs45530(csa_tree_add_51_79_groupi_n_1234 ,csa_tree_add_51_79_groupi_n_1232);
  not csa_tree_add_51_79_groupi_drc_bufs45532(csa_tree_add_51_79_groupi_n_1232 ,csa_tree_add_51_79_groupi_n_1510);
  not csa_tree_add_51_79_groupi_drc_bufs45534(csa_tree_add_51_79_groupi_n_1231 ,csa_tree_add_51_79_groupi_n_1229);
  not csa_tree_add_51_79_groupi_drc_bufs45536(csa_tree_add_51_79_groupi_n_1229 ,csa_tree_add_51_79_groupi_n_1478);
  not csa_tree_add_51_79_groupi_drc_bufs45538(csa_tree_add_51_79_groupi_n_1228 ,csa_tree_add_51_79_groupi_n_1226);
  not csa_tree_add_51_79_groupi_drc_bufs45540(csa_tree_add_51_79_groupi_n_1226 ,csa_tree_add_51_79_groupi_n_1507);
  not csa_tree_add_51_79_groupi_drc_bufs45542(csa_tree_add_51_79_groupi_n_1225 ,csa_tree_add_51_79_groupi_n_1223);
  not csa_tree_add_51_79_groupi_drc_bufs45544(csa_tree_add_51_79_groupi_n_1223 ,csa_tree_add_51_79_groupi_n_1498);
  not csa_tree_add_51_79_groupi_drc_bufs45546(csa_tree_add_51_79_groupi_n_1222 ,csa_tree_add_51_79_groupi_n_1220);
  not csa_tree_add_51_79_groupi_drc_bufs45548(csa_tree_add_51_79_groupi_n_1220 ,csa_tree_add_51_79_groupi_n_1495);
  not csa_tree_add_51_79_groupi_drc_bufs45550(csa_tree_add_51_79_groupi_n_1219 ,csa_tree_add_51_79_groupi_n_1217);
  not csa_tree_add_51_79_groupi_drc_bufs45552(csa_tree_add_51_79_groupi_n_1217 ,csa_tree_add_51_79_groupi_n_1491);
  not csa_tree_add_51_79_groupi_drc_bufs45554(csa_tree_add_51_79_groupi_n_1216 ,csa_tree_add_51_79_groupi_n_1214);
  not csa_tree_add_51_79_groupi_drc_bufs45556(csa_tree_add_51_79_groupi_n_1214 ,csa_tree_add_51_79_groupi_n_1519);
  not csa_tree_add_51_79_groupi_drc_bufs45558(csa_tree_add_51_79_groupi_n_1213 ,csa_tree_add_51_79_groupi_n_1211);
  not csa_tree_add_51_79_groupi_drc_bufs45560(csa_tree_add_51_79_groupi_n_1211 ,csa_tree_add_51_79_groupi_n_1485);
  not csa_tree_add_51_79_groupi_drc_bufs45562(csa_tree_add_51_79_groupi_n_1210 ,csa_tree_add_51_79_groupi_n_3268);
  not csa_tree_add_51_79_groupi_drc_bufs45687(csa_tree_add_51_79_groupi_n_1178 ,csa_tree_add_51_79_groupi_n_1177);
  not csa_tree_add_51_79_groupi_drc_bufs45688(csa_tree_add_51_79_groupi_n_1177 ,csa_tree_add_51_79_groupi_n_3191);
  not csa_tree_add_51_79_groupi_drc_bufs45691(csa_tree_add_51_79_groupi_n_1176 ,csa_tree_add_51_79_groupi_n_1175);
  not csa_tree_add_51_79_groupi_drc_bufs45692(csa_tree_add_51_79_groupi_n_1175 ,csa_tree_add_51_79_groupi_n_3193);
  not csa_tree_add_51_79_groupi_drc_bufs45695(csa_tree_add_51_79_groupi_n_1174 ,csa_tree_add_51_79_groupi_n_1173);
  not csa_tree_add_51_79_groupi_drc_bufs45696(csa_tree_add_51_79_groupi_n_1173 ,csa_tree_add_51_79_groupi_n_3192);
  not csa_tree_add_51_79_groupi_drc_bufs45700(csa_tree_add_51_79_groupi_n_1507 ,csa_tree_add_51_79_groupi_n_2479);
  not csa_tree_add_51_79_groupi_drc_bufs45704(csa_tree_add_51_79_groupi_n_1498 ,csa_tree_add_51_79_groupi_n_2453);
  not csa_tree_add_51_79_groupi_drc_bufs45708(csa_tree_add_51_79_groupi_n_1519 ,csa_tree_add_51_79_groupi_n_2511);
  not csa_tree_add_51_79_groupi_drc_bufs45712(csa_tree_add_51_79_groupi_n_1485 ,csa_tree_add_51_79_groupi_n_1998);
  not csa_tree_add_51_79_groupi_drc_bufs45716(csa_tree_add_51_79_groupi_n_1517 ,csa_tree_add_51_79_groupi_n_2506);
  not csa_tree_add_51_79_groupi_drc_bufs45720(csa_tree_add_51_79_groupi_n_1481 ,csa_tree_add_51_79_groupi_n_1989);
  not csa_tree_add_51_79_groupi_drc_bufs45724(csa_tree_add_51_79_groupi_n_1484 ,csa_tree_add_51_79_groupi_n_1996);
  not csa_tree_add_51_79_groupi_drc_bufs45728(csa_tree_add_51_79_groupi_n_1477 ,csa_tree_add_51_79_groupi_n_1981);
  not csa_tree_add_51_79_groupi_drc_bufs45732(csa_tree_add_51_79_groupi_n_1495 ,csa_tree_add_51_79_groupi_n_2445);
  not csa_tree_add_51_79_groupi_drc_bufs45736(csa_tree_add_51_79_groupi_n_1480 ,csa_tree_add_51_79_groupi_n_1987);
  not csa_tree_add_51_79_groupi_drc_bufs45740(csa_tree_add_51_79_groupi_n_1478 ,csa_tree_add_51_79_groupi_n_1983);
  not csa_tree_add_51_79_groupi_drc_bufs45744(csa_tree_add_51_79_groupi_n_1515 ,csa_tree_add_51_79_groupi_n_2501);
  not csa_tree_add_51_79_groupi_drc_bufs45748(csa_tree_add_51_79_groupi_n_1482 ,csa_tree_add_51_79_groupi_n_1991);
  not csa_tree_add_51_79_groupi_drc_bufs45752(csa_tree_add_51_79_groupi_n_1475 ,csa_tree_add_51_79_groupi_n_1977);
  not csa_tree_add_51_79_groupi_drc_bufs45756(csa_tree_add_51_79_groupi_n_1510 ,csa_tree_add_51_79_groupi_n_2487);
  not csa_tree_add_51_79_groupi_drc_bufs45764(csa_tree_add_51_79_groupi_n_1479 ,csa_tree_add_51_79_groupi_n_1985);
  not csa_tree_add_51_79_groupi_drc_bufs45780(csa_tree_add_51_79_groupi_n_1491 ,csa_tree_add_51_79_groupi_n_2434);
  not csa_tree_add_51_79_groupi_drc_bufs45784(csa_tree_add_51_79_groupi_n_1476 ,csa_tree_add_51_79_groupi_n_1979);
  not csa_tree_add_51_79_groupi_drc_bufs45787(csa_tree_add_51_79_groupi_n_1146 ,csa_tree_add_51_79_groupi_n_1145);
  not csa_tree_add_51_79_groupi_drc_bufs45788(csa_tree_add_51_79_groupi_n_1145 ,csa_tree_add_51_79_groupi_n_1543);
  not csa_tree_add_51_79_groupi_drc_bufs45791(csa_tree_add_51_79_groupi_n_1144 ,csa_tree_add_51_79_groupi_n_1143);
  not csa_tree_add_51_79_groupi_drc_bufs45792(csa_tree_add_51_79_groupi_n_1143 ,csa_tree_add_51_79_groupi_n_1614);
  not csa_tree_add_51_79_groupi_drc_bufs45795(csa_tree_add_51_79_groupi_n_1142 ,csa_tree_add_51_79_groupi_n_1141);
  not csa_tree_add_51_79_groupi_drc_bufs45796(csa_tree_add_51_79_groupi_n_1141 ,csa_tree_add_51_79_groupi_n_1532);
  not csa_tree_add_51_79_groupi_drc_bufs45799(csa_tree_add_51_79_groupi_n_1140 ,csa_tree_add_51_79_groupi_n_1139);
  not csa_tree_add_51_79_groupi_drc_bufs45800(csa_tree_add_51_79_groupi_n_1139 ,csa_tree_add_51_79_groupi_n_1603);
  not csa_tree_add_51_79_groupi_drc_bufs45803(csa_tree_add_51_79_groupi_n_1138 ,csa_tree_add_51_79_groupi_n_1137);
  not csa_tree_add_51_79_groupi_drc_bufs45804(csa_tree_add_51_79_groupi_n_1137 ,csa_tree_add_51_79_groupi_n_1547);
  not csa_tree_add_51_79_groupi_drc_bufs45807(csa_tree_add_51_79_groupi_n_1136 ,csa_tree_add_51_79_groupi_n_1135);
  not csa_tree_add_51_79_groupi_drc_bufs45808(csa_tree_add_51_79_groupi_n_1135 ,csa_tree_add_51_79_groupi_n_1552);
  not csa_tree_add_51_79_groupi_drc_bufs45811(csa_tree_add_51_79_groupi_n_1134 ,csa_tree_add_51_79_groupi_n_1133);
  not csa_tree_add_51_79_groupi_drc_bufs45812(csa_tree_add_51_79_groupi_n_1133 ,csa_tree_add_51_79_groupi_n_1545);
  not csa_tree_add_51_79_groupi_drc_bufs45815(csa_tree_add_51_79_groupi_n_1132 ,csa_tree_add_51_79_groupi_n_1131);
  not csa_tree_add_51_79_groupi_drc_bufs45816(csa_tree_add_51_79_groupi_n_1131 ,csa_tree_add_51_79_groupi_n_1535);
  not csa_tree_add_51_79_groupi_drc_bufs45819(csa_tree_add_51_79_groupi_n_1130 ,csa_tree_add_51_79_groupi_n_1129);
  not csa_tree_add_51_79_groupi_drc_bufs45820(csa_tree_add_51_79_groupi_n_1129 ,csa_tree_add_51_79_groupi_n_1533);
  not csa_tree_add_51_79_groupi_drc_bufs45823(csa_tree_add_51_79_groupi_n_1128 ,csa_tree_add_51_79_groupi_n_1127);
  not csa_tree_add_51_79_groupi_drc_bufs45824(csa_tree_add_51_79_groupi_n_1127 ,csa_tree_add_51_79_groupi_n_1609);
  not csa_tree_add_51_79_groupi_drc_bufs45827(csa_tree_add_51_79_groupi_n_1126 ,csa_tree_add_51_79_groupi_n_1125);
  not csa_tree_add_51_79_groupi_drc_bufs45828(csa_tree_add_51_79_groupi_n_1125 ,csa_tree_add_51_79_groupi_n_1602);
  not csa_tree_add_51_79_groupi_drc_bufs45830(csa_tree_add_51_79_groupi_n_1124 ,csa_tree_add_51_79_groupi_n_1122);
  not csa_tree_add_51_79_groupi_drc_bufs45832(csa_tree_add_51_79_groupi_n_1122 ,csa_tree_add_51_79_groupi_n_1527);
  not csa_tree_add_51_79_groupi_drc_bufs45842(csa_tree_add_51_79_groupi_n_1115 ,csa_tree_add_51_79_groupi_n_2000);
  not csa_tree_add_51_79_groupi_drc_bufs45846(csa_tree_add_51_79_groupi_n_1114 ,csa_tree_add_51_79_groupi_n_2447);
  not csa_tree_add_51_79_groupi_drc_bufs45850(csa_tree_add_51_79_groupi_n_1113 ,csa_tree_add_51_79_groupi_n_2006);
  not csa_tree_add_51_79_groupi_drc_bufs45854(csa_tree_add_51_79_groupi_n_1112 ,csa_tree_add_51_79_groupi_n_2450);
  not csa_tree_add_51_79_groupi_drc_bufs45858(csa_tree_add_51_79_groupi_n_1111 ,csa_tree_add_51_79_groupi_n_2508);
  not csa_tree_add_51_79_groupi_drc_bufs45862(csa_tree_add_51_79_groupi_n_1110 ,csa_tree_add_51_79_groupi_n_2442);
  not csa_tree_add_51_79_groupi_drc_bufs45866(csa_tree_add_51_79_groupi_n_1109 ,csa_tree_add_51_79_groupi_n_1971);
  not csa_tree_add_51_79_groupi_drc_bufs45870(csa_tree_add_51_79_groupi_n_1108 ,csa_tree_add_51_79_groupi_n_2498);
  not csa_tree_add_51_79_groupi_drc_bufs45874(csa_tree_add_51_79_groupi_n_1107 ,csa_tree_add_51_79_groupi_n_2481);
  not csa_tree_add_51_79_groupi_drc_bufs45878(csa_tree_add_51_79_groupi_n_1106 ,csa_tree_add_51_79_groupi_n_2012);
  not csa_tree_add_51_79_groupi_drc_bufs45882(csa_tree_add_51_79_groupi_n_1105 ,csa_tree_add_51_79_groupi_n_2484);
  not csa_tree_add_51_79_groupi_drc_bufs45886(csa_tree_add_51_79_groupi_n_1104 ,csa_tree_add_51_79_groupi_n_2458);
  not csa_tree_add_51_79_groupi_drc_bufs45890(csa_tree_add_51_79_groupi_n_1103 ,csa_tree_add_51_79_groupi_n_2455);
  not csa_tree_add_51_79_groupi_drc_bufs45894(csa_tree_add_51_79_groupi_n_1102 ,csa_tree_add_51_79_groupi_n_2467);
  not csa_tree_add_51_79_groupi_drc_bufs45898(csa_tree_add_51_79_groupi_n_1101 ,csa_tree_add_51_79_groupi_n_2476);
  not csa_tree_add_51_79_groupi_drc_bufs45902(csa_tree_add_51_79_groupi_n_1100 ,csa_tree_add_51_79_groupi_n_2473);
  not csa_tree_add_51_79_groupi_drc_bufs45906(csa_tree_add_51_79_groupi_n_1099 ,csa_tree_add_51_79_groupi_n_2470);
  not csa_tree_add_51_79_groupi_drc_bufs45910(csa_tree_add_51_79_groupi_n_1098 ,csa_tree_add_51_79_groupi_n_1968);
  not csa_tree_add_51_79_groupi_drc_bufs45914(csa_tree_add_51_79_groupi_n_1097 ,csa_tree_add_51_79_groupi_n_2461);
  not csa_tree_add_51_79_groupi_drc_bufs45918(csa_tree_add_51_79_groupi_n_1096 ,csa_tree_add_51_79_groupi_n_2464);
  not csa_tree_add_51_79_groupi_drc_bufs45922(csa_tree_add_51_79_groupi_n_1095 ,csa_tree_add_51_79_groupi_n_2439);
  not csa_tree_add_51_79_groupi_drc_bufs45926(csa_tree_add_51_79_groupi_n_1094 ,csa_tree_add_51_79_groupi_n_2436);
  not csa_tree_add_51_79_groupi_drc_bufs45930(csa_tree_add_51_79_groupi_n_1093 ,csa_tree_add_51_79_groupi_n_2003);
  not csa_tree_add_51_79_groupi_drc_bufs45934(csa_tree_add_51_79_groupi_n_1092 ,csa_tree_add_51_79_groupi_n_1993);
  not csa_tree_add_51_79_groupi_drc_bufs45938(csa_tree_add_51_79_groupi_n_1091 ,csa_tree_add_51_79_groupi_n_1974);
  not csa_tree_add_51_79_groupi_drc_bufs45942(csa_tree_add_51_79_groupi_n_1090 ,csa_tree_add_51_79_groupi_n_2495);
  not csa_tree_add_51_79_groupi_drc_bufs45946(csa_tree_add_51_79_groupi_n_1089 ,csa_tree_add_51_79_groupi_n_2492);
  not csa_tree_add_51_79_groupi_drc_bufs45950(csa_tree_add_51_79_groupi_n_1088 ,csa_tree_add_51_79_groupi_n_2503);
  not csa_tree_add_51_79_groupi_drc_bufs45954(csa_tree_add_51_79_groupi_n_1087 ,csa_tree_add_51_79_groupi_n_2009);
  not csa_tree_add_51_79_groupi_drc_bufs45958(csa_tree_add_51_79_groupi_n_1086 ,csa_tree_add_51_79_groupi_n_2489);
  not csa_tree_add_51_79_groupi_drc_bufs45962(csa_tree_add_51_79_groupi_n_1085 ,csa_tree_add_51_79_groupi_n_1084);
  not csa_tree_add_51_79_groupi_drc_bufs45964(csa_tree_add_51_79_groupi_n_1084 ,csa_tree_add_51_79_groupi_n_2538);
  not csa_tree_add_51_79_groupi_drc_bufs45966(csa_tree_add_51_79_groupi_n_1083 ,csa_tree_add_51_79_groupi_n_1082);
  not csa_tree_add_51_79_groupi_drc_bufs45968(csa_tree_add_51_79_groupi_n_1082 ,csa_tree_add_51_79_groupi_n_2524);
  not csa_tree_add_51_79_groupi_drc_bufs45970(csa_tree_add_51_79_groupi_n_1081 ,csa_tree_add_51_79_groupi_n_1080);
  not csa_tree_add_51_79_groupi_drc_bufs45972(csa_tree_add_51_79_groupi_n_1080 ,csa_tree_add_51_79_groupi_n_2515);
  not csa_tree_add_51_79_groupi_drc_bufs45974(csa_tree_add_51_79_groupi_n_1079 ,csa_tree_add_51_79_groupi_n_1078);
  not csa_tree_add_51_79_groupi_drc_bufs45976(csa_tree_add_51_79_groupi_n_1078 ,csa_tree_add_51_79_groupi_n_2518);
  not csa_tree_add_51_79_groupi_drc_bufs45997(csa_tree_add_51_79_groupi_n_1077 ,csa_tree_add_51_79_groupi_n_1722);
  not csa_tree_add_51_79_groupi_drc_bufs46001(csa_tree_add_51_79_groupi_n_1076 ,csa_tree_add_51_79_groupi_n_1720);
  not csa_tree_add_51_79_groupi_drc_bufs46005(csa_tree_add_51_79_groupi_n_1075 ,csa_tree_add_51_79_groupi_n_1774);
  not csa_tree_add_51_79_groupi_drc_bufs46009(csa_tree_add_51_79_groupi_n_1074 ,csa_tree_add_51_79_groupi_n_1775);
  not csa_tree_add_51_79_groupi_drc_bufs46013(csa_tree_add_51_79_groupi_n_1073 ,csa_tree_add_51_79_groupi_n_1721);
  not csa_tree_add_51_79_groupi_drc_bufs46017(csa_tree_add_51_79_groupi_n_1072 ,csa_tree_add_51_79_groupi_n_1777);
  not csa_tree_add_51_79_groupi_drc_bufs46021(csa_tree_add_51_79_groupi_n_1071 ,csa_tree_add_51_79_groupi_n_1776);
  not csa_tree_add_51_79_groupi_drc_bufs46027(csa_tree_add_51_79_groupi_n_1530 ,csa_tree_add_51_79_groupi_n_7599);
  not csa_tree_add_51_79_groupi_drc_bufs46030(csa_tree_add_51_79_groupi_n_1070 ,csa_tree_add_51_79_groupi_n_1529);
  not csa_tree_add_51_79_groupi_drc_bufs46031(csa_tree_add_51_79_groupi_n_1529 ,csa_tree_add_51_79_groupi_n_7310);
  not csa_tree_add_51_79_groupi_drc_bufs46034(csa_tree_add_51_79_groupi_n_1069 ,csa_tree_add_51_79_groupi_n_1528);
  not csa_tree_add_51_79_groupi_drc_bufs46035(csa_tree_add_51_79_groupi_n_1528 ,csa_tree_add_51_79_groupi_n_5854);
  not csa_tree_add_51_79_groupi_drc_bufs46277(csa_tree_add_51_79_groupi_n_1068 ,csa_tree_add_51_79_groupi_n_1066);
  not csa_tree_add_51_79_groupi_drc_bufs46279(csa_tree_add_51_79_groupi_n_1066 ,csa_tree_add_51_79_groupi_n_3731);
  not csa_tree_add_51_79_groupi_drc_bufs46281(csa_tree_add_51_79_groupi_n_1065 ,csa_tree_add_51_79_groupi_n_1063);
  not csa_tree_add_51_79_groupi_drc_bufs46283(csa_tree_add_51_79_groupi_n_1063 ,csa_tree_add_51_79_groupi_n_3186);
  not csa_tree_add_51_79_groupi_drc_bufs46285(csa_tree_add_51_79_groupi_n_1062 ,csa_tree_add_51_79_groupi_n_1060);
  not csa_tree_add_51_79_groupi_drc_bufs46287(csa_tree_add_51_79_groupi_n_1060 ,csa_tree_add_51_79_groupi_n_3172);
  not csa_tree_add_51_79_groupi_drc_bufs46289(csa_tree_add_51_79_groupi_n_1059 ,csa_tree_add_51_79_groupi_n_1057);
  not csa_tree_add_51_79_groupi_drc_bufs46291(csa_tree_add_51_79_groupi_n_1057 ,csa_tree_add_51_79_groupi_n_3184);
  not csa_tree_add_51_79_groupi_drc_bufs46293(csa_tree_add_51_79_groupi_n_1056 ,csa_tree_add_51_79_groupi_n_1054);
  not csa_tree_add_51_79_groupi_drc_bufs46295(csa_tree_add_51_79_groupi_n_1054 ,csa_tree_add_51_79_groupi_n_3179);
  not csa_tree_add_51_79_groupi_drc_bufs46297(csa_tree_add_51_79_groupi_n_1053 ,csa_tree_add_51_79_groupi_n_1051);
  not csa_tree_add_51_79_groupi_drc_bufs46299(csa_tree_add_51_79_groupi_n_1051 ,csa_tree_add_51_79_groupi_n_3170);
  not csa_tree_add_51_79_groupi_drc_bufs46301(csa_tree_add_51_79_groupi_n_1050 ,csa_tree_add_51_79_groupi_n_1048);
  not csa_tree_add_51_79_groupi_drc_bufs46303(csa_tree_add_51_79_groupi_n_1048 ,csa_tree_add_51_79_groupi_n_3181);
  not csa_tree_add_51_79_groupi_drc_bufs46305(csa_tree_add_51_79_groupi_n_1047 ,csa_tree_add_51_79_groupi_n_1045);
  not csa_tree_add_51_79_groupi_drc_bufs46307(csa_tree_add_51_79_groupi_n_1045 ,csa_tree_add_51_79_groupi_n_3165);
  not csa_tree_add_51_79_groupi_drc_bufs46309(csa_tree_add_51_79_groupi_n_1044 ,csa_tree_add_51_79_groupi_n_1042);
  not csa_tree_add_51_79_groupi_drc_bufs46311(csa_tree_add_51_79_groupi_n_1042 ,csa_tree_add_51_79_groupi_n_3178);
  not csa_tree_add_51_79_groupi_drc_bufs46313(csa_tree_add_51_79_groupi_n_1041 ,csa_tree_add_51_79_groupi_n_1039);
  not csa_tree_add_51_79_groupi_drc_bufs46315(csa_tree_add_51_79_groupi_n_1039 ,csa_tree_add_51_79_groupi_n_3727);
  not csa_tree_add_51_79_groupi_drc_bufs46317(csa_tree_add_51_79_groupi_n_1038 ,csa_tree_add_51_79_groupi_n_1036);
  not csa_tree_add_51_79_groupi_drc_bufs46319(csa_tree_add_51_79_groupi_n_1036 ,csa_tree_add_51_79_groupi_n_3722);
  not csa_tree_add_51_79_groupi_drc_bufs46321(csa_tree_add_51_79_groupi_n_1035 ,csa_tree_add_51_79_groupi_n_1033);
  not csa_tree_add_51_79_groupi_drc_bufs46323(csa_tree_add_51_79_groupi_n_1033 ,csa_tree_add_51_79_groupi_n_3709);
  not csa_tree_add_51_79_groupi_drc_bufs46325(csa_tree_add_51_79_groupi_n_1032 ,csa_tree_add_51_79_groupi_n_1030);
  not csa_tree_add_51_79_groupi_drc_bufs46327(csa_tree_add_51_79_groupi_n_1030 ,csa_tree_add_51_79_groupi_n_3176);
  not csa_tree_add_51_79_groupi_drc_bufs46329(csa_tree_add_51_79_groupi_n_1029 ,csa_tree_add_51_79_groupi_n_1027);
  not csa_tree_add_51_79_groupi_drc_bufs46331(csa_tree_add_51_79_groupi_n_1027 ,csa_tree_add_51_79_groupi_n_3705);
  not csa_tree_add_51_79_groupi_drc_bufs46333(csa_tree_add_51_79_groupi_n_1026 ,csa_tree_add_51_79_groupi_n_1024);
  not csa_tree_add_51_79_groupi_drc_bufs46335(csa_tree_add_51_79_groupi_n_1024 ,csa_tree_add_51_79_groupi_n_3180);
  not csa_tree_add_51_79_groupi_drc_bufs46337(csa_tree_add_51_79_groupi_n_1023 ,csa_tree_add_51_79_groupi_n_1021);
  not csa_tree_add_51_79_groupi_drc_bufs46339(csa_tree_add_51_79_groupi_n_1021 ,csa_tree_add_51_79_groupi_n_3188);
  not csa_tree_add_51_79_groupi_drc_bufs46341(csa_tree_add_51_79_groupi_n_1020 ,csa_tree_add_51_79_groupi_n_1018);
  not csa_tree_add_51_79_groupi_drc_bufs46343(csa_tree_add_51_79_groupi_n_1018 ,csa_tree_add_51_79_groupi_n_3173);
  not csa_tree_add_51_79_groupi_drc_bufs46345(csa_tree_add_51_79_groupi_n_1017 ,csa_tree_add_51_79_groupi_n_1015);
  not csa_tree_add_51_79_groupi_drc_bufs46347(csa_tree_add_51_79_groupi_n_1015 ,csa_tree_add_51_79_groupi_n_3187);
  not csa_tree_add_51_79_groupi_drc_bufs46349(csa_tree_add_51_79_groupi_n_1014 ,csa_tree_add_51_79_groupi_n_1012);
  not csa_tree_add_51_79_groupi_drc_bufs46351(csa_tree_add_51_79_groupi_n_1012 ,csa_tree_add_51_79_groupi_n_3714);
  not csa_tree_add_51_79_groupi_drc_bufs46353(csa_tree_add_51_79_groupi_n_1011 ,csa_tree_add_51_79_groupi_n_1009);
  not csa_tree_add_51_79_groupi_drc_bufs46355(csa_tree_add_51_79_groupi_n_1009 ,csa_tree_add_51_79_groupi_n_3163);
  not csa_tree_add_51_79_groupi_drc_bufs46357(csa_tree_add_51_79_groupi_n_1008 ,csa_tree_add_51_79_groupi_n_1006);
  not csa_tree_add_51_79_groupi_drc_bufs46359(csa_tree_add_51_79_groupi_n_1006 ,csa_tree_add_51_79_groupi_n_3161);
  not csa_tree_add_51_79_groupi_drc_bufs46361(csa_tree_add_51_79_groupi_n_1005 ,csa_tree_add_51_79_groupi_n_1003);
  not csa_tree_add_51_79_groupi_drc_bufs46363(csa_tree_add_51_79_groupi_n_1003 ,csa_tree_add_51_79_groupi_n_3713);
  not csa_tree_add_51_79_groupi_drc_bufs46365(csa_tree_add_51_79_groupi_n_1002 ,csa_tree_add_51_79_groupi_n_1000);
  not csa_tree_add_51_79_groupi_drc_bufs46367(csa_tree_add_51_79_groupi_n_1000 ,csa_tree_add_51_79_groupi_n_3712);
  not csa_tree_add_51_79_groupi_drc_bufs46369(csa_tree_add_51_79_groupi_n_999 ,csa_tree_add_51_79_groupi_n_997);
  not csa_tree_add_51_79_groupi_drc_bufs46371(csa_tree_add_51_79_groupi_n_997 ,csa_tree_add_51_79_groupi_n_3159);
  not csa_tree_add_51_79_groupi_drc_bufs46373(csa_tree_add_51_79_groupi_n_996 ,csa_tree_add_51_79_groupi_n_994);
  not csa_tree_add_51_79_groupi_drc_bufs46375(csa_tree_add_51_79_groupi_n_994 ,csa_tree_add_51_79_groupi_n_3711);
  not csa_tree_add_51_79_groupi_drc_bufs46377(csa_tree_add_51_79_groupi_n_993 ,csa_tree_add_51_79_groupi_n_991);
  not csa_tree_add_51_79_groupi_drc_bufs46379(csa_tree_add_51_79_groupi_n_991 ,csa_tree_add_51_79_groupi_n_3723);
  not csa_tree_add_51_79_groupi_drc_bufs46381(csa_tree_add_51_79_groupi_n_990 ,csa_tree_add_51_79_groupi_n_988);
  not csa_tree_add_51_79_groupi_drc_bufs46383(csa_tree_add_51_79_groupi_n_988 ,csa_tree_add_51_79_groupi_n_3710);
  not csa_tree_add_51_79_groupi_drc_bufs46385(csa_tree_add_51_79_groupi_n_987 ,csa_tree_add_51_79_groupi_n_985);
  not csa_tree_add_51_79_groupi_drc_bufs46387(csa_tree_add_51_79_groupi_n_985 ,csa_tree_add_51_79_groupi_n_3730);
  not csa_tree_add_51_79_groupi_drc_bufs46389(csa_tree_add_51_79_groupi_n_984 ,csa_tree_add_51_79_groupi_n_982);
  not csa_tree_add_51_79_groupi_drc_bufs46391(csa_tree_add_51_79_groupi_n_982 ,csa_tree_add_51_79_groupi_n_3183);
  not csa_tree_add_51_79_groupi_drc_bufs46393(csa_tree_add_51_79_groupi_n_981 ,csa_tree_add_51_79_groupi_n_979);
  not csa_tree_add_51_79_groupi_drc_bufs46395(csa_tree_add_51_79_groupi_n_979 ,csa_tree_add_51_79_groupi_n_3707);
  not csa_tree_add_51_79_groupi_drc_bufs46397(csa_tree_add_51_79_groupi_n_978 ,csa_tree_add_51_79_groupi_n_976);
  not csa_tree_add_51_79_groupi_drc_bufs46399(csa_tree_add_51_79_groupi_n_976 ,csa_tree_add_51_79_groupi_n_3706);
  not csa_tree_add_51_79_groupi_drc_bufs46401(csa_tree_add_51_79_groupi_n_975 ,csa_tree_add_51_79_groupi_n_973);
  not csa_tree_add_51_79_groupi_drc_bufs46403(csa_tree_add_51_79_groupi_n_973 ,csa_tree_add_51_79_groupi_n_3182);
  not csa_tree_add_51_79_groupi_drc_bufs46405(csa_tree_add_51_79_groupi_n_972 ,csa_tree_add_51_79_groupi_n_970);
  not csa_tree_add_51_79_groupi_drc_bufs46407(csa_tree_add_51_79_groupi_n_970 ,csa_tree_add_51_79_groupi_n_3732);
  not csa_tree_add_51_79_groupi_drc_bufs46409(csa_tree_add_51_79_groupi_n_969 ,csa_tree_add_51_79_groupi_n_967);
  not csa_tree_add_51_79_groupi_drc_bufs46411(csa_tree_add_51_79_groupi_n_967 ,csa_tree_add_51_79_groupi_n_3190);
  not csa_tree_add_51_79_groupi_drc_bufs46413(csa_tree_add_51_79_groupi_n_966 ,csa_tree_add_51_79_groupi_n_964);
  not csa_tree_add_51_79_groupi_drc_bufs46415(csa_tree_add_51_79_groupi_n_964 ,csa_tree_add_51_79_groupi_n_3177);
  not csa_tree_add_51_79_groupi_drc_bufs46417(csa_tree_add_51_79_groupi_n_963 ,csa_tree_add_51_79_groupi_n_961);
  not csa_tree_add_51_79_groupi_drc_bufs46419(csa_tree_add_51_79_groupi_n_961 ,csa_tree_add_51_79_groupi_n_3728);
  not csa_tree_add_51_79_groupi_drc_bufs46421(csa_tree_add_51_79_groupi_n_960 ,csa_tree_add_51_79_groupi_n_958);
  not csa_tree_add_51_79_groupi_drc_bufs46423(csa_tree_add_51_79_groupi_n_958 ,csa_tree_add_51_79_groupi_n_3189);
  not csa_tree_add_51_79_groupi_drc_bufs46425(csa_tree_add_51_79_groupi_n_957 ,csa_tree_add_51_79_groupi_n_955);
  not csa_tree_add_51_79_groupi_drc_bufs46427(csa_tree_add_51_79_groupi_n_955 ,csa_tree_add_51_79_groupi_n_3174);
  not csa_tree_add_51_79_groupi_drc_bufs46429(csa_tree_add_51_79_groupi_n_954 ,csa_tree_add_51_79_groupi_n_952);
  not csa_tree_add_51_79_groupi_drc_bufs46431(csa_tree_add_51_79_groupi_n_952 ,csa_tree_add_51_79_groupi_n_3729);
  not csa_tree_add_51_79_groupi_drc_bufs46433(csa_tree_add_51_79_groupi_n_951 ,csa_tree_add_51_79_groupi_n_949);
  not csa_tree_add_51_79_groupi_drc_bufs46435(csa_tree_add_51_79_groupi_n_949 ,csa_tree_add_51_79_groupi_n_3185);
  not csa_tree_add_51_79_groupi_drc_bufs46437(csa_tree_add_51_79_groupi_n_948 ,csa_tree_add_51_79_groupi_n_946);
  not csa_tree_add_51_79_groupi_drc_bufs46439(csa_tree_add_51_79_groupi_n_946 ,csa_tree_add_51_79_groupi_n_3721);
  not csa_tree_add_51_79_groupi_drc_bufs46441(csa_tree_add_51_79_groupi_n_945 ,csa_tree_add_51_79_groupi_n_943);
  not csa_tree_add_51_79_groupi_drc_bufs46443(csa_tree_add_51_79_groupi_n_943 ,csa_tree_add_51_79_groupi_n_3725);
  not csa_tree_add_51_79_groupi_drc_bufs46445(csa_tree_add_51_79_groupi_n_942 ,csa_tree_add_51_79_groupi_n_940);
  not csa_tree_add_51_79_groupi_drc_bufs46447(csa_tree_add_51_79_groupi_n_940 ,csa_tree_add_51_79_groupi_n_3724);
  not csa_tree_add_51_79_groupi_drc_bufs46449(csa_tree_add_51_79_groupi_n_939 ,csa_tree_add_51_79_groupi_n_937);
  not csa_tree_add_51_79_groupi_drc_bufs46451(csa_tree_add_51_79_groupi_n_937 ,csa_tree_add_51_79_groupi_n_3175);
  not csa_tree_add_51_79_groupi_drc_bufs46453(csa_tree_add_51_79_groupi_n_936 ,csa_tree_add_51_79_groupi_n_934);
  not csa_tree_add_51_79_groupi_drc_bufs46455(csa_tree_add_51_79_groupi_n_934 ,csa_tree_add_51_79_groupi_n_3720);
  not csa_tree_add_51_79_groupi_drc_bufs46457(csa_tree_add_51_79_groupi_n_933 ,csa_tree_add_51_79_groupi_n_931);
  not csa_tree_add_51_79_groupi_drc_bufs46459(csa_tree_add_51_79_groupi_n_931 ,csa_tree_add_51_79_groupi_n_3169);
  not csa_tree_add_51_79_groupi_drc_bufs46461(csa_tree_add_51_79_groupi_n_930 ,csa_tree_add_51_79_groupi_n_928);
  not csa_tree_add_51_79_groupi_drc_bufs46463(csa_tree_add_51_79_groupi_n_928 ,csa_tree_add_51_79_groupi_n_3719);
  not csa_tree_add_51_79_groupi_drc_bufs46465(csa_tree_add_51_79_groupi_n_927 ,csa_tree_add_51_79_groupi_n_925);
  not csa_tree_add_51_79_groupi_drc_bufs46467(csa_tree_add_51_79_groupi_n_925 ,csa_tree_add_51_79_groupi_n_3168);
  not csa_tree_add_51_79_groupi_drc_bufs46469(csa_tree_add_51_79_groupi_n_924 ,csa_tree_add_51_79_groupi_n_922);
  not csa_tree_add_51_79_groupi_drc_bufs46471(csa_tree_add_51_79_groupi_n_922 ,csa_tree_add_51_79_groupi_n_3167);
  not csa_tree_add_51_79_groupi_drc_bufs46473(csa_tree_add_51_79_groupi_n_921 ,csa_tree_add_51_79_groupi_n_919);
  not csa_tree_add_51_79_groupi_drc_bufs46475(csa_tree_add_51_79_groupi_n_919 ,csa_tree_add_51_79_groupi_n_3171);
  not csa_tree_add_51_79_groupi_drc_bufs46477(csa_tree_add_51_79_groupi_n_918 ,csa_tree_add_51_79_groupi_n_916);
  not csa_tree_add_51_79_groupi_drc_bufs46479(csa_tree_add_51_79_groupi_n_916 ,csa_tree_add_51_79_groupi_n_3164);
  not csa_tree_add_51_79_groupi_drc_bufs46481(csa_tree_add_51_79_groupi_n_915 ,csa_tree_add_51_79_groupi_n_913);
  not csa_tree_add_51_79_groupi_drc_bufs46483(csa_tree_add_51_79_groupi_n_913 ,csa_tree_add_51_79_groupi_n_3162);
  not csa_tree_add_51_79_groupi_drc_bufs46485(csa_tree_add_51_79_groupi_n_912 ,csa_tree_add_51_79_groupi_n_910);
  not csa_tree_add_51_79_groupi_drc_bufs46487(csa_tree_add_51_79_groupi_n_910 ,csa_tree_add_51_79_groupi_n_3718);
  not csa_tree_add_51_79_groupi_drc_bufs46489(csa_tree_add_51_79_groupi_n_909 ,csa_tree_add_51_79_groupi_n_907);
  not csa_tree_add_51_79_groupi_drc_bufs46491(csa_tree_add_51_79_groupi_n_907 ,csa_tree_add_51_79_groupi_n_3716);
  not csa_tree_add_51_79_groupi_drc_bufs46493(csa_tree_add_51_79_groupi_n_906 ,csa_tree_add_51_79_groupi_n_904);
  not csa_tree_add_51_79_groupi_drc_bufs46495(csa_tree_add_51_79_groupi_n_904 ,csa_tree_add_51_79_groupi_n_3160);
  not csa_tree_add_51_79_groupi_drc_bufs46497(csa_tree_add_51_79_groupi_n_903 ,csa_tree_add_51_79_groupi_n_901);
  not csa_tree_add_51_79_groupi_drc_bufs46499(csa_tree_add_51_79_groupi_n_901 ,csa_tree_add_51_79_groupi_n_3717);
  not csa_tree_add_51_79_groupi_drc_bufs46501(csa_tree_add_51_79_groupi_n_900 ,csa_tree_add_51_79_groupi_n_898);
  not csa_tree_add_51_79_groupi_drc_bufs46503(csa_tree_add_51_79_groupi_n_898 ,csa_tree_add_51_79_groupi_n_3708);
  not csa_tree_add_51_79_groupi_drc_bufs46505(csa_tree_add_51_79_groupi_n_897 ,csa_tree_add_51_79_groupi_n_895);
  not csa_tree_add_51_79_groupi_drc_bufs46507(csa_tree_add_51_79_groupi_n_895 ,csa_tree_add_51_79_groupi_n_3715);
  not csa_tree_add_51_79_groupi_drc_bufs46509(csa_tree_add_51_79_groupi_n_894 ,csa_tree_add_51_79_groupi_n_892);
  not csa_tree_add_51_79_groupi_drc_bufs46511(csa_tree_add_51_79_groupi_n_892 ,csa_tree_add_51_79_groupi_n_3726);
  not csa_tree_add_51_79_groupi_drc_bufs46513(csa_tree_add_51_79_groupi_n_891 ,csa_tree_add_51_79_groupi_n_889);
  not csa_tree_add_51_79_groupi_drc_bufs46515(csa_tree_add_51_79_groupi_n_889 ,csa_tree_add_51_79_groupi_n_3166);
  not csa_tree_add_51_79_groupi_drc_bufs46518(csa_tree_add_51_79_groupi_n_888 ,csa_tree_add_51_79_groupi_n_887);
  not csa_tree_add_51_79_groupi_drc_bufs46519(csa_tree_add_51_79_groupi_n_887 ,csa_tree_add_51_79_groupi_n_1643);
  not csa_tree_add_51_79_groupi_drc_bufs46522(csa_tree_add_51_79_groupi_n_886 ,csa_tree_add_51_79_groupi_n_885);
  not csa_tree_add_51_79_groupi_drc_bufs46523(csa_tree_add_51_79_groupi_n_885 ,csa_tree_add_51_79_groupi_n_1642);
  not csa_tree_add_51_79_groupi_drc_bufs46530(csa_tree_add_51_79_groupi_n_881 ,csa_tree_add_51_79_groupi_n_880);
  not csa_tree_add_51_79_groupi_drc_bufs46531(csa_tree_add_51_79_groupi_n_880 ,csa_tree_add_51_79_groupi_n_1576);
  not csa_tree_add_51_79_groupi_drc_bufs46538(csa_tree_add_51_79_groupi_n_876 ,csa_tree_add_51_79_groupi_n_875);
  not csa_tree_add_51_79_groupi_drc_bufs46539(csa_tree_add_51_79_groupi_n_875 ,csa_tree_add_51_79_groupi_n_1575);
  not csa_tree_add_51_79_groupi_drc_bufs46546(csa_tree_add_51_79_groupi_n_871 ,csa_tree_add_51_79_groupi_n_870);
  not csa_tree_add_51_79_groupi_drc_bufs46547(csa_tree_add_51_79_groupi_n_870 ,csa_tree_add_51_79_groupi_n_1573);
  not csa_tree_add_51_79_groupi_drc_bufs46550(csa_tree_add_51_79_groupi_n_869 ,csa_tree_add_51_79_groupi_n_868);
  not csa_tree_add_51_79_groupi_drc_bufs46551(csa_tree_add_51_79_groupi_n_868 ,csa_tree_add_51_79_groupi_n_1571);
  not csa_tree_add_51_79_groupi_drc_bufs46558(csa_tree_add_51_79_groupi_n_864 ,csa_tree_add_51_79_groupi_n_863);
  not csa_tree_add_51_79_groupi_drc_bufs46559(csa_tree_add_51_79_groupi_n_863 ,csa_tree_add_51_79_groupi_n_1569);
  not csa_tree_add_51_79_groupi_drc_bufs46562(csa_tree_add_51_79_groupi_n_862 ,csa_tree_add_51_79_groupi_n_861);
  not csa_tree_add_51_79_groupi_drc_bufs46563(csa_tree_add_51_79_groupi_n_861 ,csa_tree_add_51_79_groupi_n_1641);
  not csa_tree_add_51_79_groupi_drc_bufs46570(csa_tree_add_51_79_groupi_n_857 ,csa_tree_add_51_79_groupi_n_856);
  not csa_tree_add_51_79_groupi_drc_bufs46571(csa_tree_add_51_79_groupi_n_856 ,csa_tree_add_51_79_groupi_n_1570);
  not csa_tree_add_51_79_groupi_drc_bufs46578(csa_tree_add_51_79_groupi_n_852 ,csa_tree_add_51_79_groupi_n_851);
  not csa_tree_add_51_79_groupi_drc_bufs46579(csa_tree_add_51_79_groupi_n_851 ,csa_tree_add_51_79_groupi_n_1631);
  not csa_tree_add_51_79_groupi_drc_bufs46582(csa_tree_add_51_79_groupi_n_850 ,csa_tree_add_51_79_groupi_n_849);
  not csa_tree_add_51_79_groupi_drc_bufs46583(csa_tree_add_51_79_groupi_n_849 ,csa_tree_add_51_79_groupi_n_1630);
  not csa_tree_add_51_79_groupi_drc_bufs46586(csa_tree_add_51_79_groupi_n_848 ,csa_tree_add_51_79_groupi_n_847);
  not csa_tree_add_51_79_groupi_drc_bufs46587(csa_tree_add_51_79_groupi_n_847 ,csa_tree_add_51_79_groupi_n_1629);
  not csa_tree_add_51_79_groupi_drc_bufs46590(csa_tree_add_51_79_groupi_n_846 ,csa_tree_add_51_79_groupi_n_845);
  not csa_tree_add_51_79_groupi_drc_bufs46591(csa_tree_add_51_79_groupi_n_845 ,csa_tree_add_51_79_groupi_n_1628);
  not csa_tree_add_51_79_groupi_drc_bufs46594(csa_tree_add_51_79_groupi_n_844 ,csa_tree_add_51_79_groupi_n_843);
  not csa_tree_add_51_79_groupi_drc_bufs46595(csa_tree_add_51_79_groupi_n_843 ,csa_tree_add_51_79_groupi_n_1564);
  not csa_tree_add_51_79_groupi_drc_bufs46598(csa_tree_add_51_79_groupi_n_842 ,csa_tree_add_51_79_groupi_n_841);
  not csa_tree_add_51_79_groupi_drc_bufs46599(csa_tree_add_51_79_groupi_n_841 ,csa_tree_add_51_79_groupi_n_1563);
  not csa_tree_add_51_79_groupi_drc_bufs46602(csa_tree_add_51_79_groupi_n_840 ,csa_tree_add_51_79_groupi_n_839);
  not csa_tree_add_51_79_groupi_drc_bufs46603(csa_tree_add_51_79_groupi_n_839 ,csa_tree_add_51_79_groupi_n_1560);
  not csa_tree_add_51_79_groupi_drc_bufs46606(csa_tree_add_51_79_groupi_n_838 ,csa_tree_add_51_79_groupi_n_837);
  not csa_tree_add_51_79_groupi_drc_bufs46607(csa_tree_add_51_79_groupi_n_837 ,csa_tree_add_51_79_groupi_n_1558);
  not csa_tree_add_51_79_groupi_drc_bufs46610(csa_tree_add_51_79_groupi_n_836 ,csa_tree_add_51_79_groupi_n_835);
  not csa_tree_add_51_79_groupi_drc_bufs46611(csa_tree_add_51_79_groupi_n_835 ,csa_tree_add_51_79_groupi_n_1562);
  not csa_tree_add_51_79_groupi_drc_bufs46622(csa_tree_add_51_79_groupi_n_828 ,csa_tree_add_51_79_groupi_n_827);
  not csa_tree_add_51_79_groupi_drc_bufs46623(csa_tree_add_51_79_groupi_n_827 ,csa_tree_add_51_79_groupi_n_1644);
  not csa_tree_add_51_79_groupi_drc_bufs46630(csa_tree_add_51_79_groupi_n_823 ,csa_tree_add_51_79_groupi_n_822);
  not csa_tree_add_51_79_groupi_drc_bufs46631(csa_tree_add_51_79_groupi_n_822 ,csa_tree_add_51_79_groupi_n_1574);
  not csa_tree_add_51_79_groupi_drc_bufs46634(csa_tree_add_51_79_groupi_n_821 ,csa_tree_add_51_79_groupi_n_820);
  not csa_tree_add_51_79_groupi_drc_bufs46635(csa_tree_add_51_79_groupi_n_820 ,csa_tree_add_51_79_groupi_n_1572);
  not csa_tree_add_51_79_groupi_drc_bufs46649(csa_tree_add_51_79_groupi_n_810 ,csa_tree_add_51_79_groupi_n_808);
  not csa_tree_add_51_79_groupi_drc_bufs46651(csa_tree_add_51_79_groupi_n_808 ,csa_tree_add_51_79_groupi_n_1559);
  not csa_tree_add_51_79_groupi_drc_bufs46653(csa_tree_add_51_79_groupi_n_807 ,csa_tree_add_51_79_groupi_n_805);
  not csa_tree_add_51_79_groupi_drc_bufs46655(csa_tree_add_51_79_groupi_n_805 ,csa_tree_add_51_79_groupi_n_1561);
  not csa_tree_add_51_79_groupi_drc_bufs46665(csa_tree_add_51_79_groupi_n_798 ,csa_tree_add_51_79_groupi_n_796);
  not csa_tree_add_51_79_groupi_drc_bufs46667(csa_tree_add_51_79_groupi_n_796 ,csa_tree_add_51_79_groupi_n_1632);
  not csa_tree_add_51_79_groupi_drc_bufs46709(csa_tree_add_51_79_groupi_n_765 ,csa_tree_add_51_79_groupi_n_764);
  not csa_tree_add_51_79_groupi_drc_bufs46711(csa_tree_add_51_79_groupi_n_764 ,csa_tree_add_51_79_groupi_n_4793);
  not csa_tree_add_51_79_groupi_drc_bufs46714(csa_tree_add_51_79_groupi_n_763 ,csa_tree_add_51_79_groupi_n_4811);
  not csa_tree_add_51_79_groupi_drc_bufs46727(csa_tree_add_51_79_groupi_n_1521 ,csa_tree_add_51_79_groupi_n_2521);
  not csa_tree_add_51_79_groupi_drc_bufs46731(csa_tree_add_51_79_groupi_n_1527 ,csa_tree_add_51_79_groupi_n_2531);
  not csa_tree_add_51_79_groupi_drc_bufs46743(csa_tree_add_51_79_groupi_n_1524 ,csa_tree_add_51_79_groupi_n_2527);
  not csa_tree_add_51_79_groupi_drc_bufs46753(csa_tree_add_51_79_groupi_n_751 ,csa_tree_add_51_79_groupi_n_749);
  not csa_tree_add_51_79_groupi_drc_bufs46755(csa_tree_add_51_79_groupi_n_749 ,csa_tree_add_51_79_groupi_n_1213);
  not csa_tree_add_51_79_groupi_drc_bufs46757(csa_tree_add_51_79_groupi_n_748 ,csa_tree_add_51_79_groupi_n_746);
  not csa_tree_add_51_79_groupi_drc_bufs46759(csa_tree_add_51_79_groupi_n_746 ,csa_tree_add_51_79_groupi_n_1264);
  not csa_tree_add_51_79_groupi_drc_bufs46761(csa_tree_add_51_79_groupi_n_745 ,csa_tree_add_51_79_groupi_n_743);
  not csa_tree_add_51_79_groupi_drc_bufs46763(csa_tree_add_51_79_groupi_n_743 ,csa_tree_add_51_79_groupi_n_1255);
  not csa_tree_add_51_79_groupi_drc_bufs46765(csa_tree_add_51_79_groupi_n_742 ,csa_tree_add_51_79_groupi_n_740);
  not csa_tree_add_51_79_groupi_drc_bufs46767(csa_tree_add_51_79_groupi_n_740 ,csa_tree_add_51_79_groupi_n_1081);
  not csa_tree_add_51_79_groupi_drc_bufs46769(csa_tree_add_51_79_groupi_n_739 ,csa_tree_add_51_79_groupi_n_737);
  not csa_tree_add_51_79_groupi_drc_bufs46771(csa_tree_add_51_79_groupi_n_737 ,csa_tree_add_51_79_groupi_n_1228);
  not csa_tree_add_51_79_groupi_drc_bufs46773(csa_tree_add_51_79_groupi_n_736 ,csa_tree_add_51_79_groupi_n_734);
  not csa_tree_add_51_79_groupi_drc_bufs46775(csa_tree_add_51_79_groupi_n_734 ,csa_tree_add_51_79_groupi_n_1216);
  not csa_tree_add_51_79_groupi_drc_bufs46781(csa_tree_add_51_79_groupi_n_730 ,csa_tree_add_51_79_groupi_n_728);
  not csa_tree_add_51_79_groupi_drc_bufs46783(csa_tree_add_51_79_groupi_n_728 ,csa_tree_add_51_79_groupi_n_1252);
  not csa_tree_add_51_79_groupi_drc_bufs46785(csa_tree_add_51_79_groupi_n_727 ,csa_tree_add_51_79_groupi_n_725);
  not csa_tree_add_51_79_groupi_drc_bufs46787(csa_tree_add_51_79_groupi_n_725 ,csa_tree_add_51_79_groupi_n_1085);
  not csa_tree_add_51_79_groupi_drc_bufs46789(csa_tree_add_51_79_groupi_n_724 ,csa_tree_add_51_79_groupi_n_722);
  not csa_tree_add_51_79_groupi_drc_bufs46791(csa_tree_add_51_79_groupi_n_722 ,csa_tree_add_51_79_groupi_n_1222);
  not csa_tree_add_51_79_groupi_drc_bufs46797(csa_tree_add_51_79_groupi_n_718 ,csa_tree_add_51_79_groupi_n_716);
  not csa_tree_add_51_79_groupi_drc_bufs46799(csa_tree_add_51_79_groupi_n_716 ,csa_tree_add_51_79_groupi_n_1079);
  not csa_tree_add_51_79_groupi_drc_bufs46805(csa_tree_add_51_79_groupi_n_712 ,csa_tree_add_51_79_groupi_n_710);
  not csa_tree_add_51_79_groupi_drc_bufs46807(csa_tree_add_51_79_groupi_n_710 ,csa_tree_add_51_79_groupi_n_1225);
  not csa_tree_add_51_79_groupi_drc_bufs46809(csa_tree_add_51_79_groupi_n_709 ,csa_tree_add_51_79_groupi_n_707);
  not csa_tree_add_51_79_groupi_drc_bufs46811(csa_tree_add_51_79_groupi_n_707 ,csa_tree_add_51_79_groupi_n_1234);
  not csa_tree_add_51_79_groupi_drc_bufs46813(csa_tree_add_51_79_groupi_n_706 ,csa_tree_add_51_79_groupi_n_704);
  not csa_tree_add_51_79_groupi_drc_bufs46815(csa_tree_add_51_79_groupi_n_704 ,csa_tree_add_51_79_groupi_n_1240);
  not csa_tree_add_51_79_groupi_drc_bufs46821(csa_tree_add_51_79_groupi_n_700 ,csa_tree_add_51_79_groupi_n_698);
  not csa_tree_add_51_79_groupi_drc_bufs46823(csa_tree_add_51_79_groupi_n_698 ,csa_tree_add_51_79_groupi_n_1261);
  not csa_tree_add_51_79_groupi_drc_bufs46825(csa_tree_add_51_79_groupi_n_697 ,csa_tree_add_51_79_groupi_n_695);
  not csa_tree_add_51_79_groupi_drc_bufs46827(csa_tree_add_51_79_groupi_n_695 ,csa_tree_add_51_79_groupi_n_1258);
  not csa_tree_add_51_79_groupi_drc_bufs46829(csa_tree_add_51_79_groupi_n_694 ,csa_tree_add_51_79_groupi_n_692);
  not csa_tree_add_51_79_groupi_drc_bufs46831(csa_tree_add_51_79_groupi_n_692 ,csa_tree_add_51_79_groupi_n_1249);
  not csa_tree_add_51_79_groupi_drc_bufs46841(csa_tree_add_51_79_groupi_n_685 ,csa_tree_add_51_79_groupi_n_683);
  not csa_tree_add_51_79_groupi_drc_bufs46843(csa_tree_add_51_79_groupi_n_683 ,csa_tree_add_51_79_groupi_n_1246);
  not csa_tree_add_51_79_groupi_drc_bufs46845(csa_tree_add_51_79_groupi_n_682 ,csa_tree_add_51_79_groupi_n_680);
  not csa_tree_add_51_79_groupi_drc_bufs46847(csa_tree_add_51_79_groupi_n_680 ,csa_tree_add_51_79_groupi_n_1237);
  not csa_tree_add_51_79_groupi_drc_bufs46853(csa_tree_add_51_79_groupi_n_676 ,csa_tree_add_51_79_groupi_n_674);
  not csa_tree_add_51_79_groupi_drc_bufs46855(csa_tree_add_51_79_groupi_n_674 ,csa_tree_add_51_79_groupi_n_1243);
  not csa_tree_add_51_79_groupi_drc_bufs46857(csa_tree_add_51_79_groupi_n_673 ,csa_tree_add_51_79_groupi_n_671);
  not csa_tree_add_51_79_groupi_drc_bufs46859(csa_tree_add_51_79_groupi_n_671 ,csa_tree_add_51_79_groupi_n_1219);
  not csa_tree_add_51_79_groupi_drc_bufs46861(csa_tree_add_51_79_groupi_n_670 ,csa_tree_add_51_79_groupi_n_668);
  not csa_tree_add_51_79_groupi_drc_bufs46863(csa_tree_add_51_79_groupi_n_668 ,csa_tree_add_51_79_groupi_n_1083);
  not csa_tree_add_51_79_groupi_drc_bufs46877(csa_tree_add_51_79_groupi_n_658 ,csa_tree_add_51_79_groupi_n_656);
  not csa_tree_add_51_79_groupi_drc_bufs46879(csa_tree_add_51_79_groupi_n_656 ,csa_tree_add_51_79_groupi_n_1231);
  not csa_tree_add_51_79_groupi_drc_bufs46945(csa_tree_add_51_79_groupi_n_607 ,csa_tree_add_51_79_groupi_n_606);
  not csa_tree_add_51_79_groupi_drc_bufs46947(csa_tree_add_51_79_groupi_n_606 ,csa_tree_add_51_79_groupi_n_828);
  not csa_tree_add_51_79_groupi_drc_bufs46949(csa_tree_add_51_79_groupi_n_605 ,csa_tree_add_51_79_groupi_n_604);
  not csa_tree_add_51_79_groupi_drc_bufs46951(csa_tree_add_51_79_groupi_n_604 ,csa_tree_add_51_79_groupi_n_823);
  not csa_tree_add_51_79_groupi_drc_bufs46953(csa_tree_add_51_79_groupi_n_603 ,csa_tree_add_51_79_groupi_n_602);
  not csa_tree_add_51_79_groupi_drc_bufs46955(csa_tree_add_51_79_groupi_n_602 ,csa_tree_add_51_79_groupi_n_821);
  not csa_tree_add_51_79_groupi_drc_bufs46957(csa_tree_add_51_79_groupi_n_601 ,csa_tree_add_51_79_groupi_n_599);
  not csa_tree_add_51_79_groupi_drc_bufs46958(csa_tree_add_51_79_groupi_n_600 ,csa_tree_add_51_79_groupi_n_599);
  not csa_tree_add_51_79_groupi_drc_bufs46959(csa_tree_add_51_79_groupi_n_599 ,csa_tree_add_51_79_groupi_n_1572);
  not csa_tree_add_51_79_groupi_drc_bufs46961(csa_tree_add_51_79_groupi_n_598 ,csa_tree_add_51_79_groupi_n_596);
  not csa_tree_add_51_79_groupi_drc_bufs46962(csa_tree_add_51_79_groupi_n_597 ,csa_tree_add_51_79_groupi_n_596);
  not csa_tree_add_51_79_groupi_drc_bufs46963(csa_tree_add_51_79_groupi_n_596 ,csa_tree_add_51_79_groupi_n_1574);
  not csa_tree_add_51_79_groupi_drc_bufs46965(csa_tree_add_51_79_groupi_n_595 ,csa_tree_add_51_79_groupi_n_594);
  not csa_tree_add_51_79_groupi_drc_bufs46967(csa_tree_add_51_79_groupi_n_594 ,csa_tree_add_51_79_groupi_n_888);
  not csa_tree_add_51_79_groupi_drc_bufs46969(csa_tree_add_51_79_groupi_n_593 ,csa_tree_add_51_79_groupi_n_591);
  not csa_tree_add_51_79_groupi_drc_bufs46970(csa_tree_add_51_79_groupi_n_592 ,csa_tree_add_51_79_groupi_n_591);
  not csa_tree_add_51_79_groupi_drc_bufs46971(csa_tree_add_51_79_groupi_n_591 ,csa_tree_add_51_79_groupi_n_1644);
  not csa_tree_add_51_79_groupi_drc_bufs46973(csa_tree_add_51_79_groupi_n_590 ,csa_tree_add_51_79_groupi_n_589);
  not csa_tree_add_51_79_groupi_drc_bufs46975(csa_tree_add_51_79_groupi_n_589 ,csa_tree_add_51_79_groupi_n_871);
  not csa_tree_add_51_79_groupi_drc_bufs46977(csa_tree_add_51_79_groupi_n_588 ,csa_tree_add_51_79_groupi_n_587);
  not csa_tree_add_51_79_groupi_drc_bufs46979(csa_tree_add_51_79_groupi_n_587 ,csa_tree_add_51_79_groupi_n_864);
  not csa_tree_add_51_79_groupi_drc_bufs46981(csa_tree_add_51_79_groupi_n_586 ,csa_tree_add_51_79_groupi_n_584);
  not csa_tree_add_51_79_groupi_drc_bufs46982(csa_tree_add_51_79_groupi_n_585 ,csa_tree_add_51_79_groupi_n_584);
  not csa_tree_add_51_79_groupi_drc_bufs46983(csa_tree_add_51_79_groupi_n_584 ,csa_tree_add_51_79_groupi_n_1562);
  not csa_tree_add_51_79_groupi_drc_bufs46985(csa_tree_add_51_79_groupi_n_583 ,csa_tree_add_51_79_groupi_n_581);
  not csa_tree_add_51_79_groupi_drc_bufs46986(csa_tree_add_51_79_groupi_n_582 ,csa_tree_add_51_79_groupi_n_581);
  not csa_tree_add_51_79_groupi_drc_bufs46987(csa_tree_add_51_79_groupi_n_581 ,csa_tree_add_51_79_groupi_n_1558);
  not csa_tree_add_51_79_groupi_drc_bufs46989(csa_tree_add_51_79_groupi_n_580 ,csa_tree_add_51_79_groupi_n_578);
  not csa_tree_add_51_79_groupi_drc_bufs46990(csa_tree_add_51_79_groupi_n_579 ,csa_tree_add_51_79_groupi_n_578);
  not csa_tree_add_51_79_groupi_drc_bufs46991(csa_tree_add_51_79_groupi_n_578 ,csa_tree_add_51_79_groupi_n_1560);
  not csa_tree_add_51_79_groupi_drc_bufs46993(csa_tree_add_51_79_groupi_n_577 ,csa_tree_add_51_79_groupi_n_575);
  not csa_tree_add_51_79_groupi_drc_bufs46994(csa_tree_add_51_79_groupi_n_576 ,csa_tree_add_51_79_groupi_n_575);
  not csa_tree_add_51_79_groupi_drc_bufs46995(csa_tree_add_51_79_groupi_n_575 ,csa_tree_add_51_79_groupi_n_1563);
  not csa_tree_add_51_79_groupi_drc_bufs46997(csa_tree_add_51_79_groupi_n_574 ,csa_tree_add_51_79_groupi_n_572);
  not csa_tree_add_51_79_groupi_drc_bufs46998(csa_tree_add_51_79_groupi_n_573 ,csa_tree_add_51_79_groupi_n_572);
  not csa_tree_add_51_79_groupi_drc_bufs46999(csa_tree_add_51_79_groupi_n_572 ,csa_tree_add_51_79_groupi_n_1564);
  not csa_tree_add_51_79_groupi_drc_bufs47001(csa_tree_add_51_79_groupi_n_571 ,csa_tree_add_51_79_groupi_n_569);
  not csa_tree_add_51_79_groupi_drc_bufs47002(csa_tree_add_51_79_groupi_n_570 ,csa_tree_add_51_79_groupi_n_569);
  not csa_tree_add_51_79_groupi_drc_bufs47003(csa_tree_add_51_79_groupi_n_569 ,csa_tree_add_51_79_groupi_n_1628);
  not csa_tree_add_51_79_groupi_drc_bufs47005(csa_tree_add_51_79_groupi_n_568 ,csa_tree_add_51_79_groupi_n_566);
  not csa_tree_add_51_79_groupi_drc_bufs47006(csa_tree_add_51_79_groupi_n_567 ,csa_tree_add_51_79_groupi_n_566);
  not csa_tree_add_51_79_groupi_drc_bufs47007(csa_tree_add_51_79_groupi_n_566 ,csa_tree_add_51_79_groupi_n_1629);
  not csa_tree_add_51_79_groupi_drc_bufs47009(csa_tree_add_51_79_groupi_n_565 ,csa_tree_add_51_79_groupi_n_563);
  not csa_tree_add_51_79_groupi_drc_bufs47010(csa_tree_add_51_79_groupi_n_564 ,csa_tree_add_51_79_groupi_n_563);
  not csa_tree_add_51_79_groupi_drc_bufs47011(csa_tree_add_51_79_groupi_n_563 ,csa_tree_add_51_79_groupi_n_1630);
  not csa_tree_add_51_79_groupi_drc_bufs47013(csa_tree_add_51_79_groupi_n_562 ,csa_tree_add_51_79_groupi_n_560);
  not csa_tree_add_51_79_groupi_drc_bufs47014(csa_tree_add_51_79_groupi_n_561 ,csa_tree_add_51_79_groupi_n_560);
  not csa_tree_add_51_79_groupi_drc_bufs47015(csa_tree_add_51_79_groupi_n_560 ,csa_tree_add_51_79_groupi_n_1631);
  not csa_tree_add_51_79_groupi_drc_bufs47017(csa_tree_add_51_79_groupi_n_559 ,csa_tree_add_51_79_groupi_n_558);
  not csa_tree_add_51_79_groupi_drc_bufs47019(csa_tree_add_51_79_groupi_n_558 ,csa_tree_add_51_79_groupi_n_857);
  not csa_tree_add_51_79_groupi_drc_bufs47021(csa_tree_add_51_79_groupi_n_557 ,csa_tree_add_51_79_groupi_n_555);
  not csa_tree_add_51_79_groupi_drc_bufs47022(csa_tree_add_51_79_groupi_n_556 ,csa_tree_add_51_79_groupi_n_555);
  not csa_tree_add_51_79_groupi_drc_bufs47023(csa_tree_add_51_79_groupi_n_555 ,csa_tree_add_51_79_groupi_n_1570);
  not csa_tree_add_51_79_groupi_drc_bufs47025(csa_tree_add_51_79_groupi_n_554 ,csa_tree_add_51_79_groupi_n_553);
  not csa_tree_add_51_79_groupi_drc_bufs47027(csa_tree_add_51_79_groupi_n_553 ,csa_tree_add_51_79_groupi_n_862);
  not csa_tree_add_51_79_groupi_drc_bufs47029(csa_tree_add_51_79_groupi_n_552 ,csa_tree_add_51_79_groupi_n_550);
  not csa_tree_add_51_79_groupi_drc_bufs47030(csa_tree_add_51_79_groupi_n_551 ,csa_tree_add_51_79_groupi_n_550);
  not csa_tree_add_51_79_groupi_drc_bufs47031(csa_tree_add_51_79_groupi_n_550 ,csa_tree_add_51_79_groupi_n_1641);
  not csa_tree_add_51_79_groupi_drc_bufs47033(csa_tree_add_51_79_groupi_n_549 ,csa_tree_add_51_79_groupi_n_547);
  not csa_tree_add_51_79_groupi_drc_bufs47034(csa_tree_add_51_79_groupi_n_548 ,csa_tree_add_51_79_groupi_n_547);
  not csa_tree_add_51_79_groupi_drc_bufs47035(csa_tree_add_51_79_groupi_n_547 ,csa_tree_add_51_79_groupi_n_1569);
  not csa_tree_add_51_79_groupi_drc_bufs47037(csa_tree_add_51_79_groupi_n_546 ,csa_tree_add_51_79_groupi_n_545);
  not csa_tree_add_51_79_groupi_drc_bufs47039(csa_tree_add_51_79_groupi_n_545 ,csa_tree_add_51_79_groupi_n_869);
  not csa_tree_add_51_79_groupi_drc_bufs47041(csa_tree_add_51_79_groupi_n_544 ,csa_tree_add_51_79_groupi_n_542);
  not csa_tree_add_51_79_groupi_drc_bufs47042(csa_tree_add_51_79_groupi_n_543 ,csa_tree_add_51_79_groupi_n_542);
  not csa_tree_add_51_79_groupi_drc_bufs47043(csa_tree_add_51_79_groupi_n_542 ,csa_tree_add_51_79_groupi_n_1571);
  not csa_tree_add_51_79_groupi_drc_bufs47045(csa_tree_add_51_79_groupi_n_541 ,csa_tree_add_51_79_groupi_n_539);
  not csa_tree_add_51_79_groupi_drc_bufs47046(csa_tree_add_51_79_groupi_n_540 ,csa_tree_add_51_79_groupi_n_539);
  not csa_tree_add_51_79_groupi_drc_bufs47047(csa_tree_add_51_79_groupi_n_539 ,csa_tree_add_51_79_groupi_n_1573);
  not csa_tree_add_51_79_groupi_drc_bufs47049(csa_tree_add_51_79_groupi_n_538 ,csa_tree_add_51_79_groupi_n_537);
  not csa_tree_add_51_79_groupi_drc_bufs47051(csa_tree_add_51_79_groupi_n_537 ,csa_tree_add_51_79_groupi_n_876);
  not csa_tree_add_51_79_groupi_drc_bufs47053(csa_tree_add_51_79_groupi_n_536 ,csa_tree_add_51_79_groupi_n_534);
  not csa_tree_add_51_79_groupi_drc_bufs47054(csa_tree_add_51_79_groupi_n_535 ,csa_tree_add_51_79_groupi_n_534);
  not csa_tree_add_51_79_groupi_drc_bufs47055(csa_tree_add_51_79_groupi_n_534 ,csa_tree_add_51_79_groupi_n_1575);
  not csa_tree_add_51_79_groupi_drc_bufs47057(csa_tree_add_51_79_groupi_n_533 ,csa_tree_add_51_79_groupi_n_532);
  not csa_tree_add_51_79_groupi_drc_bufs47059(csa_tree_add_51_79_groupi_n_532 ,csa_tree_add_51_79_groupi_n_881);
  not csa_tree_add_51_79_groupi_drc_bufs47061(csa_tree_add_51_79_groupi_n_531 ,csa_tree_add_51_79_groupi_n_529);
  not csa_tree_add_51_79_groupi_drc_bufs47062(csa_tree_add_51_79_groupi_n_530 ,csa_tree_add_51_79_groupi_n_529);
  not csa_tree_add_51_79_groupi_drc_bufs47063(csa_tree_add_51_79_groupi_n_529 ,csa_tree_add_51_79_groupi_n_1576);
  not csa_tree_add_51_79_groupi_drc_bufs47065(csa_tree_add_51_79_groupi_n_528 ,csa_tree_add_51_79_groupi_n_527);
  not csa_tree_add_51_79_groupi_drc_bufs47067(csa_tree_add_51_79_groupi_n_527 ,csa_tree_add_51_79_groupi_n_886);
  not csa_tree_add_51_79_groupi_drc_bufs47069(csa_tree_add_51_79_groupi_n_526 ,csa_tree_add_51_79_groupi_n_524);
  not csa_tree_add_51_79_groupi_drc_bufs47070(csa_tree_add_51_79_groupi_n_525 ,csa_tree_add_51_79_groupi_n_524);
  not csa_tree_add_51_79_groupi_drc_bufs47071(csa_tree_add_51_79_groupi_n_524 ,csa_tree_add_51_79_groupi_n_1642);
  not csa_tree_add_51_79_groupi_drc_bufs47073(csa_tree_add_51_79_groupi_n_523 ,csa_tree_add_51_79_groupi_n_521);
  not csa_tree_add_51_79_groupi_drc_bufs47074(csa_tree_add_51_79_groupi_n_522 ,csa_tree_add_51_79_groupi_n_521);
  not csa_tree_add_51_79_groupi_drc_bufs47075(csa_tree_add_51_79_groupi_n_521 ,csa_tree_add_51_79_groupi_n_1643);
  not csa_tree_add_51_79_groupi_drc_bufs47077(csa_tree_add_51_79_groupi_n_520 ,csa_tree_add_51_79_groupi_n_519);
  not csa_tree_add_51_79_groupi_drc_bufs47079(csa_tree_add_51_79_groupi_n_519 ,csa_tree_add_51_79_groupi_n_891);
  not csa_tree_add_51_79_groupi_drc_bufs47081(csa_tree_add_51_79_groupi_n_518 ,csa_tree_add_51_79_groupi_n_517);
  not csa_tree_add_51_79_groupi_drc_bufs47083(csa_tree_add_51_79_groupi_n_517 ,csa_tree_add_51_79_groupi_n_894);
  not csa_tree_add_51_79_groupi_drc_bufs47085(csa_tree_add_51_79_groupi_n_516 ,csa_tree_add_51_79_groupi_n_515);
  not csa_tree_add_51_79_groupi_drc_bufs47087(csa_tree_add_51_79_groupi_n_515 ,csa_tree_add_51_79_groupi_n_897);
  not csa_tree_add_51_79_groupi_drc_bufs47089(csa_tree_add_51_79_groupi_n_514 ,csa_tree_add_51_79_groupi_n_513);
  not csa_tree_add_51_79_groupi_drc_bufs47091(csa_tree_add_51_79_groupi_n_513 ,csa_tree_add_51_79_groupi_n_900);
  not csa_tree_add_51_79_groupi_drc_bufs47093(csa_tree_add_51_79_groupi_n_512 ,csa_tree_add_51_79_groupi_n_511);
  not csa_tree_add_51_79_groupi_drc_bufs47095(csa_tree_add_51_79_groupi_n_511 ,csa_tree_add_51_79_groupi_n_903);
  not csa_tree_add_51_79_groupi_drc_bufs47097(csa_tree_add_51_79_groupi_n_510 ,csa_tree_add_51_79_groupi_n_509);
  not csa_tree_add_51_79_groupi_drc_bufs47099(csa_tree_add_51_79_groupi_n_509 ,csa_tree_add_51_79_groupi_n_906);
  not csa_tree_add_51_79_groupi_drc_bufs47101(csa_tree_add_51_79_groupi_n_508 ,csa_tree_add_51_79_groupi_n_507);
  not csa_tree_add_51_79_groupi_drc_bufs47103(csa_tree_add_51_79_groupi_n_507 ,csa_tree_add_51_79_groupi_n_909);
  not csa_tree_add_51_79_groupi_drc_bufs47105(csa_tree_add_51_79_groupi_n_506 ,csa_tree_add_51_79_groupi_n_505);
  not csa_tree_add_51_79_groupi_drc_bufs47107(csa_tree_add_51_79_groupi_n_505 ,csa_tree_add_51_79_groupi_n_912);
  not csa_tree_add_51_79_groupi_drc_bufs47109(csa_tree_add_51_79_groupi_n_504 ,csa_tree_add_51_79_groupi_n_503);
  not csa_tree_add_51_79_groupi_drc_bufs47111(csa_tree_add_51_79_groupi_n_503 ,csa_tree_add_51_79_groupi_n_915);
  not csa_tree_add_51_79_groupi_drc_bufs47113(csa_tree_add_51_79_groupi_n_502 ,csa_tree_add_51_79_groupi_n_501);
  not csa_tree_add_51_79_groupi_drc_bufs47115(csa_tree_add_51_79_groupi_n_501 ,csa_tree_add_51_79_groupi_n_918);
  not csa_tree_add_51_79_groupi_drc_bufs47117(csa_tree_add_51_79_groupi_n_500 ,csa_tree_add_51_79_groupi_n_499);
  not csa_tree_add_51_79_groupi_drc_bufs47119(csa_tree_add_51_79_groupi_n_499 ,csa_tree_add_51_79_groupi_n_921);
  not csa_tree_add_51_79_groupi_drc_bufs47121(csa_tree_add_51_79_groupi_n_498 ,csa_tree_add_51_79_groupi_n_497);
  not csa_tree_add_51_79_groupi_drc_bufs47123(csa_tree_add_51_79_groupi_n_497 ,csa_tree_add_51_79_groupi_n_924);
  not csa_tree_add_51_79_groupi_drc_bufs47125(csa_tree_add_51_79_groupi_n_496 ,csa_tree_add_51_79_groupi_n_495);
  not csa_tree_add_51_79_groupi_drc_bufs47127(csa_tree_add_51_79_groupi_n_495 ,csa_tree_add_51_79_groupi_n_927);
  not csa_tree_add_51_79_groupi_drc_bufs47129(csa_tree_add_51_79_groupi_n_494 ,csa_tree_add_51_79_groupi_n_493);
  not csa_tree_add_51_79_groupi_drc_bufs47131(csa_tree_add_51_79_groupi_n_493 ,csa_tree_add_51_79_groupi_n_930);
  not csa_tree_add_51_79_groupi_drc_bufs47133(csa_tree_add_51_79_groupi_n_492 ,csa_tree_add_51_79_groupi_n_491);
  not csa_tree_add_51_79_groupi_drc_bufs47135(csa_tree_add_51_79_groupi_n_491 ,csa_tree_add_51_79_groupi_n_933);
  not csa_tree_add_51_79_groupi_drc_bufs47137(csa_tree_add_51_79_groupi_n_490 ,csa_tree_add_51_79_groupi_n_489);
  not csa_tree_add_51_79_groupi_drc_bufs47139(csa_tree_add_51_79_groupi_n_489 ,csa_tree_add_51_79_groupi_n_936);
  not csa_tree_add_51_79_groupi_drc_bufs47141(csa_tree_add_51_79_groupi_n_488 ,csa_tree_add_51_79_groupi_n_487);
  not csa_tree_add_51_79_groupi_drc_bufs47143(csa_tree_add_51_79_groupi_n_487 ,csa_tree_add_51_79_groupi_n_939);
  not csa_tree_add_51_79_groupi_drc_bufs47145(csa_tree_add_51_79_groupi_n_486 ,csa_tree_add_51_79_groupi_n_485);
  not csa_tree_add_51_79_groupi_drc_bufs47147(csa_tree_add_51_79_groupi_n_485 ,csa_tree_add_51_79_groupi_n_942);
  not csa_tree_add_51_79_groupi_drc_bufs47149(csa_tree_add_51_79_groupi_n_484 ,csa_tree_add_51_79_groupi_n_483);
  not csa_tree_add_51_79_groupi_drc_bufs47151(csa_tree_add_51_79_groupi_n_483 ,csa_tree_add_51_79_groupi_n_945);
  not csa_tree_add_51_79_groupi_drc_bufs47153(csa_tree_add_51_79_groupi_n_482 ,csa_tree_add_51_79_groupi_n_481);
  not csa_tree_add_51_79_groupi_drc_bufs47155(csa_tree_add_51_79_groupi_n_481 ,csa_tree_add_51_79_groupi_n_948);
  not csa_tree_add_51_79_groupi_drc_bufs47157(csa_tree_add_51_79_groupi_n_480 ,csa_tree_add_51_79_groupi_n_479);
  not csa_tree_add_51_79_groupi_drc_bufs47159(csa_tree_add_51_79_groupi_n_479 ,csa_tree_add_51_79_groupi_n_951);
  not csa_tree_add_51_79_groupi_drc_bufs47161(csa_tree_add_51_79_groupi_n_478 ,csa_tree_add_51_79_groupi_n_477);
  not csa_tree_add_51_79_groupi_drc_bufs47163(csa_tree_add_51_79_groupi_n_477 ,csa_tree_add_51_79_groupi_n_954);
  not csa_tree_add_51_79_groupi_drc_bufs47165(csa_tree_add_51_79_groupi_n_476 ,csa_tree_add_51_79_groupi_n_475);
  not csa_tree_add_51_79_groupi_drc_bufs47167(csa_tree_add_51_79_groupi_n_475 ,csa_tree_add_51_79_groupi_n_957);
  not csa_tree_add_51_79_groupi_drc_bufs47169(csa_tree_add_51_79_groupi_n_474 ,csa_tree_add_51_79_groupi_n_473);
  not csa_tree_add_51_79_groupi_drc_bufs47171(csa_tree_add_51_79_groupi_n_473 ,csa_tree_add_51_79_groupi_n_960);
  not csa_tree_add_51_79_groupi_drc_bufs47173(csa_tree_add_51_79_groupi_n_472 ,csa_tree_add_51_79_groupi_n_471);
  not csa_tree_add_51_79_groupi_drc_bufs47175(csa_tree_add_51_79_groupi_n_471 ,csa_tree_add_51_79_groupi_n_963);
  not csa_tree_add_51_79_groupi_drc_bufs47177(csa_tree_add_51_79_groupi_n_470 ,csa_tree_add_51_79_groupi_n_469);
  not csa_tree_add_51_79_groupi_drc_bufs47179(csa_tree_add_51_79_groupi_n_469 ,csa_tree_add_51_79_groupi_n_966);
  not csa_tree_add_51_79_groupi_drc_bufs47181(csa_tree_add_51_79_groupi_n_468 ,csa_tree_add_51_79_groupi_n_467);
  not csa_tree_add_51_79_groupi_drc_bufs47183(csa_tree_add_51_79_groupi_n_467 ,csa_tree_add_51_79_groupi_n_969);
  not csa_tree_add_51_79_groupi_drc_bufs47185(csa_tree_add_51_79_groupi_n_466 ,csa_tree_add_51_79_groupi_n_465);
  not csa_tree_add_51_79_groupi_drc_bufs47187(csa_tree_add_51_79_groupi_n_465 ,csa_tree_add_51_79_groupi_n_972);
  not csa_tree_add_51_79_groupi_drc_bufs47189(csa_tree_add_51_79_groupi_n_464 ,csa_tree_add_51_79_groupi_n_463);
  not csa_tree_add_51_79_groupi_drc_bufs47191(csa_tree_add_51_79_groupi_n_463 ,csa_tree_add_51_79_groupi_n_975);
  not csa_tree_add_51_79_groupi_drc_bufs47193(csa_tree_add_51_79_groupi_n_462 ,csa_tree_add_51_79_groupi_n_461);
  not csa_tree_add_51_79_groupi_drc_bufs47195(csa_tree_add_51_79_groupi_n_461 ,csa_tree_add_51_79_groupi_n_978);
  not csa_tree_add_51_79_groupi_drc_bufs47197(csa_tree_add_51_79_groupi_n_460 ,csa_tree_add_51_79_groupi_n_459);
  not csa_tree_add_51_79_groupi_drc_bufs47199(csa_tree_add_51_79_groupi_n_459 ,csa_tree_add_51_79_groupi_n_981);
  not csa_tree_add_51_79_groupi_drc_bufs47201(csa_tree_add_51_79_groupi_n_458 ,csa_tree_add_51_79_groupi_n_457);
  not csa_tree_add_51_79_groupi_drc_bufs47203(csa_tree_add_51_79_groupi_n_457 ,csa_tree_add_51_79_groupi_n_984);
  not csa_tree_add_51_79_groupi_drc_bufs47205(csa_tree_add_51_79_groupi_n_456 ,csa_tree_add_51_79_groupi_n_455);
  not csa_tree_add_51_79_groupi_drc_bufs47207(csa_tree_add_51_79_groupi_n_455 ,csa_tree_add_51_79_groupi_n_987);
  not csa_tree_add_51_79_groupi_drc_bufs47209(csa_tree_add_51_79_groupi_n_454 ,csa_tree_add_51_79_groupi_n_453);
  not csa_tree_add_51_79_groupi_drc_bufs47211(csa_tree_add_51_79_groupi_n_453 ,csa_tree_add_51_79_groupi_n_990);
  not csa_tree_add_51_79_groupi_drc_bufs47213(csa_tree_add_51_79_groupi_n_452 ,csa_tree_add_51_79_groupi_n_451);
  not csa_tree_add_51_79_groupi_drc_bufs47215(csa_tree_add_51_79_groupi_n_451 ,csa_tree_add_51_79_groupi_n_993);
  not csa_tree_add_51_79_groupi_drc_bufs47217(csa_tree_add_51_79_groupi_n_450 ,csa_tree_add_51_79_groupi_n_449);
  not csa_tree_add_51_79_groupi_drc_bufs47219(csa_tree_add_51_79_groupi_n_449 ,csa_tree_add_51_79_groupi_n_996);
  not csa_tree_add_51_79_groupi_drc_bufs47221(csa_tree_add_51_79_groupi_n_448 ,csa_tree_add_51_79_groupi_n_447);
  not csa_tree_add_51_79_groupi_drc_bufs47223(csa_tree_add_51_79_groupi_n_447 ,csa_tree_add_51_79_groupi_n_999);
  not csa_tree_add_51_79_groupi_drc_bufs47225(csa_tree_add_51_79_groupi_n_446 ,csa_tree_add_51_79_groupi_n_445);
  not csa_tree_add_51_79_groupi_drc_bufs47227(csa_tree_add_51_79_groupi_n_445 ,csa_tree_add_51_79_groupi_n_1002);
  not csa_tree_add_51_79_groupi_drc_bufs47229(csa_tree_add_51_79_groupi_n_444 ,csa_tree_add_51_79_groupi_n_443);
  not csa_tree_add_51_79_groupi_drc_bufs47231(csa_tree_add_51_79_groupi_n_443 ,csa_tree_add_51_79_groupi_n_1005);
  not csa_tree_add_51_79_groupi_drc_bufs47233(csa_tree_add_51_79_groupi_n_442 ,csa_tree_add_51_79_groupi_n_441);
  not csa_tree_add_51_79_groupi_drc_bufs47235(csa_tree_add_51_79_groupi_n_441 ,csa_tree_add_51_79_groupi_n_1008);
  not csa_tree_add_51_79_groupi_drc_bufs47237(csa_tree_add_51_79_groupi_n_440 ,csa_tree_add_51_79_groupi_n_439);
  not csa_tree_add_51_79_groupi_drc_bufs47239(csa_tree_add_51_79_groupi_n_439 ,csa_tree_add_51_79_groupi_n_1011);
  not csa_tree_add_51_79_groupi_drc_bufs47241(csa_tree_add_51_79_groupi_n_438 ,csa_tree_add_51_79_groupi_n_437);
  not csa_tree_add_51_79_groupi_drc_bufs47243(csa_tree_add_51_79_groupi_n_437 ,csa_tree_add_51_79_groupi_n_1014);
  not csa_tree_add_51_79_groupi_drc_bufs47245(csa_tree_add_51_79_groupi_n_436 ,csa_tree_add_51_79_groupi_n_435);
  not csa_tree_add_51_79_groupi_drc_bufs47247(csa_tree_add_51_79_groupi_n_435 ,csa_tree_add_51_79_groupi_n_1017);
  not csa_tree_add_51_79_groupi_drc_bufs47249(csa_tree_add_51_79_groupi_n_434 ,csa_tree_add_51_79_groupi_n_433);
  not csa_tree_add_51_79_groupi_drc_bufs47251(csa_tree_add_51_79_groupi_n_433 ,csa_tree_add_51_79_groupi_n_1020);
  not csa_tree_add_51_79_groupi_drc_bufs47253(csa_tree_add_51_79_groupi_n_432 ,csa_tree_add_51_79_groupi_n_431);
  not csa_tree_add_51_79_groupi_drc_bufs47255(csa_tree_add_51_79_groupi_n_431 ,csa_tree_add_51_79_groupi_n_1023);
  not csa_tree_add_51_79_groupi_drc_bufs47257(csa_tree_add_51_79_groupi_n_430 ,csa_tree_add_51_79_groupi_n_429);
  not csa_tree_add_51_79_groupi_drc_bufs47259(csa_tree_add_51_79_groupi_n_429 ,csa_tree_add_51_79_groupi_n_1026);
  not csa_tree_add_51_79_groupi_drc_bufs47261(csa_tree_add_51_79_groupi_n_428 ,csa_tree_add_51_79_groupi_n_427);
  not csa_tree_add_51_79_groupi_drc_bufs47263(csa_tree_add_51_79_groupi_n_427 ,csa_tree_add_51_79_groupi_n_1029);
  not csa_tree_add_51_79_groupi_drc_bufs47265(csa_tree_add_51_79_groupi_n_426 ,csa_tree_add_51_79_groupi_n_425);
  not csa_tree_add_51_79_groupi_drc_bufs47267(csa_tree_add_51_79_groupi_n_425 ,csa_tree_add_51_79_groupi_n_1032);
  not csa_tree_add_51_79_groupi_drc_bufs47269(csa_tree_add_51_79_groupi_n_424 ,csa_tree_add_51_79_groupi_n_423);
  not csa_tree_add_51_79_groupi_drc_bufs47271(csa_tree_add_51_79_groupi_n_423 ,csa_tree_add_51_79_groupi_n_1035);
  not csa_tree_add_51_79_groupi_drc_bufs47273(csa_tree_add_51_79_groupi_n_422 ,csa_tree_add_51_79_groupi_n_421);
  not csa_tree_add_51_79_groupi_drc_bufs47275(csa_tree_add_51_79_groupi_n_421 ,csa_tree_add_51_79_groupi_n_1038);
  not csa_tree_add_51_79_groupi_drc_bufs47277(csa_tree_add_51_79_groupi_n_420 ,csa_tree_add_51_79_groupi_n_419);
  not csa_tree_add_51_79_groupi_drc_bufs47279(csa_tree_add_51_79_groupi_n_419 ,csa_tree_add_51_79_groupi_n_1041);
  not csa_tree_add_51_79_groupi_drc_bufs47281(csa_tree_add_51_79_groupi_n_418 ,csa_tree_add_51_79_groupi_n_417);
  not csa_tree_add_51_79_groupi_drc_bufs47283(csa_tree_add_51_79_groupi_n_417 ,csa_tree_add_51_79_groupi_n_1044);
  not csa_tree_add_51_79_groupi_drc_bufs47285(csa_tree_add_51_79_groupi_n_416 ,csa_tree_add_51_79_groupi_n_415);
  not csa_tree_add_51_79_groupi_drc_bufs47287(csa_tree_add_51_79_groupi_n_415 ,csa_tree_add_51_79_groupi_n_1047);
  not csa_tree_add_51_79_groupi_drc_bufs47289(csa_tree_add_51_79_groupi_n_414 ,csa_tree_add_51_79_groupi_n_413);
  not csa_tree_add_51_79_groupi_drc_bufs47291(csa_tree_add_51_79_groupi_n_413 ,csa_tree_add_51_79_groupi_n_1050);
  not csa_tree_add_51_79_groupi_drc_bufs47293(csa_tree_add_51_79_groupi_n_412 ,csa_tree_add_51_79_groupi_n_411);
  not csa_tree_add_51_79_groupi_drc_bufs47295(csa_tree_add_51_79_groupi_n_411 ,csa_tree_add_51_79_groupi_n_1053);
  not csa_tree_add_51_79_groupi_drc_bufs47297(csa_tree_add_51_79_groupi_n_410 ,csa_tree_add_51_79_groupi_n_409);
  not csa_tree_add_51_79_groupi_drc_bufs47299(csa_tree_add_51_79_groupi_n_409 ,csa_tree_add_51_79_groupi_n_1056);
  not csa_tree_add_51_79_groupi_drc_bufs47301(csa_tree_add_51_79_groupi_n_408 ,csa_tree_add_51_79_groupi_n_407);
  not csa_tree_add_51_79_groupi_drc_bufs47303(csa_tree_add_51_79_groupi_n_407 ,csa_tree_add_51_79_groupi_n_1059);
  not csa_tree_add_51_79_groupi_drc_bufs47305(csa_tree_add_51_79_groupi_n_406 ,csa_tree_add_51_79_groupi_n_405);
  not csa_tree_add_51_79_groupi_drc_bufs47307(csa_tree_add_51_79_groupi_n_405 ,csa_tree_add_51_79_groupi_n_1062);
  not csa_tree_add_51_79_groupi_drc_bufs47309(csa_tree_add_51_79_groupi_n_404 ,csa_tree_add_51_79_groupi_n_403);
  not csa_tree_add_51_79_groupi_drc_bufs47311(csa_tree_add_51_79_groupi_n_403 ,csa_tree_add_51_79_groupi_n_1065);
  not csa_tree_add_51_79_groupi_drc_bufs47313(csa_tree_add_51_79_groupi_n_402 ,csa_tree_add_51_79_groupi_n_401);
  not csa_tree_add_51_79_groupi_drc_bufs47315(csa_tree_add_51_79_groupi_n_401 ,csa_tree_add_51_79_groupi_n_1068);
  not csa_tree_add_51_79_groupi_drc_bufs47321(csa_tree_add_51_79_groupi_n_397 ,csa_tree_add_51_79_groupi_n_395);
  not csa_tree_add_51_79_groupi_drc_bufs47322(csa_tree_add_51_79_groupi_n_396 ,csa_tree_add_51_79_groupi_n_395);
  not csa_tree_add_51_79_groupi_drc_bufs47323(csa_tree_add_51_79_groupi_n_395 ,csa_tree_add_51_79_groupi_n_3714);
  not csa_tree_add_51_79_groupi_drc_bufs47329(csa_tree_add_51_79_groupi_n_391 ,csa_tree_add_51_79_groupi_n_389);
  not csa_tree_add_51_79_groupi_drc_bufs47330(csa_tree_add_51_79_groupi_n_390 ,csa_tree_add_51_79_groupi_n_389);
  not csa_tree_add_51_79_groupi_drc_bufs47331(csa_tree_add_51_79_groupi_n_389 ,csa_tree_add_51_79_groupi_n_3166);
  not csa_tree_add_51_79_groupi_drc_bufs47337(csa_tree_add_51_79_groupi_n_385 ,csa_tree_add_51_79_groupi_n_383);
  not csa_tree_add_51_79_groupi_drc_bufs47338(csa_tree_add_51_79_groupi_n_384 ,csa_tree_add_51_79_groupi_n_383);
  not csa_tree_add_51_79_groupi_drc_bufs47339(csa_tree_add_51_79_groupi_n_383 ,csa_tree_add_51_79_groupi_n_3188);
  not csa_tree_add_51_79_groupi_drc_bufs47345(csa_tree_add_51_79_groupi_n_379 ,csa_tree_add_51_79_groupi_n_377);
  not csa_tree_add_51_79_groupi_drc_bufs47346(csa_tree_add_51_79_groupi_n_378 ,csa_tree_add_51_79_groupi_n_377);
  not csa_tree_add_51_79_groupi_drc_bufs47347(csa_tree_add_51_79_groupi_n_377 ,csa_tree_add_51_79_groupi_n_3726);
  not csa_tree_add_51_79_groupi_drc_bufs47353(csa_tree_add_51_79_groupi_n_373 ,csa_tree_add_51_79_groupi_n_371);
  not csa_tree_add_51_79_groupi_drc_bufs47354(csa_tree_add_51_79_groupi_n_372 ,csa_tree_add_51_79_groupi_n_371);
  not csa_tree_add_51_79_groupi_drc_bufs47355(csa_tree_add_51_79_groupi_n_371 ,csa_tree_add_51_79_groupi_n_3708);
  not csa_tree_add_51_79_groupi_drc_bufs47361(csa_tree_add_51_79_groupi_n_367 ,csa_tree_add_51_79_groupi_n_365);
  not csa_tree_add_51_79_groupi_drc_bufs47362(csa_tree_add_51_79_groupi_n_366 ,csa_tree_add_51_79_groupi_n_365);
  not csa_tree_add_51_79_groupi_drc_bufs47363(csa_tree_add_51_79_groupi_n_365 ,csa_tree_add_51_79_groupi_n_3715);
  not csa_tree_add_51_79_groupi_drc_bufs47369(csa_tree_add_51_79_groupi_n_361 ,csa_tree_add_51_79_groupi_n_359);
  not csa_tree_add_51_79_groupi_drc_bufs47370(csa_tree_add_51_79_groupi_n_360 ,csa_tree_add_51_79_groupi_n_359);
  not csa_tree_add_51_79_groupi_drc_bufs47371(csa_tree_add_51_79_groupi_n_359 ,csa_tree_add_51_79_groupi_n_3160);
  not csa_tree_add_51_79_groupi_drc_bufs47377(csa_tree_add_51_79_groupi_n_355 ,csa_tree_add_51_79_groupi_n_353);
  not csa_tree_add_51_79_groupi_drc_bufs47378(csa_tree_add_51_79_groupi_n_354 ,csa_tree_add_51_79_groupi_n_353);
  not csa_tree_add_51_79_groupi_drc_bufs47379(csa_tree_add_51_79_groupi_n_353 ,csa_tree_add_51_79_groupi_n_3716);
  not csa_tree_add_51_79_groupi_drc_bufs47385(csa_tree_add_51_79_groupi_n_349 ,csa_tree_add_51_79_groupi_n_347);
  not csa_tree_add_51_79_groupi_drc_bufs47386(csa_tree_add_51_79_groupi_n_348 ,csa_tree_add_51_79_groupi_n_347);
  not csa_tree_add_51_79_groupi_drc_bufs47387(csa_tree_add_51_79_groupi_n_347 ,csa_tree_add_51_79_groupi_n_3717);
  not csa_tree_add_51_79_groupi_drc_bufs47393(csa_tree_add_51_79_groupi_n_343 ,csa_tree_add_51_79_groupi_n_341);
  not csa_tree_add_51_79_groupi_drc_bufs47394(csa_tree_add_51_79_groupi_n_342 ,csa_tree_add_51_79_groupi_n_341);
  not csa_tree_add_51_79_groupi_drc_bufs47395(csa_tree_add_51_79_groupi_n_341 ,csa_tree_add_51_79_groupi_n_3705);
  not csa_tree_add_51_79_groupi_drc_bufs47401(csa_tree_add_51_79_groupi_n_337 ,csa_tree_add_51_79_groupi_n_335);
  not csa_tree_add_51_79_groupi_drc_bufs47402(csa_tree_add_51_79_groupi_n_336 ,csa_tree_add_51_79_groupi_n_335);
  not csa_tree_add_51_79_groupi_drc_bufs47403(csa_tree_add_51_79_groupi_n_335 ,csa_tree_add_51_79_groupi_n_3176);
  not csa_tree_add_51_79_groupi_drc_bufs47409(csa_tree_add_51_79_groupi_n_331 ,csa_tree_add_51_79_groupi_n_329);
  not csa_tree_add_51_79_groupi_drc_bufs47410(csa_tree_add_51_79_groupi_n_330 ,csa_tree_add_51_79_groupi_n_329);
  not csa_tree_add_51_79_groupi_drc_bufs47411(csa_tree_add_51_79_groupi_n_329 ,csa_tree_add_51_79_groupi_n_3162);
  not csa_tree_add_51_79_groupi_drc_bufs47417(csa_tree_add_51_79_groupi_n_325 ,csa_tree_add_51_79_groupi_n_323);
  not csa_tree_add_51_79_groupi_drc_bufs47418(csa_tree_add_51_79_groupi_n_324 ,csa_tree_add_51_79_groupi_n_323);
  not csa_tree_add_51_79_groupi_drc_bufs47419(csa_tree_add_51_79_groupi_n_323 ,csa_tree_add_51_79_groupi_n_3164);
  not csa_tree_add_51_79_groupi_drc_bufs47425(csa_tree_add_51_79_groupi_n_319 ,csa_tree_add_51_79_groupi_n_317);
  not csa_tree_add_51_79_groupi_drc_bufs47426(csa_tree_add_51_79_groupi_n_318 ,csa_tree_add_51_79_groupi_n_317);
  not csa_tree_add_51_79_groupi_drc_bufs47427(csa_tree_add_51_79_groupi_n_317 ,csa_tree_add_51_79_groupi_n_3718);
  not csa_tree_add_51_79_groupi_drc_bufs47433(csa_tree_add_51_79_groupi_n_313 ,csa_tree_add_51_79_groupi_n_311);
  not csa_tree_add_51_79_groupi_drc_bufs47434(csa_tree_add_51_79_groupi_n_312 ,csa_tree_add_51_79_groupi_n_311);
  not csa_tree_add_51_79_groupi_drc_bufs47435(csa_tree_add_51_79_groupi_n_311 ,csa_tree_add_51_79_groupi_n_3167);
  not csa_tree_add_51_79_groupi_drc_bufs47441(csa_tree_add_51_79_groupi_n_307 ,csa_tree_add_51_79_groupi_n_305);
  not csa_tree_add_51_79_groupi_drc_bufs47442(csa_tree_add_51_79_groupi_n_306 ,csa_tree_add_51_79_groupi_n_305);
  not csa_tree_add_51_79_groupi_drc_bufs47443(csa_tree_add_51_79_groupi_n_305 ,csa_tree_add_51_79_groupi_n_3168);
  not csa_tree_add_51_79_groupi_drc_bufs47449(csa_tree_add_51_79_groupi_n_301 ,csa_tree_add_51_79_groupi_n_299);
  not csa_tree_add_51_79_groupi_drc_bufs47450(csa_tree_add_51_79_groupi_n_300 ,csa_tree_add_51_79_groupi_n_299);
  not csa_tree_add_51_79_groupi_drc_bufs47451(csa_tree_add_51_79_groupi_n_299 ,csa_tree_add_51_79_groupi_n_3171);
  not csa_tree_add_51_79_groupi_drc_bufs47457(csa_tree_add_51_79_groupi_n_295 ,csa_tree_add_51_79_groupi_n_293);
  not csa_tree_add_51_79_groupi_drc_bufs47458(csa_tree_add_51_79_groupi_n_294 ,csa_tree_add_51_79_groupi_n_293);
  not csa_tree_add_51_79_groupi_drc_bufs47459(csa_tree_add_51_79_groupi_n_293 ,csa_tree_add_51_79_groupi_n_3709);
  not csa_tree_add_51_79_groupi_drc_bufs47465(csa_tree_add_51_79_groupi_n_289 ,csa_tree_add_51_79_groupi_n_287);
  not csa_tree_add_51_79_groupi_drc_bufs47466(csa_tree_add_51_79_groupi_n_288 ,csa_tree_add_51_79_groupi_n_287);
  not csa_tree_add_51_79_groupi_drc_bufs47467(csa_tree_add_51_79_groupi_n_287 ,csa_tree_add_51_79_groupi_n_3169);
  not csa_tree_add_51_79_groupi_drc_bufs47473(csa_tree_add_51_79_groupi_n_283 ,csa_tree_add_51_79_groupi_n_281);
  not csa_tree_add_51_79_groupi_drc_bufs47474(csa_tree_add_51_79_groupi_n_282 ,csa_tree_add_51_79_groupi_n_281);
  not csa_tree_add_51_79_groupi_drc_bufs47475(csa_tree_add_51_79_groupi_n_281 ,csa_tree_add_51_79_groupi_n_3720);
  not csa_tree_add_51_79_groupi_drc_bufs47481(csa_tree_add_51_79_groupi_n_277 ,csa_tree_add_51_79_groupi_n_275);
  not csa_tree_add_51_79_groupi_drc_bufs47482(csa_tree_add_51_79_groupi_n_276 ,csa_tree_add_51_79_groupi_n_275);
  not csa_tree_add_51_79_groupi_drc_bufs47483(csa_tree_add_51_79_groupi_n_275 ,csa_tree_add_51_79_groupi_n_3719);
  not csa_tree_add_51_79_groupi_drc_bufs47489(csa_tree_add_51_79_groupi_n_271 ,csa_tree_add_51_79_groupi_n_269);
  not csa_tree_add_51_79_groupi_drc_bufs47490(csa_tree_add_51_79_groupi_n_270 ,csa_tree_add_51_79_groupi_n_269);
  not csa_tree_add_51_79_groupi_drc_bufs47491(csa_tree_add_51_79_groupi_n_269 ,csa_tree_add_51_79_groupi_n_3724);
  not csa_tree_add_51_79_groupi_drc_bufs47497(csa_tree_add_51_79_groupi_n_265 ,csa_tree_add_51_79_groupi_n_263);
  not csa_tree_add_51_79_groupi_drc_bufs47498(csa_tree_add_51_79_groupi_n_264 ,csa_tree_add_51_79_groupi_n_263);
  not csa_tree_add_51_79_groupi_drc_bufs47499(csa_tree_add_51_79_groupi_n_263 ,csa_tree_add_51_79_groupi_n_3725);
  not csa_tree_add_51_79_groupi_drc_bufs47505(csa_tree_add_51_79_groupi_n_259 ,csa_tree_add_51_79_groupi_n_257);
  not csa_tree_add_51_79_groupi_drc_bufs47506(csa_tree_add_51_79_groupi_n_258 ,csa_tree_add_51_79_groupi_n_257);
  not csa_tree_add_51_79_groupi_drc_bufs47507(csa_tree_add_51_79_groupi_n_257 ,csa_tree_add_51_79_groupi_n_3175);
  not csa_tree_add_51_79_groupi_drc_bufs47513(csa_tree_add_51_79_groupi_n_253 ,csa_tree_add_51_79_groupi_n_251);
  not csa_tree_add_51_79_groupi_drc_bufs47514(csa_tree_add_51_79_groupi_n_252 ,csa_tree_add_51_79_groupi_n_251);
  not csa_tree_add_51_79_groupi_drc_bufs47515(csa_tree_add_51_79_groupi_n_251 ,csa_tree_add_51_79_groupi_n_3727);
  not csa_tree_add_51_79_groupi_drc_bufs47521(csa_tree_add_51_79_groupi_n_247 ,csa_tree_add_51_79_groupi_n_245);
  not csa_tree_add_51_79_groupi_drc_bufs47522(csa_tree_add_51_79_groupi_n_246 ,csa_tree_add_51_79_groupi_n_245);
  not csa_tree_add_51_79_groupi_drc_bufs47523(csa_tree_add_51_79_groupi_n_245 ,csa_tree_add_51_79_groupi_n_3178);
  not csa_tree_add_51_79_groupi_drc_bufs47529(csa_tree_add_51_79_groupi_n_241 ,csa_tree_add_51_79_groupi_n_239);
  not csa_tree_add_51_79_groupi_drc_bufs47530(csa_tree_add_51_79_groupi_n_240 ,csa_tree_add_51_79_groupi_n_239);
  not csa_tree_add_51_79_groupi_drc_bufs47531(csa_tree_add_51_79_groupi_n_239 ,csa_tree_add_51_79_groupi_n_3181);
  not csa_tree_add_51_79_groupi_drc_bufs47537(csa_tree_add_51_79_groupi_n_235 ,csa_tree_add_51_79_groupi_n_233);
  not csa_tree_add_51_79_groupi_drc_bufs47538(csa_tree_add_51_79_groupi_n_234 ,csa_tree_add_51_79_groupi_n_233);
  not csa_tree_add_51_79_groupi_drc_bufs47539(csa_tree_add_51_79_groupi_n_233 ,csa_tree_add_51_79_groupi_n_3185);
  not csa_tree_add_51_79_groupi_drc_bufs47545(csa_tree_add_51_79_groupi_n_229 ,csa_tree_add_51_79_groupi_n_227);
  not csa_tree_add_51_79_groupi_drc_bufs47546(csa_tree_add_51_79_groupi_n_228 ,csa_tree_add_51_79_groupi_n_227);
  not csa_tree_add_51_79_groupi_drc_bufs47547(csa_tree_add_51_79_groupi_n_227 ,csa_tree_add_51_79_groupi_n_3729);
  not csa_tree_add_51_79_groupi_drc_bufs47553(csa_tree_add_51_79_groupi_n_223 ,csa_tree_add_51_79_groupi_n_221);
  not csa_tree_add_51_79_groupi_drc_bufs47554(csa_tree_add_51_79_groupi_n_222 ,csa_tree_add_51_79_groupi_n_221);
  not csa_tree_add_51_79_groupi_drc_bufs47555(csa_tree_add_51_79_groupi_n_221 ,csa_tree_add_51_79_groupi_n_3721);
  not csa_tree_add_51_79_groupi_drc_bufs47561(csa_tree_add_51_79_groupi_n_217 ,csa_tree_add_51_79_groupi_n_215);
  not csa_tree_add_51_79_groupi_drc_bufs47562(csa_tree_add_51_79_groupi_n_216 ,csa_tree_add_51_79_groupi_n_215);
  not csa_tree_add_51_79_groupi_drc_bufs47563(csa_tree_add_51_79_groupi_n_215 ,csa_tree_add_51_79_groupi_n_3189);
  not csa_tree_add_51_79_groupi_drc_bufs47569(csa_tree_add_51_79_groupi_n_211 ,csa_tree_add_51_79_groupi_n_209);
  not csa_tree_add_51_79_groupi_drc_bufs47570(csa_tree_add_51_79_groupi_n_210 ,csa_tree_add_51_79_groupi_n_209);
  not csa_tree_add_51_79_groupi_drc_bufs47571(csa_tree_add_51_79_groupi_n_209 ,csa_tree_add_51_79_groupi_n_3728);
  not csa_tree_add_51_79_groupi_drc_bufs47577(csa_tree_add_51_79_groupi_n_205 ,csa_tree_add_51_79_groupi_n_203);
  not csa_tree_add_51_79_groupi_drc_bufs47578(csa_tree_add_51_79_groupi_n_204 ,csa_tree_add_51_79_groupi_n_203);
  not csa_tree_add_51_79_groupi_drc_bufs47579(csa_tree_add_51_79_groupi_n_203 ,csa_tree_add_51_79_groupi_n_3174);
  not csa_tree_add_51_79_groupi_drc_bufs47585(csa_tree_add_51_79_groupi_n_199 ,csa_tree_add_51_79_groupi_n_197);
  not csa_tree_add_51_79_groupi_drc_bufs47586(csa_tree_add_51_79_groupi_n_198 ,csa_tree_add_51_79_groupi_n_197);
  not csa_tree_add_51_79_groupi_drc_bufs47587(csa_tree_add_51_79_groupi_n_197 ,csa_tree_add_51_79_groupi_n_3165);
  not csa_tree_add_51_79_groupi_drc_bufs47593(csa_tree_add_51_79_groupi_n_193 ,csa_tree_add_51_79_groupi_n_191);
  not csa_tree_add_51_79_groupi_drc_bufs47594(csa_tree_add_51_79_groupi_n_192 ,csa_tree_add_51_79_groupi_n_191);
  not csa_tree_add_51_79_groupi_drc_bufs47595(csa_tree_add_51_79_groupi_n_191 ,csa_tree_add_51_79_groupi_n_3190);
  not csa_tree_add_51_79_groupi_drc_bufs47601(csa_tree_add_51_79_groupi_n_187 ,csa_tree_add_51_79_groupi_n_185);
  not csa_tree_add_51_79_groupi_drc_bufs47602(csa_tree_add_51_79_groupi_n_186 ,csa_tree_add_51_79_groupi_n_185);
  not csa_tree_add_51_79_groupi_drc_bufs47603(csa_tree_add_51_79_groupi_n_185 ,csa_tree_add_51_79_groupi_n_3732);
  not csa_tree_add_51_79_groupi_drc_bufs47609(csa_tree_add_51_79_groupi_n_181 ,csa_tree_add_51_79_groupi_n_179);
  not csa_tree_add_51_79_groupi_drc_bufs47610(csa_tree_add_51_79_groupi_n_180 ,csa_tree_add_51_79_groupi_n_179);
  not csa_tree_add_51_79_groupi_drc_bufs47611(csa_tree_add_51_79_groupi_n_179 ,csa_tree_add_51_79_groupi_n_3177);
  not csa_tree_add_51_79_groupi_drc_bufs47617(csa_tree_add_51_79_groupi_n_175 ,csa_tree_add_51_79_groupi_n_173);
  not csa_tree_add_51_79_groupi_drc_bufs47618(csa_tree_add_51_79_groupi_n_174 ,csa_tree_add_51_79_groupi_n_173);
  not csa_tree_add_51_79_groupi_drc_bufs47619(csa_tree_add_51_79_groupi_n_173 ,csa_tree_add_51_79_groupi_n_3706);
  not csa_tree_add_51_79_groupi_drc_bufs47625(csa_tree_add_51_79_groupi_n_169 ,csa_tree_add_51_79_groupi_n_167);
  not csa_tree_add_51_79_groupi_drc_bufs47626(csa_tree_add_51_79_groupi_n_168 ,csa_tree_add_51_79_groupi_n_167);
  not csa_tree_add_51_79_groupi_drc_bufs47627(csa_tree_add_51_79_groupi_n_167 ,csa_tree_add_51_79_groupi_n_3707);
  not csa_tree_add_51_79_groupi_drc_bufs47633(csa_tree_add_51_79_groupi_n_163 ,csa_tree_add_51_79_groupi_n_161);
  not csa_tree_add_51_79_groupi_drc_bufs47634(csa_tree_add_51_79_groupi_n_162 ,csa_tree_add_51_79_groupi_n_161);
  not csa_tree_add_51_79_groupi_drc_bufs47635(csa_tree_add_51_79_groupi_n_161 ,csa_tree_add_51_79_groupi_n_3182);
  not csa_tree_add_51_79_groupi_drc_bufs47641(csa_tree_add_51_79_groupi_n_157 ,csa_tree_add_51_79_groupi_n_155);
  not csa_tree_add_51_79_groupi_drc_bufs47642(csa_tree_add_51_79_groupi_n_156 ,csa_tree_add_51_79_groupi_n_155);
  not csa_tree_add_51_79_groupi_drc_bufs47643(csa_tree_add_51_79_groupi_n_155 ,csa_tree_add_51_79_groupi_n_3170);
  not csa_tree_add_51_79_groupi_drc_bufs47649(csa_tree_add_51_79_groupi_n_151 ,csa_tree_add_51_79_groupi_n_149);
  not csa_tree_add_51_79_groupi_drc_bufs47650(csa_tree_add_51_79_groupi_n_150 ,csa_tree_add_51_79_groupi_n_149);
  not csa_tree_add_51_79_groupi_drc_bufs47651(csa_tree_add_51_79_groupi_n_149 ,csa_tree_add_51_79_groupi_n_3179);
  not csa_tree_add_51_79_groupi_drc_bufs47657(csa_tree_add_51_79_groupi_n_145 ,csa_tree_add_51_79_groupi_n_143);
  not csa_tree_add_51_79_groupi_drc_bufs47658(csa_tree_add_51_79_groupi_n_144 ,csa_tree_add_51_79_groupi_n_143);
  not csa_tree_add_51_79_groupi_drc_bufs47659(csa_tree_add_51_79_groupi_n_143 ,csa_tree_add_51_79_groupi_n_3730);
  not csa_tree_add_51_79_groupi_drc_bufs47665(csa_tree_add_51_79_groupi_n_139 ,csa_tree_add_51_79_groupi_n_137);
  not csa_tree_add_51_79_groupi_drc_bufs47666(csa_tree_add_51_79_groupi_n_138 ,csa_tree_add_51_79_groupi_n_137);
  not csa_tree_add_51_79_groupi_drc_bufs47667(csa_tree_add_51_79_groupi_n_137 ,csa_tree_add_51_79_groupi_n_3710);
  not csa_tree_add_51_79_groupi_drc_bufs47673(csa_tree_add_51_79_groupi_n_133 ,csa_tree_add_51_79_groupi_n_131);
  not csa_tree_add_51_79_groupi_drc_bufs47674(csa_tree_add_51_79_groupi_n_132 ,csa_tree_add_51_79_groupi_n_131);
  not csa_tree_add_51_79_groupi_drc_bufs47675(csa_tree_add_51_79_groupi_n_131 ,csa_tree_add_51_79_groupi_n_3183);
  not csa_tree_add_51_79_groupi_drc_bufs47681(csa_tree_add_51_79_groupi_n_127 ,csa_tree_add_51_79_groupi_n_125);
  not csa_tree_add_51_79_groupi_drc_bufs47682(csa_tree_add_51_79_groupi_n_126 ,csa_tree_add_51_79_groupi_n_125);
  not csa_tree_add_51_79_groupi_drc_bufs47683(csa_tree_add_51_79_groupi_n_125 ,csa_tree_add_51_79_groupi_n_3711);
  not csa_tree_add_51_79_groupi_drc_bufs47689(csa_tree_add_51_79_groupi_n_121 ,csa_tree_add_51_79_groupi_n_119);
  not csa_tree_add_51_79_groupi_drc_bufs47690(csa_tree_add_51_79_groupi_n_120 ,csa_tree_add_51_79_groupi_n_119);
  not csa_tree_add_51_79_groupi_drc_bufs47691(csa_tree_add_51_79_groupi_n_119 ,csa_tree_add_51_79_groupi_n_3723);
  not csa_tree_add_51_79_groupi_drc_bufs47697(csa_tree_add_51_79_groupi_n_115 ,csa_tree_add_51_79_groupi_n_113);
  not csa_tree_add_51_79_groupi_drc_bufs47698(csa_tree_add_51_79_groupi_n_114 ,csa_tree_add_51_79_groupi_n_113);
  not csa_tree_add_51_79_groupi_drc_bufs47699(csa_tree_add_51_79_groupi_n_113 ,csa_tree_add_51_79_groupi_n_3159);
  not csa_tree_add_51_79_groupi_drc_bufs47705(csa_tree_add_51_79_groupi_n_109 ,csa_tree_add_51_79_groupi_n_107);
  not csa_tree_add_51_79_groupi_drc_bufs47706(csa_tree_add_51_79_groupi_n_108 ,csa_tree_add_51_79_groupi_n_107);
  not csa_tree_add_51_79_groupi_drc_bufs47707(csa_tree_add_51_79_groupi_n_107 ,csa_tree_add_51_79_groupi_n_3184);
  not csa_tree_add_51_79_groupi_drc_bufs47713(csa_tree_add_51_79_groupi_n_103 ,csa_tree_add_51_79_groupi_n_101);
  not csa_tree_add_51_79_groupi_drc_bufs47714(csa_tree_add_51_79_groupi_n_102 ,csa_tree_add_51_79_groupi_n_101);
  not csa_tree_add_51_79_groupi_drc_bufs47715(csa_tree_add_51_79_groupi_n_101 ,csa_tree_add_51_79_groupi_n_3172);
  not csa_tree_add_51_79_groupi_drc_bufs47721(csa_tree_add_51_79_groupi_n_97 ,csa_tree_add_51_79_groupi_n_95);
  not csa_tree_add_51_79_groupi_drc_bufs47722(csa_tree_add_51_79_groupi_n_96 ,csa_tree_add_51_79_groupi_n_95);
  not csa_tree_add_51_79_groupi_drc_bufs47723(csa_tree_add_51_79_groupi_n_95 ,csa_tree_add_51_79_groupi_n_3712);
  not csa_tree_add_51_79_groupi_drc_bufs47729(csa_tree_add_51_79_groupi_n_91 ,csa_tree_add_51_79_groupi_n_89);
  not csa_tree_add_51_79_groupi_drc_bufs47730(csa_tree_add_51_79_groupi_n_90 ,csa_tree_add_51_79_groupi_n_89);
  not csa_tree_add_51_79_groupi_drc_bufs47731(csa_tree_add_51_79_groupi_n_89 ,csa_tree_add_51_79_groupi_n_3713);
  not csa_tree_add_51_79_groupi_drc_bufs47737(csa_tree_add_51_79_groupi_n_85 ,csa_tree_add_51_79_groupi_n_83);
  not csa_tree_add_51_79_groupi_drc_bufs47738(csa_tree_add_51_79_groupi_n_84 ,csa_tree_add_51_79_groupi_n_83);
  not csa_tree_add_51_79_groupi_drc_bufs47739(csa_tree_add_51_79_groupi_n_83 ,csa_tree_add_51_79_groupi_n_3186);
  not csa_tree_add_51_79_groupi_drc_bufs47745(csa_tree_add_51_79_groupi_n_79 ,csa_tree_add_51_79_groupi_n_77);
  not csa_tree_add_51_79_groupi_drc_bufs47746(csa_tree_add_51_79_groupi_n_78 ,csa_tree_add_51_79_groupi_n_77);
  not csa_tree_add_51_79_groupi_drc_bufs47747(csa_tree_add_51_79_groupi_n_77 ,csa_tree_add_51_79_groupi_n_3161);
  not csa_tree_add_51_79_groupi_drc_bufs47753(csa_tree_add_51_79_groupi_n_73 ,csa_tree_add_51_79_groupi_n_71);
  not csa_tree_add_51_79_groupi_drc_bufs47754(csa_tree_add_51_79_groupi_n_72 ,csa_tree_add_51_79_groupi_n_71);
  not csa_tree_add_51_79_groupi_drc_bufs47755(csa_tree_add_51_79_groupi_n_71 ,csa_tree_add_51_79_groupi_n_3163);
  not csa_tree_add_51_79_groupi_drc_bufs47761(csa_tree_add_51_79_groupi_n_67 ,csa_tree_add_51_79_groupi_n_65);
  not csa_tree_add_51_79_groupi_drc_bufs47762(csa_tree_add_51_79_groupi_n_66 ,csa_tree_add_51_79_groupi_n_65);
  not csa_tree_add_51_79_groupi_drc_bufs47763(csa_tree_add_51_79_groupi_n_65 ,csa_tree_add_51_79_groupi_n_3187);
  not csa_tree_add_51_79_groupi_drc_bufs47769(csa_tree_add_51_79_groupi_n_61 ,csa_tree_add_51_79_groupi_n_59);
  not csa_tree_add_51_79_groupi_drc_bufs47770(csa_tree_add_51_79_groupi_n_60 ,csa_tree_add_51_79_groupi_n_59);
  not csa_tree_add_51_79_groupi_drc_bufs47771(csa_tree_add_51_79_groupi_n_59 ,csa_tree_add_51_79_groupi_n_3173);
  not csa_tree_add_51_79_groupi_drc_bufs47777(csa_tree_add_51_79_groupi_n_55 ,csa_tree_add_51_79_groupi_n_53);
  not csa_tree_add_51_79_groupi_drc_bufs47778(csa_tree_add_51_79_groupi_n_54 ,csa_tree_add_51_79_groupi_n_53);
  not csa_tree_add_51_79_groupi_drc_bufs47779(csa_tree_add_51_79_groupi_n_53 ,csa_tree_add_51_79_groupi_n_3180);
  not csa_tree_add_51_79_groupi_drc_bufs47785(csa_tree_add_51_79_groupi_n_49 ,csa_tree_add_51_79_groupi_n_47);
  not csa_tree_add_51_79_groupi_drc_bufs47786(csa_tree_add_51_79_groupi_n_48 ,csa_tree_add_51_79_groupi_n_47);
  not csa_tree_add_51_79_groupi_drc_bufs47787(csa_tree_add_51_79_groupi_n_47 ,csa_tree_add_51_79_groupi_n_3722);
  not csa_tree_add_51_79_groupi_drc_bufs47789(csa_tree_add_51_79_groupi_n_46 ,csa_tree_add_51_79_groupi_n_44);
  not csa_tree_add_51_79_groupi_drc_bufs47790(csa_tree_add_51_79_groupi_n_45 ,csa_tree_add_51_79_groupi_n_44);
  not csa_tree_add_51_79_groupi_drc_bufs47791(csa_tree_add_51_79_groupi_n_44 ,csa_tree_add_51_79_groupi_n_3731);
  xor csa_tree_add_51_79_groupi_g2(csa_tree_add_51_79_groupi_n_43 ,csa_tree_add_51_79_groupi_n_11042 ,csa_tree_add_51_79_groupi_n_11085);
  xor csa_tree_add_51_79_groupi_g47793(csa_tree_add_51_79_groupi_n_42 ,csa_tree_add_51_79_groupi_n_10987 ,csa_tree_add_51_79_groupi_n_10994);
  xor csa_tree_add_51_79_groupi_g47794(csa_tree_add_51_79_groupi_n_41 ,csa_tree_add_51_79_groupi_n_10940 ,csa_tree_add_51_79_groupi_n_10989);
  xor csa_tree_add_51_79_groupi_g47795(csa_tree_add_51_79_groupi_n_40 ,csa_tree_add_51_79_groupi_n_10939 ,csa_tree_add_51_79_groupi_n_37);
  xor csa_tree_add_51_79_groupi_g47796(csa_tree_add_51_79_groupi_n_39 ,csa_tree_add_51_79_groupi_n_10937 ,csa_tree_add_51_79_groupi_n_10944);
  xor csa_tree_add_51_79_groupi_g47797(csa_tree_add_51_79_groupi_n_38 ,csa_tree_add_51_79_groupi_n_10721 ,csa_tree_add_51_79_groupi_n_10929);
  xor csa_tree_add_51_79_groupi_g47798(csa_tree_add_51_79_groupi_n_37 ,csa_tree_add_51_79_groupi_n_10720 ,csa_tree_add_51_79_groupi_n_10832);
  xor csa_tree_add_51_79_groupi_g47799(csa_tree_add_51_79_groupi_n_36 ,csa_tree_add_51_79_groupi_n_10789 ,csa_tree_add_51_79_groupi_n_10801);
  xor csa_tree_add_51_79_groupi_g47800(csa_tree_add_51_79_groupi_n_35 ,csa_tree_add_51_79_groupi_n_10725 ,csa_tree_add_51_79_groupi_n_10763);
  xor csa_tree_add_51_79_groupi_g47801(csa_tree_add_51_79_groupi_n_34 ,csa_tree_add_51_79_groupi_n_10519 ,csa_tree_add_51_79_groupi_n_10281);
  xor csa_tree_add_51_79_groupi_g47802(csa_tree_add_51_79_groupi_n_33 ,csa_tree_add_51_79_groupi_n_9609 ,csa_tree_add_51_79_groupi_n_9646);
  xor csa_tree_add_51_79_groupi_g47803(csa_tree_add_51_79_groupi_n_32 ,csa_tree_add_51_79_groupi_n_9206 ,csa_tree_add_51_79_groupi_n_9413);
  xor csa_tree_add_51_79_groupi_g47804(csa_tree_add_51_79_groupi_n_31 ,csa_tree_add_51_79_groupi_n_8967 ,csa_tree_add_51_79_groupi_n_9411);
  xor csa_tree_add_51_79_groupi_g47805(csa_tree_add_51_79_groupi_n_30 ,csa_tree_add_51_79_groupi_n_8571 ,csa_tree_add_51_79_groupi_n_8657);
  and csa_tree_add_51_79_groupi_g47806(csa_tree_add_51_79_groupi_n_29 ,csa_tree_add_51_79_groupi_n_1530 ,csa_tree_add_51_79_groupi_n_7211);
  xor csa_tree_add_51_79_groupi_g47807(csa_tree_add_51_79_groupi_n_28 ,csa_tree_add_51_79_groupi_n_6757 ,csa_tree_add_51_79_groupi_n_6935);
  xor csa_tree_add_51_79_groupi_g47808(csa_tree_add_51_79_groupi_n_27 ,csa_tree_add_51_79_groupi_n_6834 ,csa_tree_add_51_79_groupi_n_6921);
  xor csa_tree_add_51_79_groupi_g47809(csa_tree_add_51_79_groupi_n_26 ,csa_tree_add_51_79_groupi_n_6760 ,csa_tree_add_51_79_groupi_n_8028);
  xnor csa_tree_add_51_79_groupi_g47810(csa_tree_add_51_79_groupi_n_25 ,csa_tree_add_51_79_groupi_n_5107 ,csa_tree_add_51_79_groupi_n_3320);
  xor csa_tree_add_51_79_groupi_g47811(csa_tree_add_51_79_groupi_n_24 ,csa_tree_add_51_79_groupi_n_5097 ,csa_tree_add_51_79_groupi_n_5517);
  xor csa_tree_add_51_79_groupi_g47812(csa_tree_add_51_79_groupi_n_23 ,csa_tree_add_51_79_groupi_n_4301 ,csa_tree_add_51_79_groupi_n_5579);
  xor csa_tree_add_51_79_groupi_g47813(csa_tree_add_51_79_groupi_n_22 ,csa_tree_add_51_79_groupi_n_4299 ,csa_tree_add_51_79_groupi_n_5586);
  xor csa_tree_add_51_79_groupi_g47814(csa_tree_add_51_79_groupi_n_21 ,csa_tree_add_51_79_groupi_n_4298 ,csa_tree_add_51_79_groupi_n_5594);
  xor csa_tree_add_51_79_groupi_g47815(csa_tree_add_51_79_groupi_n_20 ,csa_tree_add_51_79_groupi_n_4297 ,csa_tree_add_51_79_groupi_n_5588);
  xor csa_tree_add_51_79_groupi_g47816(csa_tree_add_51_79_groupi_n_19 ,csa_tree_add_51_79_groupi_n_4296 ,csa_tree_add_51_79_groupi_n_5580);
  xor csa_tree_add_51_79_groupi_g47817(csa_tree_add_51_79_groupi_n_18 ,csa_tree_add_51_79_groupi_n_4295 ,csa_tree_add_51_79_groupi_n_5583);
  xor csa_tree_add_51_79_groupi_g47818(csa_tree_add_51_79_groupi_n_17 ,csa_tree_add_51_79_groupi_n_4294 ,csa_tree_add_51_79_groupi_n_5582);
  xor csa_tree_add_51_79_groupi_g47819(csa_tree_add_51_79_groupi_n_16 ,csa_tree_add_51_79_groupi_n_4293 ,csa_tree_add_51_79_groupi_n_5585);
  xor csa_tree_add_51_79_groupi_g47820(csa_tree_add_51_79_groupi_n_15 ,csa_tree_add_51_79_groupi_n_4291 ,csa_tree_add_51_79_groupi_n_5584);
  xor csa_tree_add_51_79_groupi_g47821(csa_tree_add_51_79_groupi_n_14 ,csa_tree_add_51_79_groupi_n_4290 ,csa_tree_add_51_79_groupi_n_5578);
  xor csa_tree_add_51_79_groupi_g47822(csa_tree_add_51_79_groupi_n_13 ,csa_tree_add_51_79_groupi_n_4289 ,csa_tree_add_51_79_groupi_n_5581);
  xor csa_tree_add_51_79_groupi_g47823(csa_tree_add_51_79_groupi_n_12 ,csa_tree_add_51_79_groupi_n_4288 ,csa_tree_add_51_79_groupi_n_5587);
  xor csa_tree_add_51_79_groupi_g47824(csa_tree_add_51_79_groupi_n_11 ,csa_tree_add_51_79_groupi_n_3735 ,csa_tree_add_51_79_groupi_n_3273);
  xor csa_tree_add_51_79_groupi_g47825(csa_tree_add_51_79_groupi_n_10 ,csa_tree_add_51_79_groupi_n_3256 ,csa_tree_add_51_79_groupi_n_6181);
  xor csa_tree_add_51_79_groupi_g47826(csa_tree_add_51_79_groupi_n_9 ,csa_tree_add_51_79_groupi_n_3239 ,csa_tree_add_51_79_groupi_n_6333);
  xor csa_tree_add_51_79_groupi_g47827(csa_tree_add_51_79_groupi_n_8 ,csa_tree_add_51_79_groupi_n_4 ,csa_tree_add_51_79_groupi_n_1777);
  xor csa_tree_add_51_79_groupi_g47828(csa_tree_add_51_79_groupi_n_7 ,csa_tree_add_51_79_groupi_n_3282 ,csa_tree_add_51_79_groupi_n_1776);
  xor csa_tree_add_51_79_groupi_g47829(csa_tree_add_51_79_groupi_n_6 ,csa_tree_add_51_79_groupi_n_5 ,csa_tree_add_51_79_groupi_n_1775);
  xor csa_tree_add_51_79_groupi_g47830(csa_tree_add_51_79_groupi_n_5 ,csa_tree_add_51_79_groupi_n_1787 ,csa_tree_add_51_79_groupi_n_1774);
  xor csa_tree_add_51_79_groupi_g47831(csa_tree_add_51_79_groupi_n_4 ,csa_tree_add_51_79_groupi_n_1781 ,csa_tree_add_51_79_groupi_n_1722);
  xor csa_tree_add_51_79_groupi_g47832(csa_tree_add_51_79_groupi_n_3 ,csa_tree_add_51_79_groupi_n_1783 ,csa_tree_add_51_79_groupi_n_1721);
  xor csa_tree_add_51_79_groupi_g47833(csa_tree_add_51_79_groupi_n_2 ,csa_tree_add_51_79_groupi_n_3 ,csa_tree_add_51_79_groupi_n_1720);
  xor csa_tree_add_51_79_groupi_g47834(csa_tree_add_51_79_groupi_n_1 ,csa_tree_add_51_79_groupi_n_1210 ,csa_tree_add_51_79_groupi_n_4811);
  xor csa_tree_add_51_79_groupi_g47835(csa_tree_add_51_79_groupi_n_0 ,csa_tree_add_51_79_groupi_n_6161 ,csa_tree_add_51_79_groupi_n_764);
  buf g47848(csa_tree_add_51_79_groupi_n_1905 ,in11[0]);
  buf g47849(csa_tree_add_51_79_groupi_n_2337 ,in3[0]);
  buf g47850(csa_tree_add_51_79_groupi_n_2326 ,in19[0]);
  buf g47851(csa_tree_add_51_79_groupi_n_2344 ,in1[0]);
  buf g47852(csa_tree_add_51_79_groupi_n_1852 ,in9[0]);

endmodule

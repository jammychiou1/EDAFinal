module top(in1, in2, in3, in4, out1, out2, out3, out4);

  input [33:0] in1;

  input [34:0] in2, in3, in4;

  output out1, out2, out3, out4;
  wire [33:0] in1;
  wire [34:0] in2, in3, in4;
  wire out1, out2, out3, out4;
  wire w__1, w__2, w__3, w__4, w__5, w__6, w__7, w__8;
  wire w__9, w__10, w__12, w__12, w__13, w__14, w__15, w__16;
  wire w__17, w__18, w__19, w__20, w__683, w__22, w__23, w__24;
  wire w__25, w__26, w__27, w__28, w__29, w__30, w__31, w__32;
  wire w__33, w__34, w__35, w__36, w__37, w__38, w__39, w__40;
  wire w__41, w__42, w__43, w__44, w__45, w__46, w__47, w__48;
  wire w__49, w__50, w__51, w__52, w__53, w__54, w__55, w__56;
  wire w__57, w__58, w__59, w__60, w__61, w__62, w__63, w__64;
  wire w__65, w__66, w__67, w__68, w__69, w__70, w__71, w__72;
  wire w__73, w__74, w__75, w__76, w__77, w__78, w__79, w__80;
  wire w__81, w__82, w__83, w__84, w__85, w__86, w__87, w__88;
  wire w__89, w__90, w__91, w__92, w__93, w__94, w__95, w__96;
  wire w__97, w__98, w__99, w__100, w__101, w__102, w__103, w__104;
  wire w__105, w__106, w__107, w__108, w__109, w__110, w__111, w__112;
  wire w__113, w__114, w__115, w__116, w__117, w__118, w__119, w__120;
  wire w__121, w__122, w__123, w__124, w__125, w__126, w__127, w__128;
  wire w__129, w__130, w__131, w__132, w__133, w__134, w__135, w__136;
  wire w__137, w__138, w__479, w__480, w__493, w__494, w__491, w__492;
  wire w__485, w__486, w__495, w__496, w__497, w__498, w__487, w__488;
  wire w__489, w__490, w__527, w__519, w__515, w__529, w__501, w__533;
  wire w__541, w__523, w__543, w__531, w__513, w__499, w__503, w__535;
  wire w__539, w__521, w__517, w__507, w__511, w__537, w__509, w__525;
  wire w__505, w__178, w__179, w__180, w__181, w__182, w__183, w__481;
  wire w__185, w__186, w__483, w__188, w__189, w__190, w__191, w__192;
  wire w__193, w__194, w__195, w__196, w__197, w__198, w__199, w__200;
  wire w__201, w__202, w__203, w__204, w__205, w__206, w__207, w__208;
  wire w__209, w__210, w__211, w__212, w__213, w__214, w__215, w__216;
  wire w__217, w__218, w__219, w__220, w__221, w__222, w__223, w__224;
  wire w__225, w__226, w__227, w__228, w__229, w__230, w__231, w__232;
  wire w__233, w__234, w__235, w__236, w__237, w__238, w__239, w__240;
  wire w__241, w__242, w__243, w__244, w__245, w__246, w__247, w__248;
  wire w__249, w__250, w__251, w__252, w__253, w__254, w__255, w__256;
  wire w__257, w__258, w__259, w__260, w__261, w__262, w__263, w__264;
  wire w__265, w__266, w__267, w__268, w__269, w__270, w__271, w__272;
  wire w__273, w__274, w__275, w__276, w__277, w__278, w__279, w__280;
  wire w__281, w__282, w__283, w__284, w__285, w__286, w__287, w__288;
  wire w__289, w__290, w__291, w__292, w__293, w__294, w__295, w__296;
  wire w__297, w__298, w__299, w__300, w__301, w__302, w__303, w__304;
  wire w__305, w__306, w__307, w__308, w__309, w__310, w__311, w__312;
  wire w__313, w__314, w__315, w__316, w__317, w__318, w__319, w__320;
  wire w__321, w__322, w__323, w__324, w__325, w__326, w__327, w__328;
  wire w__329, w__330, w__331, w__332, w__333, w__334, w__335, w__336;
  wire w__337, w__338, w__339, w__340, w__341, w__342, w__343, w__344;
  wire w__345, w__346, w__347, w__348, w__349, w__350, w__351, w__352;
  wire w__353, w__354, w__355, w__356, w__357, w__358, w__359, w__360;
  wire w__361, w__362, w__363, w__364, w__365, w__366, w__367, w__368;
  wire w__369, w__370, w__371, w__372, w__373, w__374, w__375, w__376;
  wire w__377, w__378, w__379, w__380, w__381, w__382, w__383, w__384;
  wire w__385, w__386, w__387, w__388, w__389, w__390, w__391, w__392;
  wire w__393, w__394, w__395, w__396, w__397, w__398, w__399, w__400;
  wire w__401, w__402, w__403, w__404, w__405, w__406, w__407, w__408;
  wire w__409, w__410, w__411, w__412, w__413, w__414, w__415, w__416;
  wire w__417, w__418, w__419, w__420, w__421, w__422, w__423, w__424;
  wire w__425, w__426, w__427, w__428, w__429, w__430, w__431, w__432;
  wire w__433, w__434, w__435, w__436, w__437, w__438, w__439, w__440;
  wire w__441, w__442, w__443, w__444, w__445, w__446, w__447, w__448;
  wire w__449, w__450, w__451, w__452, w__453, w__454, w__455, w__456;
  wire w__457, w__458, w__459, w__460, w__461, w__462, w__463, w__464;
  wire w__465, w__466, w__467, w__468, w__469, w__470, w__471, w__472;
  wire w__473, w__474, w__475, w__476, w__477, w__478, w__479, w__480;
  wire w__481, w__482, w__483, w__484, w__485, w__486, w__487, w__488;
  wire w__489, w__490, w__491, w__492, w__493, w__494, w__495, w__496;
  wire w__497, w__498, w__499, w__500, w__501, w__502, w__503, w__504;
  wire w__505, w__506, w__507, w__508, w__509, w__510, w__511, w__512;
  wire w__513, w__514, w__515, w__516, w__517, w__518, w__519, w__520;
  wire w__521, w__522, w__523, w__524, w__525, w__526, w__527, w__528;
  wire w__529, w__530, w__531, w__532, w__533, w__534, w__535, w__536;
  wire w__537, w__538, w__539, w__540, w__541, w__542, w__543, w__544;
  wire w__545, w__546, w__547, w__548, w__549, w__550, w__551, w__552;
  wire w__553, w__554, w__555, w__556, w__557, w__558, w__559, w__560;
  wire w__561, w__562, w__563, w__564, w__565, w__566, w__567, w__568;
  wire w__569, w__570, w__571, w__572, w__573, w__574, w__575, w__576;
  wire w__577, w__578, w__579, w__580, w__581, w__582, w__583, w__584;
  wire w__585, w__586, w__587, w__588, w__589, w__590, w__591, w__592;
  wire w__593, w__594, w__595, w__596, w__597, w__598, w__599, w__600;
  wire w__601, w__602, w__603, w__604, w__605, w__606, w__607, w__608;
  wire w__609, w__610, w__611, w__612, w__613, w__614, w__615, w__616;
  wire w__617, w__618, w__619, w__620, w__621, w__622, w__623, w__624;
  wire w__625, w__626, w__627, w__628, w__629, w__630, w__631, w__632;
  wire w__633, w__634, w__635, w__636, w__637, w__638, w__639, w__640;
  wire w__641, w__642, w__643, w__644, w__645, w__646, w__647, w__648;
  wire w__649, w__650, w__651, w__652, w__653, w__654, w__655, w__656;
  wire w__657, w__658, w__659, w__660, w__661, w__662, w__663, w__664;
  wire w__665, w__666, w__667, w__668, w__669, w__670, w__671, w__672;
  wire w__673, w__674, w__675, w__676, w__677, w__678, w__679, w__680;
  wire w__681, w__682, w__683, w__684, w__685, w__686, w__687, w__688;
  wire w__689, w__690, w__691, w__692, w__693, w__694, w__695, w__696;
  wire w__697, w__698, w__699, w__700, w__701, w__702, w__703, w__704;
  wire w__705, w__706, w__707, w__708, w__709, w__710, w__711, w__712;
  wire w__713, w__714, w__715, w__716, w__717;
  not g__1(w__683 ,in1[0]);
  nor g__2(w__682 ,w__672 ,w__680);
  nor g__3(w__681 ,w__669 ,w__679);
  or g__4(w__680 ,w__668 ,w__677);
  or g__5(w__679 ,w__667 ,w__678);
  or g__6(w__678 ,w__664 ,w__676);
  or g__7(w__677 ,w__655 ,w__675);
  or g__8(w__676 ,w__673 ,w__671);
  or g__9(w__675 ,w__670 ,w__674);
  or g__10(w__674 ,w__660 ,w__666);
  or g__11(w__673 ,w__662 ,w__661);
  or g__12(w__672 ,w__656 ,w__654);
  or g__13(w__671 ,w__659 ,w__649);
  or g__14(w__670 ,w__650 ,w__658);
  or g__15(w__669 ,w__652 ,w__651);
  or g__16(w__668 ,w__653 ,w__663);
  or g__17(w__667 ,w__657 ,w__665);
  or g__18(w__666 ,w__627 ,w__626);
  or g__19(w__665 ,w__646 ,w__644);
  or g__20(w__664 ,w__548 ,w__640);
  or g__21(w__663 ,w__641 ,w__636);
  or g__22(w__662 ,w__638 ,w__637);
  or g__23(w__661 ,w__635 ,w__633);
  or g__24(w__660 ,w__634 ,w__629);
  or g__25(w__659 ,w__632 ,w__631);
  or g__26(w__658 ,w__645 ,w__639);
  or g__27(w__657 ,w__615 ,w__648);
  or g__28(w__656 ,w__643 ,w__620);
  or g__29(w__655 ,w__546 ,w__623);
  or g__30(w__654 ,w__625 ,w__642);
  or g__31(w__653 ,w__624 ,w__616);
  or g__32(w__652 ,w__622 ,w__621);
  or g__33(w__651 ,w__619 ,w__617);
  or g__34(w__650 ,w__618 ,w__647);
  or g__35(w__649 ,w__630 ,w__628);
  or g__36(w__648 ,w__609 ,w__608);
  or g__37(w__647 ,w__610 ,w__607);
  or g__38(w__646 ,w__606 ,w__605);
  or g__39(w__645 ,w__602 ,w__599);
  or g__40(w__644 ,w__603 ,w__601);
  or g__41(w__643 ,w__587 ,w__583);
  or g__42(w__642 ,w__594 ,w__576);
  or g__43(w__641 ,w__596 ,w__588);
  or g__44(w__640 ,w__598 ,w__597);
  or g__45(w__639 ,w__595 ,w__591);
  or g__46(w__638 ,w__593 ,w__592);
  or g__47(w__637 ,w__590 ,w__589);
  or g__48(w__636 ,w__578 ,w__569);
  or g__49(w__635 ,w__586 ,w__584);
  or g__50(w__634 ,w__585 ,w__582);
  or g__51(w__633 ,w__581 ,w__614);
  or g__52(w__632 ,w__577 ,w__575);
  or g__53(w__631 ,w__573 ,w__572);
  or g__54(w__630 ,w__600 ,w__570);
  or g__55(w__629 ,w__574 ,w__571);
  or g__56(w__628 ,w__547 ,w__567);
  or g__57(w__627 ,w__568 ,w__566);
  or g__58(w__626 ,w__579 ,w__565);
  or g__59(w__625 ,w__557 ,w__611);
  or g__60(w__624 ,w__563 ,w__555);
  or g__61(w__623 ,w__564 ,w__560);
  or g__62(w__622 ,w__562 ,w__561);
  or g__63(w__621 ,w__559 ,w__558);
  or g__64(w__620 ,w__580 ,w__545);
  or g__65(w__619 ,w__556 ,w__554);
  or g__66(w__618 ,w__553 ,w__550);
  or g__67(w__617 ,w__552 ,w__551);
  or g__68(w__616 ,w__613 ,w__604);
  or g__69(w__615 ,w__549 ,w__612);
  xor g__70(w__614 ,w__524 ,in4[8]);
  xor g__71(w__613 ,w__496 ,in3[21]);
  xor g__72(w__612 ,w__482 ,in4[22]);
  xor g__73(w__611 ,w__540 ,in3[26]);
  xor g__74(w__610 ,w__528 ,in3[13]);
  xor g__75(w__609 ,w__496 ,in4[21]);
  xor g__76(w__608 ,w__514 ,in4[20]);
  xor g__77(w__607 ,w__526 ,in3[12]);
  xor g__78(w__606 ,w__538 ,in4[19]);
  xor g__79(w__605 ,w__498 ,in4[18]);
  xor g__80(w__604 ,w__514 ,in3[20]);
  xor g__81(w__603 ,w__536 ,in4[17]);
  xor g__82(w__602 ,w__520 ,in3[11]);
  xor g__83(w__601 ,w__488 ,in4[16]);
  xor g__84(w__600 ,w__508 ,in4[3]);
  xor g__85(w__599 ,w__518 ,in3[10]);
  xor g__86(w__598 ,w__490 ,in4[33]);
  xor g__87(w__597 ,w__502 ,in4[32]);
  xor g__88(w__596 ,w__538 ,in3[19]);
  xor g__89(w__595 ,w__516 ,in3[9]);
  xor g__90(w__594 ,w__534 ,in3[25]);
  xor g__91(w__593 ,w__504 ,in4[15]);
  xor g__92(w__592 ,w__532 ,in4[14]);
  xor g__93(w__591 ,w__524 ,in3[8]);
  xor g__94(w__590 ,w__528 ,in4[13]);
  xor g__95(w__589 ,w__526 ,in4[12]);
  xor g__96(w__588 ,w__498 ,in3[18]);
  xor g__97(w__587 ,w__494 ,in3[31]);
  xor g__98(w__586 ,w__520 ,in4[11]);
  xor g__99(w__585 ,w__506 ,in3[7]);
  xor g__100(w__584 ,w__518 ,in4[10]);
  xor g__101(w__583 ,w__480 ,in3[30]);
  xor g__102(w__582 ,w__512 ,in3[6]);
  xor g__103(w__581 ,w__516 ,in4[9]);
  xor g__104(w__580 ,w__544 ,in3[29]);
  xnor g__105(w__579 ,in1[0] ,in3[0]);
  xor g__106(w__578 ,w__536 ,in3[17]);
  xor g__107(w__577 ,w__506 ,in4[7]);
  xor g__108(w__576 ,w__530 ,in3[24]);
  xor g__109(w__575 ,w__512 ,in4[6]);
  xor g__110(w__574 ,w__510 ,in3[5]);
  xor g__111(w__573 ,w__510 ,in4[5]);
  xor g__112(w__572 ,w__484 ,in4[4]);
  xor g__113(w__571 ,w__484 ,in3[4]);
  xor g__114(w__570 ,w__486 ,in4[2]);
  xor g__115(w__569 ,w__488 ,in3[16]);
  xor g__116(w__568 ,w__508 ,in3[3]);
  xor g__117(w__567 ,w__478 ,in4[1]);
  xor g__118(w__566 ,w__486 ,in3[2]);
  xor g__119(w__565 ,w__478 ,in3[1]);
  xor g__120(w__564 ,w__500 ,in3[34]);
  xor g__121(w__563 ,w__522 ,in3[23]);
  xor g__122(w__562 ,w__494 ,in4[31]);
  xor g__123(w__561 ,w__480 ,in4[30]);
  xor g__124(w__560 ,w__490 ,in3[33]);
  xor g__125(w__559 ,w__544 ,in4[29]);
  xor g__126(w__558 ,w__492 ,in4[28]);
  xor g__127(w__557 ,w__542 ,in3[27]);
  xor g__128(w__556 ,w__542 ,in4[27]);
  xor g__129(w__555 ,w__482 ,in3[22]);
  xor g__130(w__554 ,w__540 ,in4[26]);
  xor g__131(w__553 ,w__504 ,in3[15]);
  xor g__132(w__552 ,w__534 ,in4[25]);
  xor g__133(w__551 ,w__530 ,in4[24]);
  xor g__134(w__550 ,w__532 ,in3[14]);
  xor g__135(w__549 ,w__522 ,in4[23]);
  xor g__136(w__548 ,w__500 ,in4[34]);
  xnor g__137(w__547 ,in1[0] ,in4[0]);
  xor g__138(w__546 ,w__502 ,in3[32]);
  xor g__139(w__545 ,w__492 ,in3[28]);
  not g__140(w__544 ,w__543);
  not g__141(w__543 ,w__712);
  not g__142(w__542 ,w__541);
  not g__143(w__541 ,w__710);
  not g__144(w__540 ,w__539);
  not g__145(w__539 ,w__709);
  not g__146(w__538 ,w__537);
  not g__147(w__537 ,w__702);
  not g__148(w__536 ,w__535);
  not g__149(w__535 ,w__700);
  not g__150(w__534 ,w__533);
  not g__151(w__533 ,w__708);
  not g__152(w__532 ,w__531);
  not g__153(w__531 ,w__697);
  not g__154(w__530 ,w__529);
  not g__155(w__529 ,w__707);
  not g__156(w__528 ,w__527);
  not g__157(w__527 ,w__696);
  not g__158(w__526 ,w__525);
  not g__159(w__525 ,w__695);
  not g__160(w__524 ,w__523);
  not g__161(w__523 ,w__691);
  not g__162(w__522 ,w__521);
  not g__163(w__521 ,w__706);
  not g__164(w__520 ,w__519);
  not g__165(w__519 ,w__694);
  not g__166(w__518 ,w__517);
  not g__167(w__517 ,w__693);
  not g__168(w__516 ,w__515);
  not g__169(w__515 ,w__692);
  not g__170(w__514 ,w__513);
  not g__171(w__513 ,w__703);
  not g__172(w__512 ,w__511);
  not g__173(w__511 ,w__689);
  not g__174(w__510 ,w__509);
  not g__175(w__509 ,w__688);
  not g__176(w__508 ,w__507);
  not g__177(w__507 ,w__686);
  not g__178(w__506 ,w__505);
  not g__179(w__505 ,w__690);
  not g__180(w__504 ,w__503);
  not g__181(w__503 ,w__698);
  not g__182(w__502 ,w__501);
  not g__183(w__501 ,w__715);
  not g__184(w__500 ,w__499);
  not g__185(w__499 ,w__717);
  not g__186(w__498 ,w__497);
  not g__187(w__497 ,w__701);
  not g__188(w__496 ,w__495);
  not g__189(w__495 ,w__704);
  not g__190(w__494 ,w__493);
  not g__191(w__493 ,w__714);
  not g__192(w__492 ,w__491);
  not g__193(w__491 ,w__711);
  not g__194(w__490 ,w__489);
  not g__195(w__489 ,w__716);
  not g__196(w__488 ,w__487);
  not g__197(w__487 ,w__699);
  not g__198(w__486 ,w__485);
  not g__199(w__485 ,w__685);
  not g__200(w__484 ,w__483);
  not g__201(w__483 ,w__687);
  not g__202(w__482 ,w__481);
  not g__203(w__481 ,w__705);
  not g__204(w__480 ,w__479);
  not g__205(w__479 ,w__713);
  not g__206(w__478 ,w__477);
  not g__207(w__477 ,w__684);
  buf g__208(out3 ,w__681);
  buf g__209(out2 ,w__682);
  and g__210(w__115 ,w__23 ,w__112);
  or g__211(w__114 ,w__113 ,w__112);
  and g__212(w__113 ,in1[32] ,w__111);
  and g__213(w__112 ,w__15 ,w__110);
  not g__214(w__111 ,w__110);
  and g__215(w__110 ,w__18 ,w__104);
  or g__216(w__109 ,w__105 ,w__104);
  xnor g__217(w__108 ,w__95 ,in1[29]);
  xnor g__218(w__107 ,w__94 ,in1[27]);
  xnor g__219(w__106 ,w__93 ,in1[23]);
  and g__220(w__105 ,in1[30] ,w__97);
  and g__221(w__104 ,w__22 ,w__96);
  xnor g__222(w__103 ,w__87 ,in1[28]);
  xnor g__223(w__102 ,w__89 ,in1[26]);
  xnor g__224(w__101 ,w__85 ,in1[22]);
  xnor g__225(w__100 ,w__88 ,in1[25]);
  xnor g__226(w__99 ,w__84 ,in1[21]);
  xnor g__227(w__98 ,w__83 ,in1[19]);
  not g__228(w__97 ,w__96);
  and g__229(w__96 ,w__26 ,w__86);
  or g__230(w__95 ,in1[28] ,w__87);
  or g__231(w__94 ,in1[26] ,w__89);
  or g__232(w__93 ,in1[22] ,w__85);
  xnor g__233(w__92 ,w__80 ,in1[20]);
  xnor g__234(w__91 ,w__79 ,in1[18]);
  xnor g__235(w__90 ,w__81 ,in1[17]);
  or g__236(w__89 ,w__34 ,w__7);
  or g__237(w__88 ,in1[24] ,w__7);
  not g__238(w__87 ,w__86);
  and g__239(w__86 ,w__44 ,w__78);
  or g__240(w__85 ,w__28 ,w__80);
  or g__241(w__84 ,in1[20] ,w__80);
  or g__242(w__83 ,in1[18] ,w__79);
  xnor g__243(w__82 ,w__12 ,in1[16]);
  or g__244(w__81 ,in1[16] ,w__12);
  or g__245(w__80 ,w__41 ,w__12);
  or g__246(w__79 ,w__30 ,w__12);
  and g__247(w__78 ,w__54 ,w__76);
  or g__248(w__77 ,w__74 ,w__76);
  not g__249(w__75 ,w__76);
  and g__250(w__76 ,w__13 ,w__71);
  nor g__251(w__74 ,w__13 ,w__71);
  xnor g__252(w__73 ,w__66 ,in1[11]);
  xnor g__253(w__72 ,w__67 ,in1[13]);
  and g__254(w__71 ,w__16 ,w__65);
  xnor g__255(w__70 ,w__61 ,in1[12]);
  xnor g__256(w__69 ,w__62 ,in1[10]);
  xnor g__257(w__68 ,w__63 ,in1[9]);
  or g__258(w__67 ,in1[12] ,w__61);
  or g__259(w__66 ,in1[10] ,w__62);
  and g__260(w__65 ,w__32 ,w__60);
  xnor g__261(w__64 ,w__56 ,in1[8]);
  or g__262(w__63 ,in1[8] ,w__9);
  or g__263(w__62 ,w__27 ,w__9);
  not g__264(w__61 ,w__60);
  and g__265(w__60 ,w__45 ,w__57);
  or g__266(w__59 ,w__58 ,w__57);
  and g__267(w__58 ,in1[7] ,w__53);
  not g__268(w__56 ,w__57);
  and g__269(w__57 ,w__17 ,w__52);
  xnor g__270(w__55 ,w__50 ,in1[5]);
  nor g__271(w__54 ,w__29 ,w__49);
  not g__272(w__53 ,w__52);
  and g__273(w__52 ,w__14 ,w__48);
  xnor g__274(w__51 ,w__42 ,in1[4]);
  or g__275(w__50 ,in1[4] ,w__42);
  or g__276(w__49 ,w__28 ,w__41);
  and g__277(w__48 ,w__25 ,w__43);
  or g__278(w__47 ,w__46 ,w__43);
  and g__279(w__46 ,in1[3] ,w__39);
  nor g__280(w__45 ,in1[10] ,w__37);
  nor g__281(w__44 ,in1[26] ,w__36);
  not g__282(w__42 ,w__43);
  and g__283(w__43 ,w__20 ,w__38);
  or g__284(w__41 ,in1[18] ,w__40);
  or g__285(w__40 ,in1[19] ,w__30);
  not g__286(w__39 ,w__38);
  and g__287(w__38 ,w__24 ,w__31);
  or g__288(w__37 ,in1[11] ,w__27);
  or g__289(w__36 ,in1[27] ,w__34);
  or g__290(w__35 ,w__33 ,w__31);
  or g__291(w__34 ,in1[25] ,in1[24]);
  and g__292(w__33 ,in1[1] ,in1[0]);
  nor g__293(w__32 ,in1[13] ,in1[12]);
  and g__294(w__31 ,w__19 ,w__683);
  or g__295(w__30 ,in1[17] ,in1[16]);
  or g__296(w__29 ,in1[23] ,in1[22]);
  or g__297(w__28 ,in1[21] ,in1[20]);
  or g__298(w__27 ,in1[9] ,in1[8]);
  nor g__299(w__26 ,in1[29] ,in1[28]);
  nor g__300(w__25 ,in1[5] ,in1[4]);
  not g__301(w__24 ,in1[2]);
  not g__302(w__23 ,in1[33]);
  not g__303(w__22 ,in1[30]);
  not g__305(w__20 ,in1[3]);
  not g__306(w__19 ,in1[1]);
  not g__307(w__18 ,in1[31]);
  not g__308(w__17 ,in1[7]);
  not g__309(w__16 ,in1[14]);
  not g__310(w__15 ,in1[32]);
  not g__311(w__14 ,in1[6]);
  not g__312(w__13 ,in1[15]);
  not g__313(w__12 ,w__10);
  not g__315(w__10 ,w__75);
  not g__316(w__9 ,w__8);
  not g__317(w__8 ,w__56);
  buf g__318(w__685 ,w__1);
  buf g__319(w__716 ,w__6);
  buf g__320(w__687 ,w__51);
  buf g__321(w__706 ,w__106);
  buf g__322(w__701 ,w__91);
  buf g__323(w__703 ,w__92);
  buf g__324(w__689 ,w__2);
  buf g__325(w__691 ,w__64);
  buf g__326(w__692 ,w__68);
  buf g__327(w__693 ,w__69);
  buf g__328(w__695 ,w__70);
  buf g__329(w__688 ,w__55);
  buf g__330(w__707 ,w__4);
  buf g__331(w__697 ,w__3);
  buf g__332(w__705 ,w__101);
  buf g__333(w__711 ,w__103);
  buf g__334(w__700 ,w__90);
  buf g__335(w__699 ,w__82);
  buf g__336(w__714 ,w__5);
  buf g__337(w__709 ,w__102);
  buf g__338(w__708 ,w__100);
  buf g__339(w__710 ,w__107);
  buf g__340(w__702 ,w__98);
  buf g__341(w__704 ,w__99);
  buf g__342(w__694 ,w__73);
  buf g__343(w__696 ,w__72);
  buf g__344(w__712 ,w__108);
  buf g__345(w__698 ,w__77);
  buf g__346(w__690 ,w__59);
  buf g__347(w__715 ,w__114);
  buf g__348(w__686 ,w__47);
  buf g__349(w__684 ,w__35);
  buf g__350(w__713 ,w__109);
  buf g__351(w__717 ,w__115);
  not g__352(w__7 ,w__78);
  xor g__353(w__6 ,w__112 ,in1[33]);
  xor g__354(w__5 ,w__104 ,in1[31]);
  xor g__355(w__4 ,w__78 ,in1[24]);
  xor g__356(w__3 ,w__65 ,in1[14]);
  xor g__357(w__2 ,w__48 ,in1[6]);
  xor g__358(w__1 ,w__31 ,in1[2]);
  or g__359(out4 ,w__131 ,w__301);
  nor g__360(w__301 ,w__193 ,w__300);
  or g__361(w__300 ,w__226 ,w__299);
  nor g__362(w__299 ,w__198 ,w__298);
  nor g__363(w__298 ,w__124 ,w__297);
  nor g__364(w__297 ,w__220 ,w__296);
  nor g__365(w__296 ,w__212 ,w__295);
  nor g__366(w__295 ,w__200 ,w__294);
  nor g__367(w__294 ,w__225 ,w__293);
  nor g__368(w__293 ,w__190 ,w__292);
  nor g__369(w__292 ,w__119 ,w__291);
  nor g__370(w__291 ,w__222 ,w__290);
  nor g__371(w__290 ,w__219 ,w__289);
  nor g__372(w__289 ,w__209 ,w__288);
  nor g__373(w__288 ,w__123 ,w__287);
  nor g__374(w__287 ,w__201 ,w__286);
  nor g__375(w__286 ,w__134 ,w__285);
  nor g__376(w__285 ,w__195 ,w__284);
  nor g__377(w__284 ,w__130 ,w__283);
  nor g__378(w__283 ,w__191 ,w__282);
  nor g__379(w__282 ,w__132 ,w__281);
  nor g__380(w__281 ,w__229 ,w__280);
  nor g__381(w__280 ,w__126 ,w__279);
  nor g__382(w__279 ,w__223 ,w__278);
  nor g__383(w__278 ,w__205 ,w__277);
  nor g__384(w__277 ,w__216 ,w__276);
  nor g__385(w__276 ,w__215 ,w__275);
  nor g__386(w__275 ,w__210 ,w__274);
  nor g__387(w__274 ,w__117 ,w__273);
  nor g__388(w__273 ,w__206 ,w__272);
  nor g__389(w__272 ,w__125 ,w__271);
  nor g__390(w__271 ,w__202 ,w__270);
  nor g__391(w__270 ,w__214 ,w__269);
  nor g__392(w__269 ,w__204 ,w__268);
  nor g__393(w__268 ,w__135 ,w__267);
  nor g__394(w__267 ,w__196 ,w__266);
  nor g__395(w__266 ,w__213 ,w__265);
  nor g__396(w__265 ,w__194 ,w__264);
  nor g__397(w__264 ,w__120 ,w__263);
  nor g__398(w__263 ,w__192 ,w__262);
  nor g__399(w__262 ,w__137 ,w__261);
  nor g__400(w__261 ,w__189 ,w__260);
  nor g__401(w__260 ,w__116 ,w__259);
  nor g__402(w__259 ,w__230 ,w__258);
  nor g__403(w__258 ,w__127 ,w__257);
  nor g__404(w__257 ,w__227 ,w__256);
  nor g__405(w__256 ,w__133 ,w__255);
  nor g__406(w__255 ,w__224 ,w__254);
  nor g__407(w__254 ,w__136 ,w__253);
  nor g__408(w__253 ,w__221 ,w__252);
  nor g__409(w__252 ,w__129 ,w__251);
  nor g__410(w__251 ,w__217 ,w__250);
  nor g__411(w__250 ,w__128 ,w__249);
  nor g__412(w__249 ,w__231 ,w__248);
  nor g__413(w__248 ,w__138 ,w__247);
  nor g__414(w__247 ,w__211 ,w__246);
  nor g__415(w__246 ,w__118 ,w__245);
  nor g__416(w__245 ,w__199 ,w__244);
  nor g__417(w__244 ,w__122 ,w__243);
  nor g__418(w__243 ,w__207 ,w__242);
  nor g__419(w__242 ,w__208 ,w__241);
  nor g__420(w__241 ,w__218 ,w__240);
  nor g__421(w__240 ,w__121 ,w__239);
  nor g__422(w__239 ,w__203 ,w__238);
  nor g__423(w__238 ,w__228 ,w__237);
  nor g__424(w__237 ,w__197 ,w__236);
  nor g__425(w__236 ,w__234 ,w__235);
  nor g__426(w__235 ,w__684 ,w__233);
  and g__427(w__234 ,in4[1] ,w__232);
  nor g__428(w__233 ,in4[1] ,w__232);
  nor g__429(w__231 ,w__523 ,in4[8]);
  nor g__430(w__230 ,w__527 ,in4[13]);
  nor g__431(w__229 ,w__529 ,in4[24]);
  nor g__432(w__228 ,w__185 ,w__486);
  nor g__433(w__227 ,w__525 ,in4[12]);
  nor g__434(w__226 ,w__183 ,w__490);
  nor g__435(w__225 ,w__178 ,w__480);
  nor g__436(w__224 ,w__519 ,in4[11]);
  nor g__437(w__223 ,w__521 ,in4[23]);
  nor g__438(w__222 ,w__543 ,in4[29]);
  nor g__439(w__221 ,w__517 ,in4[10]);
  nor g__440(w__220 ,w__501 ,in4[32]);
  nor g__441(w__219 ,w__179 ,w__492);
  nor g__442(w__218 ,w__483 ,in4[4]);
  nor g__443(w__217 ,w__515 ,in4[9]);
  nor g__444(w__216 ,w__481 ,in4[22]);
  nor g__445(w__215 ,w__181 ,w__496);
  nor g__446(w__214 ,w__186 ,w__498);
  nor g__447(w__213 ,w__182 ,w__488);
  nor g__448(w__212 ,w__180 ,w__494);
  nor g__449(w__211 ,w__505 ,in4[7]);
  or g__450(w__232 ,w__188 ,in4[0]);
  and g__451(w__210 ,w__496 ,w__181);
  and g__452(w__209 ,w__492 ,w__179);
  and g__453(w__208 ,in4[4] ,w__483);
  nor g__454(w__207 ,w__509 ,in4[5]);
  nor g__455(w__206 ,w__513 ,in4[20]);
  and g__456(w__205 ,in4[22] ,w__481);
  and g__457(w__204 ,w__498 ,w__186);
  nor g__458(w__203 ,w__507 ,in4[3]);
  nor g__459(w__202 ,w__537 ,in4[19]);
  nor g__460(w__201 ,w__541 ,in4[27]);
  and g__461(w__200 ,w__494 ,w__180);
  nor g__462(w__199 ,w__511 ,in4[6]);
  and g__463(w__198 ,w__490 ,w__183);
  and g__464(w__197 ,w__486 ,w__185);
  nor g__465(w__196 ,w__535 ,in4[17]);
  nor g__466(w__195 ,w__539 ,in4[26]);
  and g__467(w__194 ,w__488 ,w__182);
  nor g__468(w__193 ,w__499 ,in4[34]);
  nor g__469(w__192 ,w__503 ,in4[15]);
  nor g__470(w__191 ,w__533 ,in4[25]);
  and g__471(w__190 ,w__480 ,w__178);
  nor g__472(w__189 ,w__531 ,in4[14]);
  not g__473(w__188 ,w__683);
  not g__475(w__186 ,in4[18]);
  not g__476(w__185 ,in4[2]);
  not g__478(w__183 ,in4[33]);
  not g__479(w__182 ,in4[16]);
  not g__480(w__181 ,in4[21]);
  not g__481(w__180 ,in4[31]);
  not g__482(w__179 ,in4[28]);
  not g__483(w__178 ,in4[30]);
  and g__523(w__138 ,in4[7] ,w__505);
  and g__524(w__137 ,in4[14] ,w__531);
  and g__525(w__136 ,in4[10] ,w__517);
  and g__526(w__135 ,in4[17] ,w__535);
  and g__527(w__134 ,in4[26] ,w__539);
  and g__528(w__133 ,in4[11] ,w__519);
  and g__529(w__132 ,in4[24] ,w__529);
  and g__530(w__131 ,in4[34] ,w__499);
  and g__531(w__130 ,in4[25] ,w__533);
  and g__532(w__129 ,in4[9] ,w__515);
  and g__533(w__128 ,in4[8] ,w__523);
  and g__534(w__127 ,in4[12] ,w__525);
  and g__535(w__126 ,in4[23] ,w__521);
  and g__536(w__125 ,in4[19] ,w__537);
  and g__537(w__124 ,in4[32] ,w__501);
  and g__538(w__123 ,in4[27] ,w__541);
  and g__539(w__122 ,in4[5] ,w__509);
  and g__540(w__121 ,in4[3] ,w__507);
  and g__541(w__120 ,in4[15] ,w__503);
  and g__542(w__119 ,in4[29] ,w__543);
  and g__543(w__118 ,in4[6] ,w__511);
  and g__544(w__117 ,in4[20] ,w__513);
  and g__545(w__116 ,in4[13] ,w__527);
  or g__546(out1 ,w__316 ,w__476);
  nor g__547(w__476 ,w__366 ,w__475);
  nor g__548(w__475 ,w__399 ,w__474);
  nor g__549(w__474 ,w__372 ,w__473);
  nor g__550(w__473 ,w__393 ,w__472);
  nor g__551(w__472 ,w__306 ,w__471);
  nor g__552(w__471 ,w__385 ,w__470);
  nor g__553(w__470 ,w__375 ,w__469);
  nor g__554(w__469 ,w__398 ,w__468);
  nor g__555(w__468 ,w__363 ,w__467);
  nor g__556(w__467 ,w__404 ,w__466);
  nor g__557(w__466 ,w__310 ,w__465);
  nor g__558(w__465 ,w__392 ,w__464);
  nor g__559(w__464 ,w__383 ,w__463);
  nor g__560(w__463 ,w__380 ,w__462);
  nor g__561(w__462 ,w__308 ,w__461);
  nor g__562(w__461 ,w__374 ,w__460);
  nor g__563(w__460 ,w__315 ,w__459);
  nor g__564(w__459 ,w__370 ,w__458);
  nor g__565(w__458 ,w__307 ,w__457);
  nor g__566(w__457 ,w__397 ,w__456);
  nor g__567(w__456 ,w__305 ,w__455);
  nor g__568(w__455 ,w__402 ,w__454);
  nor g__569(w__454 ,w__317 ,w__453);
  nor g__570(w__453 ,w__379 ,w__452);
  nor g__571(w__452 ,w__390 ,w__451);
  nor g__572(w__451 ,w__389 ,w__450);
  nor g__573(w__450 ,w__384 ,w__449);
  nor g__574(w__449 ,w__368 ,w__448);
  nor g__575(w__448 ,w__312 ,w__447);
  nor g__576(w__447 ,w__378 ,w__446);
  nor g__577(w__446 ,w__321 ,w__445);
  nor g__578(w__445 ,w__388 ,w__444);
  nor g__579(w__444 ,w__376 ,w__443);
  nor g__580(w__443 ,w__373 ,w__442);
  nor g__581(w__442 ,w__314 ,w__441);
  nor g__582(w__441 ,w__386 ,w__440);
  nor g__583(w__440 ,w__369 ,w__439);
  nor g__584(w__439 ,w__367 ,w__438);
  nor g__585(w__438 ,w__313 ,w__437);
  nor g__586(w__437 ,w__365 ,w__436);
  nor g__587(w__436 ,w__311 ,w__435);
  nor g__588(w__435 ,w__405 ,w__434);
  nor g__589(w__434 ,w__302 ,w__433);
  nor g__590(w__433 ,w__403 ,w__432);
  nor g__591(w__432 ,w__323 ,w__431);
  nor g__592(w__431 ,w__400 ,w__430);
  nor g__593(w__430 ,w__303 ,w__429);
  nor g__594(w__429 ,w__396 ,w__428);
  nor g__595(w__428 ,w__318 ,w__427);
  nor g__596(w__427 ,w__394 ,w__426);
  nor g__597(w__426 ,w__304 ,w__425);
  nor g__598(w__425 ,w__395 ,w__424);
  nor g__599(w__424 ,w__309 ,w__423);
  nor g__600(w__423 ,w__387 ,w__422);
  nor g__601(w__422 ,w__324 ,w__421);
  nor g__602(w__421 ,w__364 ,w__420);
  nor g__603(w__420 ,w__320 ,w__419);
  nor g__604(w__419 ,w__381 ,w__418);
  nor g__605(w__418 ,w__322 ,w__417);
  nor g__606(w__417 ,w__382 ,w__416);
  nor g__607(w__416 ,w__391 ,w__415);
  nor g__608(w__415 ,w__377 ,w__414);
  nor g__609(w__414 ,w__319 ,w__413);
  nor g__610(w__413 ,w__401 ,w__412);
  nor g__611(w__412 ,w__371 ,w__411);
  nor g__612(w__411 ,w__409 ,w__410);
  and g__613(w__410 ,w__684 ,w__408);
  nor g__614(w__409 ,in2[1] ,w__407);
  or g__615(w__408 ,w__359 ,w__406);
  not g__616(w__407 ,w__406);
  nor g__617(w__405 ,w__329 ,in2[13]);
  nor g__618(w__404 ,w__332 ,in2[29]);
  nor g__619(w__403 ,w__340 ,in2[12]);
  nor g__620(w__402 ,w__339 ,in2[23]);
  nor g__621(w__401 ,w__358 ,in2[2]);
  nor g__622(w__400 ,w__345 ,in2[11]);
  nor g__623(w__399 ,w__356 ,in2[33]);
  nor g__624(w__398 ,w__351 ,in2[30]);
  nor g__625(w__397 ,w__344 ,in2[24]);
  nor g__626(w__396 ,w__348 ,in2[10]);
  nor g__627(w__395 ,w__341 ,in2[8]);
  nor g__628(w__394 ,w__342 ,in2[9]);
  nor g__629(w__393 ,w__337 ,in2[32]);
  nor g__630(w__392 ,w__352 ,in2[28]);
  nor g__631(w__391 ,w__361 ,w__328);
  nor g__632(w__390 ,w__357 ,w__326);
  nor g__633(w__389 ,w__354 ,in2[21]);
  nor g__634(w__388 ,w__360 ,in2[18]);
  nor g__635(w__387 ,w__350 ,in2[7]);
  nor g__636(w__386 ,w__355 ,in2[16]);
  nor g__637(w__385 ,w__353 ,in2[31]);
  or g__638(w__406 ,w__362 ,w__683);
  and g__639(w__384 ,in2[21] ,w__354);
  and g__640(w__383 ,in2[28] ,w__352);
  and g__641(w__382 ,w__328 ,w__361);
  nor g__642(w__381 ,w__335 ,in2[5]);
  nor g__643(w__380 ,w__336 ,in2[27]);
  and g__644(w__379 ,w__326 ,w__357);
  nor g__645(w__378 ,w__338 ,in2[19]);
  nor g__646(w__377 ,w__334 ,in2[3]);
  and g__647(w__376 ,in2[18] ,w__360);
  and g__648(w__375 ,in2[31] ,w__353);
  nor g__649(w__374 ,w__346 ,in2[26]);
  nor g__650(w__373 ,w__347 ,in2[17]);
  and g__651(w__372 ,in2[33] ,w__356);
  and g__652(w__371 ,in2[2] ,w__358);
  nor g__653(w__370 ,w__343 ,in2[25]);
  and g__654(w__369 ,in2[16] ,w__355);
  nor g__655(w__368 ,w__330 ,in2[20]);
  nor g__656(w__367 ,w__333 ,in2[15]);
  nor g__657(w__365 ,w__349 ,in2[14]);
  nor g__658(w__364 ,w__331 ,in2[6]);
  and g__659(w__363 ,in2[30] ,w__351);
  not g__660(w__362 ,in2[0]);
  not g__661(w__361 ,in2[4]);
  not g__662(w__360 ,w__701);
  not g__663(w__359 ,in2[1]);
  not g__664(w__358 ,w__685);
  not g__665(w__357 ,in2[22]);
  not g__666(w__356 ,w__716);
  not g__667(w__355 ,w__699);
  not g__668(w__354 ,w__704);
  not g__669(w__353 ,w__714);
  not g__670(w__352 ,w__711);
  not g__671(w__351 ,w__713);
  not g__672(w__335 ,w__688);
  not g__673(w__341 ,w__691);
  not g__674(w__342 ,w__692);
  not g__675(w__347 ,w__700);
  not g__676(w__338 ,w__702);
  not g__677(w__348 ,w__693);
  not g__678(w__330 ,w__703);
  not g__679(w__345 ,w__694);
  not g__680(w__339 ,w__706);
  not g__681(w__331 ,w__689);
  not g__682(w__340 ,w__695);
  not g__683(w__344 ,w__707);
  not g__684(w__343 ,w__708);
  not g__685(w__329 ,w__696);
  not g__686(w__346 ,w__709);
  not g__687(w__336 ,w__710);
  not g__688(w__349 ,w__697);
  not g__689(w__332 ,w__712);
  not g__690(w__337 ,w__715);
  not g__691(w__334 ,w__686);
  not g__692(w__350 ,w__690);
  not g__693(w__333 ,w__698);
  not g__694(w__328 ,w__327);
  not g__695(w__327 ,w__687);
  not g__696(w__326 ,w__325);
  not g__697(w__325 ,w__705);
  and g__698(w__324 ,in2[7] ,w__350);
  and g__699(w__323 ,in2[12] ,w__340);
  and g__700(w__322 ,in2[5] ,w__335);
  and g__701(w__321 ,in2[19] ,w__338);
  and g__702(w__320 ,in2[6] ,w__331);
  and g__703(w__319 ,in2[3] ,w__334);
  and g__704(w__318 ,in2[10] ,w__348);
  and g__705(w__317 ,in2[23] ,w__339);
  and g__706(w__315 ,in2[26] ,w__346);
  and g__707(w__314 ,in2[17] ,w__347);
  and g__708(w__313 ,in2[15] ,w__333);
  and g__709(w__312 ,in2[20] ,w__330);
  and g__710(w__311 ,in2[14] ,w__349);
  and g__711(w__310 ,in2[29] ,w__332);
  and g__712(w__309 ,in2[8] ,w__341);
  and g__713(w__308 ,in2[27] ,w__336);
  and g__714(w__307 ,in2[25] ,w__343);
  and g__715(w__306 ,in2[32] ,w__337);
  and g__716(w__305 ,in2[24] ,w__344);
  and g__717(w__304 ,in2[9] ,w__342);
  and g__718(w__303 ,in2[11] ,w__345);
  and g__719(w__302 ,in2[13] ,w__329);
  buf g__720(w__316 ,in2[34]);
  buf g__721(w__366 ,w__717);

endmodule

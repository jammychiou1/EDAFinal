module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, out1, out2, out3);

  input [12:0] in1;

  input [17:0] in2;

  input [31:0] in3, in7, in9;

  input in4, in5, in6, in8;

  input [4:0] in10;

  input [15:0] in11;

  output [32:0] out1;

  output [31:0] out2, out3;
  wire [12:0] in1;
  wire [17:0] in2;
  wire [31:0] in3, in7, in9;
  wire in4, in5, in6, in8;
  wire [4:0] in10;
  wire [15:0] in11;
  wire [32:0] out1;
  wire [31:0] out2, out3;
  wire add_25_22_n_23, add_25_22_n_24, add_25_22_n_25, add_25_22_n_26, add_25_22_n_27, add_25_22_n_28, add_25_22_n_29, add_25_22_n_30;
  wire add_25_22_n_31, add_25_22_n_32, add_25_22_n_33, add_25_22_n_34, add_25_22_n_35, add_25_22_n_36, out2[6], add_25_22_n_38;
  wire add_25_22_n_39, add_25_22_n_40, add_25_22_n_41, add_25_22_n_42, add_25_22_n_43, add_25_22_n_44, add_25_22_n_45, add_25_22_n_46;
  wire add_25_22_n_47, add_25_22_n_48, add_25_22_n_49, add_25_22_n_51, add_25_22_n_52, add_25_22_n_54, add_25_22_n_55, add_25_22_n_56;
  wire add_25_22_n_57, add_25_22_n_58, add_25_22_n_59, add_25_22_n_60, add_25_22_n_61, add_25_22_n_62, add_25_22_n_63, add_25_22_n_64;
  wire add_25_22_n_65, add_25_22_n_66, add_25_22_n_67, add_25_22_n_68, add_25_22_n_69, add_25_22_n_70, add_25_22_n_71, add_25_22_n_72;
  wire add_25_22_n_73, add_25_22_n_74, add_25_22_n_75, add_25_22_n_76, csa_tree_add_22_22_n_0, csa_tree_add_22_22_n_1, csa_tree_add_22_22_n_2, csa_tree_add_22_22_n_3;
  wire csa_tree_add_22_22_n_4, csa_tree_add_22_22_n_5, csa_tree_add_22_22_n_6, csa_tree_add_22_22_n_7, csa_tree_add_22_22_n_8, csa_tree_add_22_22_n_9, csa_tree_add_22_22_n_8, csa_tree_add_22_22_n_9;
  wire csa_tree_add_22_22_n_12, csa_tree_add_22_22_n_13, csa_tree_add_22_22_n_12, csa_tree_add_22_22_n_13, csa_tree_add_22_22_n_16, csa_tree_add_22_22_n_17, csa_tree_add_22_22_n_18, csa_tree_add_22_22_n_72;
  wire csa_tree_add_22_22_n_74, csa_tree_add_22_22_n_74, csa_tree_add_22_22_n_22, csa_tree_add_22_22_n_23, csa_tree_add_22_22_n_22, csa_tree_add_22_22_n_23, csa_tree_add_22_22_n_26, csa_tree_add_22_22_n_27;
  wire csa_tree_add_22_22_n_28, csa_tree_add_22_22_n_69, csa_tree_add_22_22_n_71, csa_tree_add_22_22_n_71, csa_tree_add_22_22_n_32, csa_tree_add_22_22_n_33, csa_tree_add_22_22_n_34, csa_tree_add_22_22_n_35;
  wire csa_tree_add_22_22_n_36, csa_tree_add_22_22_n_75, csa_tree_add_22_22_n_77, csa_tree_add_22_22_n_77, csa_tree_add_22_22_n_78, csa_tree_add_22_22_n_80, csa_tree_add_22_22_n_80, csa_tree_add_22_22_n_43;
  wire csa_tree_add_22_22_n_45, csa_tree_add_22_22_n_45, csa_tree_add_22_22_n_46, csa_tree_add_22_22_n_48, csa_tree_add_22_22_n_48, csa_tree_add_22_22_n_49, csa_tree_add_22_22_n_51, csa_tree_add_22_22_n_51;
  wire csa_tree_add_22_22_n_52, csa_tree_add_22_22_n_54, csa_tree_add_22_22_n_54, csa_tree_add_22_22_n_55, csa_tree_add_22_22_n_57, csa_tree_add_22_22_n_57, csa_tree_add_22_22_n_58, csa_tree_add_22_22_n_60;
  wire csa_tree_add_22_22_n_60, csa_tree_add_22_22_n_61, csa_tree_add_22_22_n_63, csa_tree_add_22_22_n_63, csa_tree_add_22_22_n_67, csa_tree_add_22_22_n_68, csa_tree_add_22_22_n_68, csa_tree_add_22_22_n_67;
  wire csa_tree_add_22_22_n_68, csa_tree_add_22_22_n_69, csa_tree_add_22_22_n_71, csa_tree_add_22_22_n_71, csa_tree_add_22_22_n_72, csa_tree_add_22_22_n_74, csa_tree_add_22_22_n_74, csa_tree_add_22_22_n_75;
  wire csa_tree_add_22_22_n_77, csa_tree_add_22_22_n_77, csa_tree_add_22_22_n_78, csa_tree_add_22_22_n_80, csa_tree_add_22_22_n_80, csa_tree_add_22_22_n_81, csa_tree_add_22_22_n_82, csa_tree_add_22_22_n_83;
  wire csa_tree_add_22_22_n_84, csa_tree_add_22_22_n_85, csa_tree_add_22_22_n_86, csa_tree_add_22_22_n_87, csa_tree_add_22_22_n_88, csa_tree_add_22_22_n_89, csa_tree_add_22_22_n_90, csa_tree_add_22_22_n_91;
  wire csa_tree_add_22_22_n_92, csa_tree_add_22_22_n_94, csa_tree_add_22_22_n_95, csa_tree_add_22_22_n_96, csa_tree_add_22_22_n_97, csa_tree_add_22_22_n_98, csa_tree_add_22_22_n_99, csa_tree_add_22_22_n_100;
  wire csa_tree_add_22_22_n_101, csa_tree_add_22_22_n_102, csa_tree_add_22_22_n_103, csa_tree_add_22_22_n_104, csa_tree_add_22_22_n_105, csa_tree_add_22_22_n_106, csa_tree_add_22_22_n_107, csa_tree_add_22_22_n_108;
  wire csa_tree_add_22_22_n_109, csa_tree_add_22_22_n_110, csa_tree_add_22_22_n_111, csa_tree_add_22_22_n_112, csa_tree_add_22_22_n_113, csa_tree_add_22_22_n_114, csa_tree_add_22_22_n_115, csa_tree_add_22_22_n_116;
  wire csa_tree_add_22_22_n_117, csa_tree_add_22_22_n_118, csa_tree_add_22_22_n_119, csa_tree_add_22_22_n_120, csa_tree_add_22_22_n_121, csa_tree_add_22_22_n_122, csa_tree_add_22_22_n_123, csa_tree_add_22_22_n_124;
  wire csa_tree_add_22_22_n_125, csa_tree_add_22_22_n_126, csa_tree_add_22_22_n_127, csa_tree_add_22_22_n_128, csa_tree_add_22_22_n_129, csa_tree_add_22_22_n_130, csa_tree_add_22_22_n_131, csa_tree_add_22_22_n_132;
  wire csa_tree_add_22_22_n_133, csa_tree_add_22_22_n_134, csa_tree_add_22_22_n_135, csa_tree_add_22_22_n_136, csa_tree_add_22_22_n_137, csa_tree_add_22_22_n_138, csa_tree_add_22_22_n_139, csa_tree_add_22_22_n_140;
  wire csa_tree_add_22_22_n_141, csa_tree_add_22_22_n_142, csa_tree_add_22_22_n_143, csa_tree_add_22_22_n_144, csa_tree_add_22_22_n_145, csa_tree_add_22_22_n_146, csa_tree_add_22_22_n_147, csa_tree_add_22_22_n_148;
  wire csa_tree_add_22_22_n_149, csa_tree_add_22_22_n_150, csa_tree_add_22_22_n_151, csa_tree_add_22_22_n_152, csa_tree_add_22_22_n_153, csa_tree_add_22_22_n_154, csa_tree_add_22_22_n_155, csa_tree_add_22_22_n_156;
  wire csa_tree_add_22_22_n_157, csa_tree_add_22_22_n_158, csa_tree_add_22_22_n_159, csa_tree_add_22_22_n_160, csa_tree_add_22_22_n_161, csa_tree_add_22_22_n_162, csa_tree_add_22_22_n_163, csa_tree_add_22_22_n_164;
  wire csa_tree_add_22_22_n_165, csa_tree_add_22_22_n_166, csa_tree_add_22_22_n_167, csa_tree_add_22_22_n_170, csa_tree_add_22_22_n_171, csa_tree_add_22_22_n_172, csa_tree_add_22_22_n_173, csa_tree_add_22_22_n_174;
  wire csa_tree_add_22_22_n_175, csa_tree_add_22_22_n_176, csa_tree_add_22_22_n_177, csa_tree_add_22_22_n_178, csa_tree_add_22_22_n_179, csa_tree_add_22_22_n_180, csa_tree_add_22_22_n_181, csa_tree_add_22_22_n_182;
  wire csa_tree_add_22_22_n_183, csa_tree_add_22_22_n_184, csa_tree_add_22_22_n_185, csa_tree_add_22_22_n_186, csa_tree_add_22_22_n_187, csa_tree_add_22_22_n_188, csa_tree_add_22_22_n_189, csa_tree_add_22_22_n_190;
  wire csa_tree_add_22_22_n_191, csa_tree_add_22_22_n_192, csa_tree_add_22_22_n_193, csa_tree_add_22_22_n_194, csa_tree_add_22_22_n_195, csa_tree_add_22_22_n_196, csa_tree_add_22_22_n_197, csa_tree_add_22_22_n_198;
  wire csa_tree_add_22_22_n_199, csa_tree_add_22_22_n_200, csa_tree_add_22_22_n_201, csa_tree_add_22_22_n_202, csa_tree_add_22_22_n_203, csa_tree_add_22_22_n_204, csa_tree_add_22_22_n_205, csa_tree_add_22_22_n_206;
  wire csa_tree_add_22_22_n_207, csa_tree_add_22_22_n_208, csa_tree_add_22_22_n_209, csa_tree_add_22_22_n_210, csa_tree_add_22_22_n_211, csa_tree_add_22_22_n_212, csa_tree_add_22_22_n_213, csa_tree_add_22_22_n_214;
  wire csa_tree_add_22_22_n_215, csa_tree_add_22_22_n_216, csa_tree_add_22_22_n_217, csa_tree_add_22_22_n_218, csa_tree_add_22_22_n_219, csa_tree_add_22_22_n_220, csa_tree_add_22_22_n_221, csa_tree_add_22_22_n_222;
  wire csa_tree_add_22_22_n_223, csa_tree_add_22_22_n_224, csa_tree_add_22_22_n_225, csa_tree_add_22_22_n_226, csa_tree_add_22_22_n_227, csa_tree_add_22_22_n_228, csa_tree_add_22_22_n_229, csa_tree_add_22_22_n_230;
  wire csa_tree_add_22_22_n_232, csa_tree_add_22_22_n_233, csa_tree_add_22_22_n_234, csa_tree_add_22_22_n_235, csa_tree_add_22_22_n_236, csa_tree_add_22_22_n_237, csa_tree_add_22_22_n_238, csa_tree_add_22_22_n_239;
  wire csa_tree_add_22_22_n_240, csa_tree_add_22_22_n_241, csa_tree_add_22_22_n_242, csa_tree_add_22_22_n_243, csa_tree_add_22_22_n_244, csa_tree_add_22_22_n_245, csa_tree_add_22_22_n_246, csa_tree_add_22_22_n_247;
  wire csa_tree_add_22_22_n_248, csa_tree_add_22_22_n_249, csa_tree_add_22_22_n_250, csa_tree_add_22_22_n_251, csa_tree_add_22_22_n_252, csa_tree_add_22_22_n_253, csa_tree_add_22_22_n_254, csa_tree_add_22_22_n_255;
  wire csa_tree_add_22_22_n_256, csa_tree_add_22_22_n_257, csa_tree_add_22_22_n_258, csa_tree_add_22_22_n_259, csa_tree_add_22_22_n_260, csa_tree_add_22_22_n_261, csa_tree_add_22_22_n_262, csa_tree_add_22_22_n_263;
  wire csa_tree_add_22_22_n_264, csa_tree_add_22_22_n_265, csa_tree_add_22_22_n_266, csa_tree_add_22_22_n_267, csa_tree_add_22_22_n_268, csa_tree_add_22_22_n_269, csa_tree_add_22_22_n_270, csa_tree_add_22_22_n_271;
  wire csa_tree_add_22_22_n_272, csa_tree_add_22_22_n_273, csa_tree_add_22_22_n_274, csa_tree_add_22_22_n_275, csa_tree_add_22_22_n_276, csa_tree_add_22_22_n_277, csa_tree_add_22_22_n_278, csa_tree_add_22_22_n_279;
  wire csa_tree_add_22_22_n_280, csa_tree_add_22_22_n_281, csa_tree_add_22_22_n_282, csa_tree_add_22_22_n_283, csa_tree_add_22_22_n_284, csa_tree_add_22_22_n_285, csa_tree_add_22_22_n_287, csa_tree_add_22_22_n_288;
  wire csa_tree_add_22_22_n_289, csa_tree_add_22_22_n_290, csa_tree_add_22_22_n_291, csa_tree_add_22_22_n_292, csa_tree_add_22_22_n_293, csa_tree_add_22_22_n_294, csa_tree_add_22_22_n_295, csa_tree_add_22_22_n_296;
  wire csa_tree_add_22_22_n_297, csa_tree_add_22_22_n_298, csa_tree_add_22_22_n_299, csa_tree_add_22_22_n_300, csa_tree_add_22_22_n_301, csa_tree_add_22_22_n_302, csa_tree_add_22_22_n_303, csa_tree_add_22_22_n_304;
  wire csa_tree_add_22_22_n_305, csa_tree_add_22_22_n_306, csa_tree_add_22_22_n_307, csa_tree_add_22_22_n_308, csa_tree_add_22_22_n_309, csa_tree_add_22_22_n_310, csa_tree_add_22_22_n_311, csa_tree_add_22_22_n_312;
  wire csa_tree_add_22_22_n_313, csa_tree_add_22_22_n_314, csa_tree_add_22_22_n_315, csa_tree_add_22_22_n_316, csa_tree_add_22_22_n_317, csa_tree_add_22_22_n_318, csa_tree_add_22_22_n_319, csa_tree_add_22_22_n_320;
  wire csa_tree_add_22_22_n_321, csa_tree_add_22_22_n_322, csa_tree_add_22_22_n_323, csa_tree_add_22_22_n_324, csa_tree_add_22_22_n_325, csa_tree_add_22_22_n_326, csa_tree_add_22_22_n_327, csa_tree_add_22_22_n_328;
  wire csa_tree_add_22_22_n_329, csa_tree_add_22_22_n_330, csa_tree_add_22_22_n_331, csa_tree_add_22_22_n_332, csa_tree_add_22_22_n_333, csa_tree_add_22_22_n_334, csa_tree_add_22_22_n_335, csa_tree_add_22_22_n_336;
  wire csa_tree_add_22_22_n_337, csa_tree_add_22_22_n_338, csa_tree_add_22_22_n_339, csa_tree_add_22_22_n_340, csa_tree_add_22_22_n_341, csa_tree_add_22_22_n_342, csa_tree_add_22_22_n_343, csa_tree_add_22_22_n_344;
  wire csa_tree_add_22_22_n_345, csa_tree_add_22_22_n_346, csa_tree_add_22_22_n_347, csa_tree_add_22_22_n_348, csa_tree_add_22_22_n_349, csa_tree_add_22_22_n_350, csa_tree_add_22_22_n_351, csa_tree_add_22_22_n_352;
  wire csa_tree_add_22_22_n_353, csa_tree_add_22_22_n_354, csa_tree_add_22_22_n_355, csa_tree_add_22_22_n_356, csa_tree_add_22_22_n_357, csa_tree_add_22_22_n_358, csa_tree_add_22_22_n_359, csa_tree_add_22_22_n_360;
  wire csa_tree_add_22_22_n_361, csa_tree_add_22_22_n_362, csa_tree_add_22_22_n_363, csa_tree_add_22_22_n_364, csa_tree_add_22_22_n_365, csa_tree_add_22_22_n_366, csa_tree_add_22_22_n_367, csa_tree_add_22_22_n_368;
  wire csa_tree_add_22_22_n_369, csa_tree_add_22_22_n_370, csa_tree_add_22_22_n_371, csa_tree_add_22_22_n_373, csa_tree_add_22_22_n_375, csa_tree_add_22_22_n_376, csa_tree_add_22_22_n_377, csa_tree_add_22_22_n_378;
  wire csa_tree_add_22_22_n_379, csa_tree_add_22_22_n_380, csa_tree_add_22_22_n_381, csa_tree_add_22_22_n_382, csa_tree_add_22_22_n_383, csa_tree_add_22_22_n_384, csa_tree_add_22_22_n_385, csa_tree_add_22_22_n_386;
  wire csa_tree_add_22_22_n_387, csa_tree_add_22_22_n_388, csa_tree_add_22_22_n_389, csa_tree_add_22_22_n_390, csa_tree_add_22_22_n_391, csa_tree_add_22_22_n_392, csa_tree_add_22_22_n_393, csa_tree_add_22_22_n_394;
  wire csa_tree_add_22_22_n_395, csa_tree_add_22_22_n_396, csa_tree_add_22_22_n_397, csa_tree_add_22_22_n_398, csa_tree_add_22_22_n_399, csa_tree_add_22_22_n_400, csa_tree_add_22_22_n_401, csa_tree_add_22_22_n_402;
  wire csa_tree_add_22_22_n_403, csa_tree_add_22_22_n_405, csa_tree_add_22_22_n_407, csa_tree_add_22_22_n_408, csa_tree_add_22_22_n_409, csa_tree_add_22_22_n_410, csa_tree_add_22_22_n_411, csa_tree_add_22_22_n_412;
  wire csa_tree_add_22_22_n_413, csa_tree_add_22_22_n_414, csa_tree_add_22_22_n_415, csa_tree_add_22_22_n_416, csa_tree_add_22_22_n_417, csa_tree_add_22_22_n_418, csa_tree_add_22_22_n_419, csa_tree_add_22_22_n_420;
  wire csa_tree_add_22_22_n_421, csa_tree_add_22_22_n_422, csa_tree_add_22_22_n_423, csa_tree_add_22_22_n_424, csa_tree_add_22_22_n_425, csa_tree_add_22_22_n_426, csa_tree_add_22_22_n_427, csa_tree_add_22_22_n_428;
  wire csa_tree_add_22_22_n_429, csa_tree_add_22_22_n_430, csa_tree_add_22_22_n_431, csa_tree_add_22_22_n_432, csa_tree_add_22_22_n_434, csa_tree_add_22_22_n_435, csa_tree_add_22_22_n_436, csa_tree_add_22_22_n_438;
  wire csa_tree_add_22_22_n_439, csa_tree_add_22_22_n_440, csa_tree_add_22_22_n_441, csa_tree_add_22_22_n_442, csa_tree_add_22_22_n_443, csa_tree_add_22_22_n_444, csa_tree_add_22_22_n_445, csa_tree_add_22_22_n_446;
  wire csa_tree_add_22_22_n_447, csa_tree_add_22_22_n_448, csa_tree_add_22_22_n_449, csa_tree_add_22_22_n_450, csa_tree_add_22_22_n_451, csa_tree_add_22_22_n_452, csa_tree_add_22_22_n_453, csa_tree_add_22_22_n_454;
  wire csa_tree_add_22_22_n_455, csa_tree_add_22_22_n_456, csa_tree_add_22_22_n_457, csa_tree_add_22_22_n_458, csa_tree_add_22_22_n_459, csa_tree_add_22_22_n_460, csa_tree_add_22_22_n_461, csa_tree_add_22_22_n_462;
  wire csa_tree_add_22_22_n_463, csa_tree_add_22_22_n_464, csa_tree_add_22_22_n_466, csa_tree_add_22_22_n_467, csa_tree_add_22_22_n_468, csa_tree_add_22_22_n_469, csa_tree_add_22_22_n_473, csa_tree_add_22_22_n_474;
  wire csa_tree_add_22_22_n_475, csa_tree_add_22_22_n_476, csa_tree_add_22_22_n_477, csa_tree_add_22_22_n_478, csa_tree_add_22_22_n_479, csa_tree_add_22_22_n_480, csa_tree_add_22_22_n_481, csa_tree_add_22_22_n_482;
  wire csa_tree_add_22_22_n_483, csa_tree_add_22_22_n_484, csa_tree_add_22_22_n_485, csa_tree_add_22_22_n_486, csa_tree_add_22_22_n_487, csa_tree_add_22_22_n_488, csa_tree_add_22_22_n_489, csa_tree_add_22_22_n_490;
  wire csa_tree_add_22_22_n_491, csa_tree_add_22_22_n_492, csa_tree_add_22_22_n_493, csa_tree_add_22_22_n_494, csa_tree_add_22_22_n_495, csa_tree_add_22_22_n_496, csa_tree_add_22_22_n_497, csa_tree_add_22_22_n_498;
  wire csa_tree_add_22_22_n_501, csa_tree_add_22_22_n_503, csa_tree_add_22_22_n_504, csa_tree_add_22_22_n_505, csa_tree_add_22_22_n_506, csa_tree_add_22_22_n_507, csa_tree_add_22_22_n_508, csa_tree_add_22_22_n_510;
  wire csa_tree_add_24_21_groupi_n_0, csa_tree_add_24_21_groupi_n_1, csa_tree_add_24_21_groupi_n_2, csa_tree_add_24_21_groupi_n_3, csa_tree_add_24_21_groupi_n_58, csa_tree_add_24_21_groupi_n_60, csa_tree_add_24_21_groupi_n_61, csa_tree_add_24_21_groupi_n_63;
  wire csa_tree_add_24_21_groupi_n_52, csa_tree_add_24_21_groupi_n_54, csa_tree_add_24_21_groupi_n_64, csa_tree_add_24_21_groupi_n_66, csa_tree_add_24_21_groupi_n_66, csa_tree_add_24_21_groupi_n_61, csa_tree_add_24_21_groupi_n_63, csa_tree_add_24_21_groupi_n_63;
  wire csa_tree_add_24_21_groupi_n_70, csa_tree_add_24_21_groupi_n_72, csa_tree_add_24_21_groupi_n_72, csa_tree_add_24_21_groupi_n_70, csa_tree_add_24_21_groupi_n_72, csa_tree_add_24_21_groupi_n_58, csa_tree_add_24_21_groupi_n_60, csa_tree_add_24_21_groupi_n_60;
  wire csa_tree_add_24_21_groupi_n_67, csa_tree_add_24_21_groupi_n_69, csa_tree_add_24_21_groupi_n_69, csa_tree_add_24_21_groupi_n_55, csa_tree_add_24_21_groupi_n_57, csa_tree_add_24_21_groupi_n_29, csa_tree_add_24_21_groupi_n_30, csa_tree_add_24_21_groupi_n_64;
  wire csa_tree_add_24_21_groupi_n_66, csa_tree_add_24_21_groupi_n_33, csa_tree_add_24_21_groupi_n_34, csa_tree_add_24_21_groupi_n_55, csa_tree_add_24_21_groupi_n_57, csa_tree_add_24_21_groupi_n_57, csa_tree_add_24_21_groupi_n_38, csa_tree_add_24_21_groupi_n_39;
  wire csa_tree_add_24_21_groupi_n_40, csa_tree_add_24_21_groupi_n_41, csa_tree_add_24_21_groupi_n_42, csa_tree_add_24_21_groupi_n_43, csa_tree_add_24_21_groupi_n_67, csa_tree_add_24_21_groupi_n_69, csa_tree_add_22_22_n_85, csa_tree_add_22_22_n_86;
  wire csa_tree_add_22_22_n_86, csa_tree_add_24_21_groupi_n_52, csa_tree_add_24_21_groupi_n_54, csa_tree_add_24_21_groupi_n_54, csa_tree_add_24_21_groupi_n_52, csa_tree_add_24_21_groupi_n_54, csa_tree_add_24_21_groupi_n_54, csa_tree_add_24_21_groupi_n_55;
  wire csa_tree_add_24_21_groupi_n_57, csa_tree_add_24_21_groupi_n_57, csa_tree_add_24_21_groupi_n_58, csa_tree_add_24_21_groupi_n_60, csa_tree_add_24_21_groupi_n_60, csa_tree_add_24_21_groupi_n_61, csa_tree_add_24_21_groupi_n_63, csa_tree_add_24_21_groupi_n_63;
  wire csa_tree_add_24_21_groupi_n_64, csa_tree_add_24_21_groupi_n_66, csa_tree_add_24_21_groupi_n_66, csa_tree_add_24_21_groupi_n_67, csa_tree_add_24_21_groupi_n_69, csa_tree_add_24_21_groupi_n_69, csa_tree_add_24_21_groupi_n_70, csa_tree_add_24_21_groupi_n_72;
  wire csa_tree_add_24_21_groupi_n_72, csa_tree_add_24_21_groupi_n_73, csa_tree_add_24_21_groupi_n_74, csa_tree_add_24_21_groupi_n_75, csa_tree_add_24_21_groupi_n_76, csa_tree_add_24_21_groupi_n_77, csa_tree_add_24_21_groupi_n_78, csa_tree_add_24_21_groupi_n_79;
  wire csa_tree_add_24_21_groupi_n_80, csa_tree_add_24_21_groupi_n_81, csa_tree_add_24_21_groupi_n_55, csa_tree_add_24_21_groupi_n_57, csa_tree_add_24_21_groupi_n_84, csa_tree_add_24_21_groupi_n_85, csa_tree_add_24_21_groupi_n_86, csa_tree_add_24_21_groupi_n_203;
  wire csa_tree_add_24_21_groupi_n_205, csa_tree_add_24_21_groupi_n_205, csa_tree_add_24_21_groupi_n_90, csa_tree_add_24_21_groupi_n_91, csa_tree_add_24_21_groupi_n_92, csa_tree_add_24_21_groupi_n_218, csa_tree_add_24_21_groupi_n_220, csa_tree_add_24_21_groupi_n_220;
  wire csa_tree_add_24_21_groupi_n_67, csa_tree_add_24_21_groupi_n_69, csa_tree_add_24_21_groupi_n_58, csa_tree_add_24_21_groupi_n_60, csa_tree_add_24_21_groupi_n_206, csa_tree_add_24_21_groupi_n_208, csa_tree_add_24_21_groupi_n_208, csa_tree_add_24_21_groupi_n_70;
  wire csa_tree_add_24_21_groupi_n_72, csa_tree_add_24_21_groupi_n_61, csa_tree_add_24_21_groupi_n_63, csa_tree_add_24_21_groupi_n_64, csa_tree_add_24_21_groupi_n_66, csa_tree_add_22_22_n_85, csa_tree_add_22_22_n_86, csa_tree_add_22_22_n_86;
  wire csa_tree_add_24_21_groupi_n_215, csa_tree_add_24_21_groupi_n_217, csa_tree_add_24_21_groupi_n_217, csa_tree_add_24_21_groupi_n_209, csa_tree_add_24_21_groupi_n_211, csa_tree_add_24_21_groupi_n_211, csa_tree_add_24_21_groupi_n_118, csa_tree_add_24_21_groupi_n_119;
  wire csa_tree_add_24_21_groupi_n_120, csa_tree_add_24_21_groupi_n_212, csa_tree_add_24_21_groupi_n_214, csa_tree_add_24_21_groupi_n_214, csa_tree_add_24_21_groupi_n_172, csa_tree_add_24_21_groupi_n_173, csa_tree_add_24_21_groupi_n_173, csa_tree_add_24_21_groupi_n_146;
  wire csa_tree_add_24_21_groupi_n_148, csa_tree_add_24_21_groupi_n_164, csa_tree_add_24_21_groupi_n_166, csa_tree_add_24_21_groupi_n_158, csa_tree_add_24_21_groupi_n_160, csa_tree_add_24_21_groupi_n_149, csa_tree_add_24_21_groupi_n_151, csa_tree_add_24_21_groupi_n_152;
  wire csa_tree_add_24_21_groupi_n_154, csa_tree_add_24_21_groupi_n_152, csa_tree_add_24_21_groupi_n_154, csa_tree_add_24_21_groupi_n_154, csa_tree_add_24_21_groupi_n_149, csa_tree_add_24_21_groupi_n_151, csa_tree_add_24_21_groupi_n_151, csa_tree_add_24_21_groupi_n_146;
  wire csa_tree_add_24_21_groupi_n_148, csa_tree_add_24_21_groupi_n_148, csa_tree_add_24_21_groupi_n_146, csa_tree_add_24_21_groupi_n_148, csa_tree_add_24_21_groupi_n_148, csa_tree_add_24_21_groupi_n_149, csa_tree_add_24_21_groupi_n_151, csa_tree_add_24_21_groupi_n_151;
  wire csa_tree_add_24_21_groupi_n_152, csa_tree_add_24_21_groupi_n_154, csa_tree_add_24_21_groupi_n_154, csa_tree_add_24_21_groupi_n_158, csa_tree_add_24_21_groupi_n_160, csa_tree_add_24_21_groupi_n_160, csa_tree_add_24_21_groupi_n_158, csa_tree_add_24_21_groupi_n_160;
  wire csa_tree_add_24_21_groupi_n_160, csa_tree_add_24_21_groupi_n_164, csa_tree_add_24_21_groupi_n_166, csa_tree_add_24_21_groupi_n_166, csa_tree_add_24_21_groupi_n_164, csa_tree_add_24_21_groupi_n_166, csa_tree_add_24_21_groupi_n_166, csa_tree_add_24_21_groupi_n_270;
  wire csa_tree_add_24_21_groupi_n_261, csa_tree_add_24_21_groupi_n_264, csa_tree_add_24_21_groupi_n_267, csa_tree_add_24_21_groupi_n_258, csa_tree_add_24_21_groupi_n_172, csa_tree_add_24_21_groupi_n_173, csa_tree_add_24_21_groupi_n_258, csa_tree_add_24_21_groupi_n_261;
  wire csa_tree_add_24_21_groupi_n_264, csa_tree_add_24_21_groupi_n_267, csa_tree_add_24_21_groupi_n_270, csa_tree_add_24_21_groupi_n_200, csa_tree_add_24_21_groupi_n_146, csa_tree_add_24_21_groupi_n_148, csa_tree_add_24_21_groupi_n_148, csa_tree_add_24_21_groupi_n_149;
  wire csa_tree_add_24_21_groupi_n_151, csa_tree_add_24_21_groupi_n_151, csa_tree_add_24_21_groupi_n_164, csa_tree_add_24_21_groupi_n_166, csa_tree_add_24_21_groupi_n_166, csa_tree_add_24_21_groupi_n_152, csa_tree_add_24_21_groupi_n_154, csa_tree_add_24_21_groupi_n_154;
  wire csa_tree_add_24_21_groupi_n_158, csa_tree_add_24_21_groupi_n_160, csa_tree_add_24_21_groupi_n_160, csa_tree_add_24_21_groupi_n_593, csa_tree_add_24_21_groupi_n_279, csa_tree_add_24_21_groupi_n_279, csa_tree_add_24_21_groupi_n_198, csa_tree_add_24_21_groupi_n_200;
  wire csa_tree_add_24_21_groupi_n_200, csa_tree_add_22_22_n_85, csa_tree_add_22_22_n_86, csa_tree_add_24_21_groupi_n_203, csa_tree_add_24_21_groupi_n_205, csa_tree_add_24_21_groupi_n_205, csa_tree_add_24_21_groupi_n_206, csa_tree_add_24_21_groupi_n_208;
  wire csa_tree_add_24_21_groupi_n_208, csa_tree_add_24_21_groupi_n_209, csa_tree_add_24_21_groupi_n_211, csa_tree_add_24_21_groupi_n_211, csa_tree_add_24_21_groupi_n_212, csa_tree_add_24_21_groupi_n_214, csa_tree_add_24_21_groupi_n_214, csa_tree_add_24_21_groupi_n_215;
  wire csa_tree_add_24_21_groupi_n_217, csa_tree_add_24_21_groupi_n_217, csa_tree_add_24_21_groupi_n_218, csa_tree_add_24_21_groupi_n_220, csa_tree_add_24_21_groupi_n_220, csa_tree_add_24_21_groupi_n_253, csa_tree_add_24_21_groupi_n_254, csa_tree_add_22_22_n_81;
  wire csa_tree_add_22_22_n_82, csa_tree_add_24_21_groupi_n_257, csa_tree_add_24_21_groupi_n_258, csa_tree_add_24_21_groupi_n_260, csa_tree_add_24_21_groupi_n_260, csa_tree_add_24_21_groupi_n_261, csa_tree_add_24_21_groupi_n_263, csa_tree_add_24_21_groupi_n_263;
  wire csa_tree_add_24_21_groupi_n_264, csa_tree_add_24_21_groupi_n_266, csa_tree_add_24_21_groupi_n_266, csa_tree_add_24_21_groupi_n_267, csa_tree_add_24_21_groupi_n_269, csa_tree_add_24_21_groupi_n_269, csa_tree_add_24_21_groupi_n_270, csa_tree_add_24_21_groupi_n_272;
  wire csa_tree_add_24_21_groupi_n_272, csa_tree_add_24_21_groupi_n_279, csa_tree_add_24_21_groupi_n_281, csa_tree_add_24_21_groupi_n_281, csa_tree_add_24_21_groupi_n_276, csa_tree_add_24_21_groupi_n_277, csa_tree_add_24_21_groupi_n_278, csa_tree_add_24_21_groupi_n_279;
  wire csa_tree_add_24_21_groupi_n_281, csa_tree_add_24_21_groupi_n_281, csa_tree_add_24_21_groupi_n_200, csa_tree_add_24_21_groupi_n_404, csa_tree_add_24_21_groupi_n_404, csa_tree_add_24_21_groupi_n_291, csa_tree_add_24_21_groupi_n_293, csa_tree_add_24_21_groupi_n_293;
  wire csa_tree_add_24_21_groupi_n_291, csa_tree_add_24_21_groupi_n_293, csa_tree_add_24_21_groupi_n_293, csa_tree_add_24_21_groupi_n_291, csa_tree_add_24_21_groupi_n_293, csa_tree_add_24_21_groupi_n_293, csa_tree_add_24_21_groupi_n_258, csa_tree_add_24_21_groupi_n_260;
  wire csa_tree_add_24_21_groupi_n_260, csa_tree_add_24_21_groupi_n_261, csa_tree_add_24_21_groupi_n_263, csa_tree_add_24_21_groupi_n_263, csa_tree_add_24_21_groupi_n_270, csa_tree_add_24_21_groupi_n_272, csa_tree_add_24_21_groupi_n_272, csa_tree_add_24_21_groupi_n_264;
  wire csa_tree_add_24_21_groupi_n_266, csa_tree_add_24_21_groupi_n_266, csa_tree_add_24_21_groupi_n_267, csa_tree_add_24_21_groupi_n_269, csa_tree_add_24_21_groupi_n_269, csa_tree_add_24_21_groupi_n_309, csa_tree_add_24_21_groupi_n_309, csa_tree_add_24_21_groupi_n_311;
  wire csa_tree_add_24_21_groupi_n_311, csa_tree_add_24_21_groupi_n_198, csa_tree_add_24_21_groupi_n_314, csa_tree_add_24_21_groupi_n_314, csa_tree_add_24_21_groupi_n_316, csa_tree_add_24_21_groupi_n_316, csa_tree_add_24_21_groupi_n_318, csa_tree_add_24_21_groupi_n_318;
  wire csa_tree_add_24_21_groupi_n_320, csa_tree_add_24_21_groupi_n_321, csa_tree_add_22_22_n_103, csa_tree_add_22_22_n_102, csa_tree_add_22_22_n_118, csa_tree_add_24_21_groupi_n_325, csa_tree_add_22_22_n_99, csa_tree_add_24_21_groupi_n_327;
  wire csa_tree_add_24_21_groupi_n_328, csa_tree_add_24_21_groupi_n_329, csa_tree_add_24_21_groupi_n_330, csa_tree_add_24_21_groupi_n_331, csa_tree_add_24_21_groupi_n_332, csa_tree_add_24_21_groupi_n_333, csa_tree_add_24_21_groupi_n_334, csa_tree_add_24_21_groupi_n_335;
  wire csa_tree_add_24_21_groupi_n_336, csa_tree_add_24_21_groupi_n_337, csa_tree_add_24_21_groupi_n_338, csa_tree_add_22_22_n_117, csa_tree_add_24_21_groupi_n_340, csa_tree_add_24_21_groupi_n_341, csa_tree_add_24_21_groupi_n_342, csa_tree_add_22_22_n_114;
  wire csa_tree_add_22_22_n_100, csa_tree_add_22_22_n_101, csa_tree_add_24_21_groupi_n_346, csa_tree_add_24_21_groupi_n_347, csa_tree_add_24_21_groupi_n_348, csa_tree_add_24_21_groupi_n_349, csa_tree_add_22_22_n_116, csa_tree_add_22_22_n_97;
  wire csa_tree_add_22_22_n_115, csa_tree_add_22_22_n_96, csa_tree_add_22_22_n_98, csa_tree_add_24_21_groupi_n_355, csa_tree_add_24_21_groupi_n_356, csa_tree_add_24_21_groupi_n_357, csa_tree_add_24_21_groupi_n_358, csa_tree_add_24_21_groupi_n_359;
  wire csa_tree_add_24_21_groupi_n_360, csa_tree_add_24_21_groupi_n_361, csa_tree_add_24_21_groupi_n_362, csa_tree_add_24_21_groupi_n_363, csa_tree_add_24_21_groupi_n_364, csa_tree_add_24_21_groupi_n_365, csa_tree_add_24_21_groupi_n_366, csa_tree_add_24_21_groupi_n_367;
  wire csa_tree_add_24_21_groupi_n_368, csa_tree_add_24_21_groupi_n_369, csa_tree_add_24_21_groupi_n_370, csa_tree_add_24_21_groupi_n_371, csa_tree_add_24_21_groupi_n_372, csa_tree_add_24_21_groupi_n_373, csa_tree_add_24_21_groupi_n_374, csa_tree_add_24_21_groupi_n_375;
  wire csa_tree_add_24_21_groupi_n_376, csa_tree_add_24_21_groupi_n_377, csa_tree_add_24_21_groupi_n_378, csa_tree_add_24_21_groupi_n_379, csa_tree_add_24_21_groupi_n_380, csa_tree_add_24_21_groupi_n_381, csa_tree_add_24_21_groupi_n_382, csa_tree_add_24_21_groupi_n_383;
  wire csa_tree_add_24_21_groupi_n_384, csa_tree_add_24_21_groupi_n_385, csa_tree_add_24_21_groupi_n_386, csa_tree_add_24_21_groupi_n_387, csa_tree_add_24_21_groupi_n_388, csa_tree_add_24_21_groupi_n_389, csa_tree_add_24_21_groupi_n_390, csa_tree_add_24_21_groupi_n_391;
  wire csa_tree_add_24_21_groupi_n_392, csa_tree_add_24_21_groupi_n_393, csa_tree_add_24_21_groupi_n_394, csa_tree_add_24_21_groupi_n_395, csa_tree_add_24_21_groupi_n_396, csa_tree_add_24_21_groupi_n_397, csa_tree_add_24_21_groupi_n_266, csa_tree_add_24_21_groupi_n_399;
  wire csa_tree_add_24_21_groupi_n_269, csa_tree_add_24_21_groupi_n_404, csa_tree_add_24_21_groupi_n_402, csa_tree_add_24_21_groupi_n_404, csa_tree_add_24_21_groupi_n_404, csa_tree_add_24_21_groupi_n_405, csa_tree_add_24_21_groupi_n_406, csa_tree_add_24_21_groupi_n_407;
  wire csa_tree_add_24_21_groupi_n_408, csa_tree_add_24_21_groupi_n_409, csa_tree_add_24_21_groupi_n_410, csa_tree_add_24_21_groupi_n_411, csa_tree_add_24_21_groupi_n_412, csa_tree_add_24_21_groupi_n_413, csa_tree_add_24_21_groupi_n_414, csa_tree_add_24_21_groupi_n_415;
  wire csa_tree_add_24_21_groupi_n_416, csa_tree_add_24_21_groupi_n_417, csa_tree_add_24_21_groupi_n_418, csa_tree_add_24_21_groupi_n_419, csa_tree_add_24_21_groupi_n_420, csa_tree_add_24_21_groupi_n_421, csa_tree_add_24_21_groupi_n_422, csa_tree_add_24_21_groupi_n_423;
  wire csa_tree_add_24_21_groupi_n_424, csa_tree_add_24_21_groupi_n_425, csa_tree_add_24_21_groupi_n_426, csa_tree_add_24_21_groupi_n_427, csa_tree_add_24_21_groupi_n_428, csa_tree_add_24_21_groupi_n_429, csa_tree_add_24_21_groupi_n_430, csa_tree_add_24_21_groupi_n_431;
  wire csa_tree_add_24_21_groupi_n_432, csa_tree_add_24_21_groupi_n_433, csa_tree_add_24_21_groupi_n_434, csa_tree_add_24_21_groupi_n_435, csa_tree_add_24_21_groupi_n_436, csa_tree_add_24_21_groupi_n_437, csa_tree_add_24_21_groupi_n_438, csa_tree_add_24_21_groupi_n_439;
  wire csa_tree_add_24_21_groupi_n_440, csa_tree_add_24_21_groupi_n_441, csa_tree_add_24_21_groupi_n_442, csa_tree_add_24_21_groupi_n_443, csa_tree_add_24_21_groupi_n_444, csa_tree_add_24_21_groupi_n_445, csa_tree_add_24_21_groupi_n_446, csa_tree_add_24_21_groupi_n_447;
  wire csa_tree_add_24_21_groupi_n_448, csa_tree_add_24_21_groupi_n_449, csa_tree_add_24_21_groupi_n_450, csa_tree_add_24_21_groupi_n_451, csa_tree_add_24_21_groupi_n_452, csa_tree_add_24_21_groupi_n_453, csa_tree_add_24_21_groupi_n_454, csa_tree_add_24_21_groupi_n_455;
  wire csa_tree_add_24_21_groupi_n_456, csa_tree_add_24_21_groupi_n_457, csa_tree_add_24_21_groupi_n_458, csa_tree_add_24_21_groupi_n_459, csa_tree_add_24_21_groupi_n_460, csa_tree_add_24_21_groupi_n_461, csa_tree_add_24_21_groupi_n_462, csa_tree_add_24_21_groupi_n_463;
  wire csa_tree_add_24_21_groupi_n_464, csa_tree_add_24_21_groupi_n_465, csa_tree_add_24_21_groupi_n_466, csa_tree_add_24_21_groupi_n_467, csa_tree_add_24_21_groupi_n_468, csa_tree_add_24_21_groupi_n_469, csa_tree_add_24_21_groupi_n_470, csa_tree_add_24_21_groupi_n_471;
  wire csa_tree_add_24_21_groupi_n_472, csa_tree_add_24_21_groupi_n_473, csa_tree_add_24_21_groupi_n_474, csa_tree_add_24_21_groupi_n_475, csa_tree_add_24_21_groupi_n_272, csa_tree_add_24_21_groupi_n_477, csa_tree_add_24_21_groupi_n_260, csa_tree_add_24_21_groupi_n_479;
  wire csa_tree_add_24_21_groupi_n_263, csa_tree_add_24_21_groupi_n_481, csa_tree_add_24_21_groupi_n_482, csa_tree_add_24_21_groupi_n_483, csa_tree_add_24_21_groupi_n_484, csa_tree_add_24_21_groupi_n_485, csa_tree_add_24_21_groupi_n_486, csa_tree_add_24_21_groupi_n_487;
  wire csa_tree_add_24_21_groupi_n_488, csa_tree_add_24_21_groupi_n_489, csa_tree_add_24_21_groupi_n_490, csa_tree_add_24_21_groupi_n_491, csa_tree_add_24_21_groupi_n_492, csa_tree_add_24_21_groupi_n_493, csa_tree_add_24_21_groupi_n_494, csa_tree_add_24_21_groupi_n_495;
  wire csa_tree_add_24_21_groupi_n_496, csa_tree_add_24_21_groupi_n_497, csa_tree_add_24_21_groupi_n_498, csa_tree_add_24_21_groupi_n_499, csa_tree_add_24_21_groupi_n_500, csa_tree_add_24_21_groupi_n_501, csa_tree_add_24_21_groupi_n_502, csa_tree_add_24_21_groupi_n_503;
  wire csa_tree_add_24_21_groupi_n_504, csa_tree_add_24_21_groupi_n_505, csa_tree_add_24_21_groupi_n_506, csa_tree_add_24_21_groupi_n_507, csa_tree_add_24_21_groupi_n_508, csa_tree_add_24_21_groupi_n_509, csa_tree_add_24_21_groupi_n_510, csa_tree_add_24_21_groupi_n_511;
  wire csa_tree_add_24_21_groupi_n_512, csa_tree_add_24_21_groupi_n_513, csa_tree_add_24_21_groupi_n_514, csa_tree_add_24_21_groupi_n_515, csa_tree_add_24_21_groupi_n_516, csa_tree_add_24_21_groupi_n_517, csa_tree_add_24_21_groupi_n_518, csa_tree_add_24_21_groupi_n_519;
  wire csa_tree_add_24_21_groupi_n_520, csa_tree_add_24_21_groupi_n_521, csa_tree_add_24_21_groupi_n_522, csa_tree_add_24_21_groupi_n_523, csa_tree_add_24_21_groupi_n_524, csa_tree_add_24_21_groupi_n_525, csa_tree_add_24_21_groupi_n_526, csa_tree_add_24_21_groupi_n_527;
  wire csa_tree_add_24_21_groupi_n_528, csa_tree_add_24_21_groupi_n_529, csa_tree_add_24_21_groupi_n_530, csa_tree_add_24_21_groupi_n_531, csa_tree_add_24_21_groupi_n_532, csa_tree_add_24_21_groupi_n_533, csa_tree_add_24_21_groupi_n_534, csa_tree_add_24_21_groupi_n_535;
  wire csa_tree_add_24_21_groupi_n_536, csa_tree_add_24_21_groupi_n_537, csa_tree_add_24_21_groupi_n_538, csa_tree_add_24_21_groupi_n_539, csa_tree_add_24_21_groupi_n_540, csa_tree_add_24_21_groupi_n_541, csa_tree_add_24_21_groupi_n_542, csa_tree_add_24_21_groupi_n_543;
  wire csa_tree_add_24_21_groupi_n_544, csa_tree_add_24_21_groupi_n_545, csa_tree_add_24_21_groupi_n_546, csa_tree_add_24_21_groupi_n_547, csa_tree_add_24_21_groupi_n_548, csa_tree_add_24_21_groupi_n_549, csa_tree_add_24_21_groupi_n_550, csa_tree_add_24_21_groupi_n_551;
  wire csa_tree_add_24_21_groupi_n_552, csa_tree_add_24_21_groupi_n_553, csa_tree_add_24_21_groupi_n_554, csa_tree_add_24_21_groupi_n_555, csa_tree_add_24_21_groupi_n_556, csa_tree_add_24_21_groupi_n_557, csa_tree_add_24_21_groupi_n_558, csa_tree_add_24_21_groupi_n_559;
  wire csa_tree_add_24_21_groupi_n_560, csa_tree_add_24_21_groupi_n_561, csa_tree_add_24_21_groupi_n_562, csa_tree_add_24_21_groupi_n_563, csa_tree_add_24_21_groupi_n_564, csa_tree_add_24_21_groupi_n_565, csa_tree_add_24_21_groupi_n_566, csa_tree_add_24_21_groupi_n_567;
  wire csa_tree_add_24_21_groupi_n_568, csa_tree_add_24_21_groupi_n_569, csa_tree_add_24_21_groupi_n_570, csa_tree_add_24_21_groupi_n_571, csa_tree_add_24_21_groupi_n_572, csa_tree_add_24_21_groupi_n_573, csa_tree_add_24_21_groupi_n_574, csa_tree_add_24_21_groupi_n_575;
  wire csa_tree_add_24_21_groupi_n_576, csa_tree_add_24_21_groupi_n_577, csa_tree_add_24_21_groupi_n_578, csa_tree_add_24_21_groupi_n_579, csa_tree_add_24_21_groupi_n_580, csa_tree_add_24_21_groupi_n_581, csa_tree_add_24_21_groupi_n_582, csa_tree_add_24_21_groupi_n_583;
  wire csa_tree_add_24_21_groupi_n_584, csa_tree_add_24_21_groupi_n_585, csa_tree_add_24_21_groupi_n_586, csa_tree_add_24_21_groupi_n_587, csa_tree_add_24_21_groupi_n_588, csa_tree_add_24_21_groupi_n_589, csa_tree_add_24_21_groupi_n_590, csa_tree_add_24_21_groupi_n_281;
  wire csa_tree_add_24_21_groupi_n_592, csa_tree_add_24_21_groupi_n_593, csa_tree_add_24_21_groupi_n_594, csa_tree_add_24_21_groupi_n_595, csa_tree_add_24_21_groupi_n_596, csa_tree_add_24_21_groupi_n_597, csa_tree_add_24_21_groupi_n_598, csa_tree_add_24_21_groupi_n_599;
  wire csa_tree_add_24_21_groupi_n_600, csa_tree_add_24_21_groupi_n_601, csa_tree_add_24_21_groupi_n_602, csa_tree_add_24_21_groupi_n_603, csa_tree_add_24_21_groupi_n_604, csa_tree_add_24_21_groupi_n_605, csa_tree_add_24_21_groupi_n_606, csa_tree_add_24_21_groupi_n_607;
  wire csa_tree_add_24_21_groupi_n_608, csa_tree_add_24_21_groupi_n_609, csa_tree_add_24_21_groupi_n_610, csa_tree_add_24_21_groupi_n_611, csa_tree_add_24_21_groupi_n_612, csa_tree_add_24_21_groupi_n_613, csa_tree_add_24_21_groupi_n_614, csa_tree_add_24_21_groupi_n_615;
  wire csa_tree_add_24_21_groupi_n_616, csa_tree_add_24_21_groupi_n_617, csa_tree_add_24_21_groupi_n_618, csa_tree_add_24_21_groupi_n_619, csa_tree_add_24_21_groupi_n_620, csa_tree_add_24_21_groupi_n_621, csa_tree_add_24_21_groupi_n_622, csa_tree_add_24_21_groupi_n_623;
  wire csa_tree_add_24_21_groupi_n_624, csa_tree_add_24_21_groupi_n_625, csa_tree_add_24_21_groupi_n_626, csa_tree_add_24_21_groupi_n_627, csa_tree_add_24_21_groupi_n_628, csa_tree_add_24_21_groupi_n_629, csa_tree_add_24_21_groupi_n_630, csa_tree_add_24_21_groupi_n_631;
  wire csa_tree_add_24_21_groupi_n_632, csa_tree_add_24_21_groupi_n_633, csa_tree_add_24_21_groupi_n_634, csa_tree_add_24_21_groupi_n_635, csa_tree_add_24_21_groupi_n_636, csa_tree_add_24_21_groupi_n_637, csa_tree_add_24_21_groupi_n_638, csa_tree_add_24_21_groupi_n_639;
  wire csa_tree_add_24_21_groupi_n_640, csa_tree_add_24_21_groupi_n_641, csa_tree_add_24_21_groupi_n_642, csa_tree_add_24_21_groupi_n_643, csa_tree_add_24_21_groupi_n_644, csa_tree_add_24_21_groupi_n_645, csa_tree_add_24_21_groupi_n_646, csa_tree_add_24_21_groupi_n_647;
  wire csa_tree_add_24_21_groupi_n_648, csa_tree_add_24_21_groupi_n_649, csa_tree_add_24_21_groupi_n_650, csa_tree_add_24_21_groupi_n_651, csa_tree_add_24_21_groupi_n_652, csa_tree_add_24_21_groupi_n_653, csa_tree_add_24_21_groupi_n_654, csa_tree_add_24_21_groupi_n_655;
  wire csa_tree_add_24_21_groupi_n_656, csa_tree_add_24_21_groupi_n_657, csa_tree_add_24_21_groupi_n_658, csa_tree_add_24_21_groupi_n_659, csa_tree_add_24_21_groupi_n_660, csa_tree_add_24_21_groupi_n_661, csa_tree_add_24_21_groupi_n_662, csa_tree_add_24_21_groupi_n_663;
  wire csa_tree_add_24_21_groupi_n_664, csa_tree_add_24_21_groupi_n_665, csa_tree_add_24_21_groupi_n_666, csa_tree_add_24_21_groupi_n_667, csa_tree_add_24_21_groupi_n_668, csa_tree_add_24_21_groupi_n_669, csa_tree_add_24_21_groupi_n_670, csa_tree_add_24_21_groupi_n_671;
  wire csa_tree_add_24_21_groupi_n_672, csa_tree_add_24_21_groupi_n_673, csa_tree_add_24_21_groupi_n_674, csa_tree_add_24_21_groupi_n_675, csa_tree_add_24_21_groupi_n_676, csa_tree_add_24_21_groupi_n_677, csa_tree_add_24_21_groupi_n_678, csa_tree_add_24_21_groupi_n_679;
  wire csa_tree_add_24_21_groupi_n_680, csa_tree_add_24_21_groupi_n_681, csa_tree_add_24_21_groupi_n_682, csa_tree_add_24_21_groupi_n_683, csa_tree_add_24_21_groupi_n_684, csa_tree_add_24_21_groupi_n_685, csa_tree_add_24_21_groupi_n_686, csa_tree_add_24_21_groupi_n_687;
  wire csa_tree_add_24_21_groupi_n_688, csa_tree_add_24_21_groupi_n_689, csa_tree_add_24_21_groupi_n_690, csa_tree_add_24_21_groupi_n_691, csa_tree_add_24_21_groupi_n_692, csa_tree_add_24_21_groupi_n_693, csa_tree_add_24_21_groupi_n_694, csa_tree_add_24_21_groupi_n_695;
  wire csa_tree_add_24_21_groupi_n_696, csa_tree_add_24_21_groupi_n_697, csa_tree_add_24_21_groupi_n_698, csa_tree_add_24_21_groupi_n_699, csa_tree_add_24_21_groupi_n_700, csa_tree_add_24_21_groupi_n_701, csa_tree_add_24_21_groupi_n_702, csa_tree_add_24_21_groupi_n_703;
  wire csa_tree_add_24_21_groupi_n_704, csa_tree_add_24_21_groupi_n_705, csa_tree_add_24_21_groupi_n_706, csa_tree_add_24_21_groupi_n_707, csa_tree_add_24_21_groupi_n_708, csa_tree_add_24_21_groupi_n_709, csa_tree_add_24_21_groupi_n_710, csa_tree_add_24_21_groupi_n_711;
  wire csa_tree_add_24_21_groupi_n_712, csa_tree_add_24_21_groupi_n_713, csa_tree_add_24_21_groupi_n_714, csa_tree_add_24_21_groupi_n_715, csa_tree_add_24_21_groupi_n_716, csa_tree_add_24_21_groupi_n_717, csa_tree_add_24_21_groupi_n_718, csa_tree_add_24_21_groupi_n_719;
  wire csa_tree_add_24_21_groupi_n_720, csa_tree_add_24_21_groupi_n_721, csa_tree_add_24_21_groupi_n_722, csa_tree_add_24_21_groupi_n_723, csa_tree_add_24_21_groupi_n_724, csa_tree_add_24_21_groupi_n_725, csa_tree_add_24_21_groupi_n_726, csa_tree_add_24_21_groupi_n_727;
  wire csa_tree_add_24_21_groupi_n_728, csa_tree_add_24_21_groupi_n_729, csa_tree_add_24_21_groupi_n_730, csa_tree_add_24_21_groupi_n_731, csa_tree_add_24_21_groupi_n_732, csa_tree_add_24_21_groupi_n_733, csa_tree_add_24_21_groupi_n_734, csa_tree_add_24_21_groupi_n_735;
  wire csa_tree_add_24_21_groupi_n_736, csa_tree_add_24_21_groupi_n_737, csa_tree_add_24_21_groupi_n_738, csa_tree_add_24_21_groupi_n_739, csa_tree_add_24_21_groupi_n_740, csa_tree_add_24_21_groupi_n_741, csa_tree_add_24_21_groupi_n_742, csa_tree_add_24_21_groupi_n_743;
  wire csa_tree_add_24_21_groupi_n_744, csa_tree_add_24_21_groupi_n_745, csa_tree_add_24_21_groupi_n_746, csa_tree_add_24_21_groupi_n_747, csa_tree_add_24_21_groupi_n_748, csa_tree_add_24_21_groupi_n_749, csa_tree_add_24_21_groupi_n_750, csa_tree_add_24_21_groupi_n_751;
  wire csa_tree_add_24_21_groupi_n_752, csa_tree_add_24_21_groupi_n_753, csa_tree_add_24_21_groupi_n_754, csa_tree_add_24_21_groupi_n_755, csa_tree_add_24_21_groupi_n_756, csa_tree_add_24_21_groupi_n_757, csa_tree_add_24_21_groupi_n_758, csa_tree_add_24_21_groupi_n_759;
  wire csa_tree_add_24_21_groupi_n_760, csa_tree_add_24_21_groupi_n_761, csa_tree_add_24_21_groupi_n_762, csa_tree_add_24_21_groupi_n_763, csa_tree_add_24_21_groupi_n_764, csa_tree_add_24_21_groupi_n_765, csa_tree_add_24_21_groupi_n_766, csa_tree_add_24_21_groupi_n_767;
  wire csa_tree_add_24_21_groupi_n_768, csa_tree_add_24_21_groupi_n_769, csa_tree_add_24_21_groupi_n_770, csa_tree_add_24_21_groupi_n_771, csa_tree_add_24_21_groupi_n_772, csa_tree_add_24_21_groupi_n_773, csa_tree_add_24_21_groupi_n_774, csa_tree_add_24_21_groupi_n_775;
  wire csa_tree_add_24_21_groupi_n_776, csa_tree_add_24_21_groupi_n_777, csa_tree_add_24_21_groupi_n_778, csa_tree_add_24_21_groupi_n_779, csa_tree_add_24_21_groupi_n_780, csa_tree_add_24_21_groupi_n_781, csa_tree_add_24_21_groupi_n_782, csa_tree_add_24_21_groupi_n_783;
  wire csa_tree_add_24_21_groupi_n_784, csa_tree_add_24_21_groupi_n_785, csa_tree_add_24_21_groupi_n_786, csa_tree_add_24_21_groupi_n_787, csa_tree_add_24_21_groupi_n_788, csa_tree_add_24_21_groupi_n_789, csa_tree_add_24_21_groupi_n_790, csa_tree_add_24_21_groupi_n_791;
  wire csa_tree_add_24_21_groupi_n_792, csa_tree_add_24_21_groupi_n_793, csa_tree_add_24_21_groupi_n_794, csa_tree_add_24_21_groupi_n_795, csa_tree_add_24_21_groupi_n_796, csa_tree_add_24_21_groupi_n_797, csa_tree_add_24_21_groupi_n_798, csa_tree_add_24_21_groupi_n_799;
  wire csa_tree_add_24_21_groupi_n_800, csa_tree_add_24_21_groupi_n_801, csa_tree_add_24_21_groupi_n_802, csa_tree_add_24_21_groupi_n_803, csa_tree_add_24_21_groupi_n_804, csa_tree_add_24_21_groupi_n_805, csa_tree_add_24_21_groupi_n_806, csa_tree_add_24_21_groupi_n_807;
  wire csa_tree_add_24_21_groupi_n_808, csa_tree_add_24_21_groupi_n_809, csa_tree_add_24_21_groupi_n_810, csa_tree_add_24_21_groupi_n_811, csa_tree_add_24_21_groupi_n_812, csa_tree_add_24_21_groupi_n_813, csa_tree_add_24_21_groupi_n_814, csa_tree_add_24_21_groupi_n_815;
  wire csa_tree_add_24_21_groupi_n_816, csa_tree_add_24_21_groupi_n_817, csa_tree_add_24_21_groupi_n_818, csa_tree_add_24_21_groupi_n_819, csa_tree_add_24_21_groupi_n_820, csa_tree_add_24_21_groupi_n_821, csa_tree_add_24_21_groupi_n_822, csa_tree_add_24_21_groupi_n_823;
  wire csa_tree_add_24_21_groupi_n_824, csa_tree_add_24_21_groupi_n_825, csa_tree_add_24_21_groupi_n_826, csa_tree_add_24_21_groupi_n_827, csa_tree_add_24_21_groupi_n_828, csa_tree_add_24_21_groupi_n_829, csa_tree_add_24_21_groupi_n_830, csa_tree_add_24_21_groupi_n_831;
  wire csa_tree_add_24_21_groupi_n_832, csa_tree_add_24_21_groupi_n_833, csa_tree_add_24_21_groupi_n_834, csa_tree_add_24_21_groupi_n_835, csa_tree_add_24_21_groupi_n_836, csa_tree_add_24_21_groupi_n_837, csa_tree_add_24_21_groupi_n_838, csa_tree_add_24_21_groupi_n_839;
  wire csa_tree_add_24_21_groupi_n_840, csa_tree_add_24_21_groupi_n_841, csa_tree_add_24_21_groupi_n_842, csa_tree_add_24_21_groupi_n_843, csa_tree_add_24_21_groupi_n_844, csa_tree_add_24_21_groupi_n_845, csa_tree_add_24_21_groupi_n_846, csa_tree_add_24_21_groupi_n_847;
  wire csa_tree_add_24_21_groupi_n_848, csa_tree_add_24_21_groupi_n_849, csa_tree_add_24_21_groupi_n_850, csa_tree_add_24_21_groupi_n_851, csa_tree_add_24_21_groupi_n_852, csa_tree_add_24_21_groupi_n_853, csa_tree_add_24_21_groupi_n_854, csa_tree_add_24_21_groupi_n_855;
  wire csa_tree_add_24_21_groupi_n_856, csa_tree_add_24_21_groupi_n_857, csa_tree_add_24_21_groupi_n_858, csa_tree_add_24_21_groupi_n_859, csa_tree_add_24_21_groupi_n_860, csa_tree_add_24_21_groupi_n_861, csa_tree_add_24_21_groupi_n_862, csa_tree_add_24_21_groupi_n_863;
  wire csa_tree_add_24_21_groupi_n_864, csa_tree_add_24_21_groupi_n_865, csa_tree_add_24_21_groupi_n_866, csa_tree_add_24_21_groupi_n_867, csa_tree_add_24_21_groupi_n_868, csa_tree_add_24_21_groupi_n_869, csa_tree_add_24_21_groupi_n_870, csa_tree_add_24_21_groupi_n_871;
  wire csa_tree_add_24_21_groupi_n_872, csa_tree_add_24_21_groupi_n_873, csa_tree_add_24_21_groupi_n_874, csa_tree_add_24_21_groupi_n_875, csa_tree_add_24_21_groupi_n_876, csa_tree_add_24_21_groupi_n_877, csa_tree_add_24_21_groupi_n_878, csa_tree_add_24_21_groupi_n_879;
  wire csa_tree_add_24_21_groupi_n_880, csa_tree_add_24_21_groupi_n_881, csa_tree_add_24_21_groupi_n_882, csa_tree_add_24_21_groupi_n_883, csa_tree_add_24_21_groupi_n_884, csa_tree_add_24_21_groupi_n_885, csa_tree_add_24_21_groupi_n_886, csa_tree_add_24_21_groupi_n_887;
  wire csa_tree_add_24_21_groupi_n_888, csa_tree_add_24_21_groupi_n_889, csa_tree_add_24_21_groupi_n_890, csa_tree_add_24_21_groupi_n_891, csa_tree_add_24_21_groupi_n_892, csa_tree_add_24_21_groupi_n_893, csa_tree_add_24_21_groupi_n_894, csa_tree_add_24_21_groupi_n_895;
  wire csa_tree_add_24_21_groupi_n_896, csa_tree_add_24_21_groupi_n_897, csa_tree_add_24_21_groupi_n_898, csa_tree_add_24_21_groupi_n_899, csa_tree_add_24_21_groupi_n_900, csa_tree_add_24_21_groupi_n_901, csa_tree_add_24_21_groupi_n_902, csa_tree_add_24_21_groupi_n_903;
  wire csa_tree_add_24_21_groupi_n_904, csa_tree_add_24_21_groupi_n_905, csa_tree_add_24_21_groupi_n_906, csa_tree_add_24_21_groupi_n_907, csa_tree_add_24_21_groupi_n_908, csa_tree_add_24_21_groupi_n_909, csa_tree_add_24_21_groupi_n_910, csa_tree_add_24_21_groupi_n_911;
  wire csa_tree_add_24_21_groupi_n_912, csa_tree_add_24_21_groupi_n_913, csa_tree_add_24_21_groupi_n_914, csa_tree_add_24_21_groupi_n_915, csa_tree_add_24_21_groupi_n_916, csa_tree_add_24_21_groupi_n_917, csa_tree_add_24_21_groupi_n_918, csa_tree_add_24_21_groupi_n_919;
  wire csa_tree_add_24_21_groupi_n_920, csa_tree_add_24_21_groupi_n_921, csa_tree_add_24_21_groupi_n_922, csa_tree_add_24_21_groupi_n_923, csa_tree_add_24_21_groupi_n_924, csa_tree_add_24_21_groupi_n_925, csa_tree_add_24_21_groupi_n_926, csa_tree_add_24_21_groupi_n_927;
  wire csa_tree_add_24_21_groupi_n_928, csa_tree_add_24_21_groupi_n_929, csa_tree_add_24_21_groupi_n_930, csa_tree_add_24_21_groupi_n_931, csa_tree_add_24_21_groupi_n_932, csa_tree_add_24_21_groupi_n_933, csa_tree_add_24_21_groupi_n_934, csa_tree_add_24_21_groupi_n_935;
  wire csa_tree_add_24_21_groupi_n_936, csa_tree_add_24_21_groupi_n_937, csa_tree_add_24_21_groupi_n_938, csa_tree_add_24_21_groupi_n_939, csa_tree_add_24_21_groupi_n_940, csa_tree_add_24_21_groupi_n_941, csa_tree_add_24_21_groupi_n_942, csa_tree_add_24_21_groupi_n_943;
  wire csa_tree_add_24_21_groupi_n_944, csa_tree_add_24_21_groupi_n_945, csa_tree_add_24_21_groupi_n_946, csa_tree_add_24_21_groupi_n_947, csa_tree_add_24_21_groupi_n_948, csa_tree_add_24_21_groupi_n_949, csa_tree_add_24_21_groupi_n_950, csa_tree_add_24_21_groupi_n_951;
  wire csa_tree_add_24_21_groupi_n_952, csa_tree_add_24_21_groupi_n_953, csa_tree_add_24_21_groupi_n_954, csa_tree_add_24_21_groupi_n_955, csa_tree_add_24_21_groupi_n_956, csa_tree_add_24_21_groupi_n_957, csa_tree_add_24_21_groupi_n_958, csa_tree_add_24_21_groupi_n_959;
  wire csa_tree_add_24_21_groupi_n_960, csa_tree_add_24_21_groupi_n_961, csa_tree_add_24_21_groupi_n_962, csa_tree_add_24_21_groupi_n_963, csa_tree_add_24_21_groupi_n_964, csa_tree_add_24_21_groupi_n_965, csa_tree_add_24_21_groupi_n_966, csa_tree_add_24_21_groupi_n_967;
  wire csa_tree_add_24_21_groupi_n_968, csa_tree_add_24_21_groupi_n_969, csa_tree_add_24_21_groupi_n_970, csa_tree_add_24_21_groupi_n_971, csa_tree_add_24_21_groupi_n_972, csa_tree_add_24_21_groupi_n_973, csa_tree_add_24_21_groupi_n_974, csa_tree_add_24_21_groupi_n_975;
  wire csa_tree_add_24_21_groupi_n_976, csa_tree_add_24_21_groupi_n_977, csa_tree_add_24_21_groupi_n_978, csa_tree_add_24_21_groupi_n_979, csa_tree_add_24_21_groupi_n_980, csa_tree_add_24_21_groupi_n_981, csa_tree_add_24_21_groupi_n_982, csa_tree_add_24_21_groupi_n_983;
  wire csa_tree_add_24_21_groupi_n_984, csa_tree_add_24_21_groupi_n_985, csa_tree_add_24_21_groupi_n_986, csa_tree_add_24_21_groupi_n_987, csa_tree_add_24_21_groupi_n_988, csa_tree_add_24_21_groupi_n_989, csa_tree_add_24_21_groupi_n_990, csa_tree_add_24_21_groupi_n_991;
  wire csa_tree_add_24_21_groupi_n_992, csa_tree_add_24_21_groupi_n_993, csa_tree_add_24_21_groupi_n_994, csa_tree_add_24_21_groupi_n_995, csa_tree_add_24_21_groupi_n_996, csa_tree_add_24_21_groupi_n_997, csa_tree_add_24_21_groupi_n_998, csa_tree_add_24_21_groupi_n_999;
  wire csa_tree_add_24_21_groupi_n_1000, csa_tree_add_24_21_groupi_n_1001, csa_tree_add_24_21_groupi_n_1002, csa_tree_add_24_21_groupi_n_1003, csa_tree_add_24_21_groupi_n_1004, csa_tree_add_24_21_groupi_n_1005, csa_tree_add_24_21_groupi_n_1006, csa_tree_add_24_21_groupi_n_1007;
  wire csa_tree_add_24_21_groupi_n_1008, csa_tree_add_24_21_groupi_n_1009, csa_tree_add_24_21_groupi_n_1010, csa_tree_add_24_21_groupi_n_1011, csa_tree_add_24_21_groupi_n_1012, csa_tree_add_24_21_groupi_n_1013, csa_tree_add_24_21_groupi_n_1014, csa_tree_add_24_21_groupi_n_1015;
  wire csa_tree_add_24_21_groupi_n_1016, csa_tree_add_24_21_groupi_n_1017, csa_tree_add_24_21_groupi_n_1018, csa_tree_add_24_21_groupi_n_1019, csa_tree_add_24_21_groupi_n_1020, csa_tree_add_24_21_groupi_n_1021, csa_tree_add_24_21_groupi_n_1022, csa_tree_add_24_21_groupi_n_1023;
  wire csa_tree_add_24_21_groupi_n_1024, csa_tree_add_24_21_groupi_n_1025, csa_tree_add_24_21_groupi_n_1026, csa_tree_add_24_21_groupi_n_1027, csa_tree_add_24_21_groupi_n_1028, csa_tree_add_24_21_groupi_n_1029, csa_tree_add_24_21_groupi_n_1030, csa_tree_add_24_21_groupi_n_1031;
  wire csa_tree_add_24_21_groupi_n_1032, csa_tree_add_24_21_groupi_n_1033, csa_tree_add_24_21_groupi_n_1034, csa_tree_add_24_21_groupi_n_1035, csa_tree_add_24_21_groupi_n_1036, csa_tree_add_24_21_groupi_n_1037, csa_tree_add_24_21_groupi_n_1038, csa_tree_add_24_21_groupi_n_1039;
  wire csa_tree_add_24_21_groupi_n_1040, csa_tree_add_24_21_groupi_n_1041, csa_tree_add_24_21_groupi_n_1042, csa_tree_add_24_21_groupi_n_1043, csa_tree_add_24_21_groupi_n_1044, csa_tree_add_24_21_groupi_n_1045, csa_tree_add_24_21_groupi_n_1046, csa_tree_add_24_21_groupi_n_1047;
  wire csa_tree_add_24_21_groupi_n_1048, csa_tree_add_24_21_groupi_n_1049, csa_tree_add_24_21_groupi_n_1050, csa_tree_add_24_21_groupi_n_1051, csa_tree_add_24_21_groupi_n_1052, csa_tree_add_24_21_groupi_n_1053, csa_tree_add_24_21_groupi_n_1054, csa_tree_add_24_21_groupi_n_1055;
  wire csa_tree_add_24_21_groupi_n_1056, csa_tree_add_24_21_groupi_n_1057, csa_tree_add_24_21_groupi_n_1058, csa_tree_add_24_21_groupi_n_1059, csa_tree_add_24_21_groupi_n_1060, csa_tree_add_24_21_groupi_n_1061, csa_tree_add_24_21_groupi_n_1062, csa_tree_add_24_21_groupi_n_1063;
  wire csa_tree_add_24_21_groupi_n_1064, csa_tree_add_24_21_groupi_n_1065, csa_tree_add_24_21_groupi_n_1066, csa_tree_add_24_21_groupi_n_1067, csa_tree_add_24_21_groupi_n_1068, csa_tree_add_24_21_groupi_n_1069, csa_tree_add_24_21_groupi_n_1070, csa_tree_add_24_21_groupi_n_1071;
  wire csa_tree_add_24_21_groupi_n_1072, csa_tree_add_24_21_groupi_n_1073, csa_tree_add_24_21_groupi_n_1074, csa_tree_add_24_21_groupi_n_1075, csa_tree_add_24_21_groupi_n_1076, csa_tree_add_24_21_groupi_n_1077, csa_tree_add_24_21_groupi_n_1078, csa_tree_add_24_21_groupi_n_1079;
  wire csa_tree_add_24_21_groupi_n_1080, csa_tree_add_24_21_groupi_n_1081, csa_tree_add_24_21_groupi_n_1082, csa_tree_add_24_21_groupi_n_1083, csa_tree_add_24_21_groupi_n_1084, csa_tree_add_24_21_groupi_n_1085, csa_tree_add_24_21_groupi_n_1086, csa_tree_add_24_21_groupi_n_1087;
  wire csa_tree_add_24_21_groupi_n_1088, csa_tree_add_24_21_groupi_n_1089, csa_tree_add_24_21_groupi_n_1090, csa_tree_add_24_21_groupi_n_1091, csa_tree_add_24_21_groupi_n_1092, csa_tree_add_24_21_groupi_n_1093, csa_tree_add_24_21_groupi_n_1094, csa_tree_add_24_21_groupi_n_1095;
  wire csa_tree_add_24_21_groupi_n_1096, csa_tree_add_24_21_groupi_n_1097, csa_tree_add_24_21_groupi_n_1098, csa_tree_add_24_21_groupi_n_1099, csa_tree_add_24_21_groupi_n_1100, csa_tree_add_24_21_groupi_n_1101, csa_tree_add_24_21_groupi_n_1102, csa_tree_add_24_21_groupi_n_1103;
  wire csa_tree_add_24_21_groupi_n_1104, csa_tree_add_24_21_groupi_n_1105, csa_tree_add_24_21_groupi_n_1106, csa_tree_add_24_21_groupi_n_1107, csa_tree_add_24_21_groupi_n_1108, csa_tree_add_24_21_groupi_n_1109, csa_tree_add_24_21_groupi_n_1110, csa_tree_add_24_21_groupi_n_1111;
  wire csa_tree_add_24_21_groupi_n_1112, csa_tree_add_24_21_groupi_n_1113, csa_tree_add_24_21_groupi_n_1114, csa_tree_add_24_21_groupi_n_1115, csa_tree_add_24_21_groupi_n_1116, csa_tree_add_24_21_groupi_n_1117, csa_tree_add_24_21_groupi_n_1118, csa_tree_add_24_21_groupi_n_1119;
  wire csa_tree_add_24_21_groupi_n_1120, csa_tree_add_24_21_groupi_n_1121, csa_tree_add_24_21_groupi_n_1122, csa_tree_add_24_21_groupi_n_1123, csa_tree_add_24_21_groupi_n_1124, csa_tree_add_24_21_groupi_n_1125, csa_tree_add_24_21_groupi_n_1126, csa_tree_add_24_21_groupi_n_1127;
  wire csa_tree_add_24_21_groupi_n_1128, csa_tree_add_24_21_groupi_n_1129, csa_tree_add_24_21_groupi_n_1130, csa_tree_add_24_21_groupi_n_1131, csa_tree_add_24_21_groupi_n_1132, csa_tree_add_24_21_groupi_n_1133, csa_tree_add_24_21_groupi_n_1134, csa_tree_add_24_21_groupi_n_1135;
  wire csa_tree_add_24_21_groupi_n_1136, csa_tree_add_24_21_groupi_n_1137, csa_tree_add_24_21_groupi_n_1138, csa_tree_add_24_21_groupi_n_1139, csa_tree_add_24_21_groupi_n_1140, csa_tree_add_24_21_groupi_n_1141, csa_tree_add_24_21_groupi_n_1142, csa_tree_add_24_21_groupi_n_1143;
  wire csa_tree_add_24_21_groupi_n_1144, csa_tree_add_24_21_groupi_n_1145, csa_tree_add_24_21_groupi_n_1146, csa_tree_add_24_21_groupi_n_1147, csa_tree_add_24_21_groupi_n_1148, csa_tree_add_24_21_groupi_n_1149, csa_tree_add_24_21_groupi_n_1150, csa_tree_add_24_21_groupi_n_1151;
  wire csa_tree_add_24_21_groupi_n_1152, csa_tree_add_24_21_groupi_n_1153, csa_tree_add_24_21_groupi_n_1154, csa_tree_add_24_21_groupi_n_1155, csa_tree_add_24_21_groupi_n_1156, csa_tree_add_24_21_groupi_n_1157, csa_tree_add_24_21_groupi_n_1158, csa_tree_add_24_21_groupi_n_1159;
  wire csa_tree_add_24_21_groupi_n_1160, csa_tree_add_24_21_groupi_n_1161, csa_tree_add_24_21_groupi_n_1162, csa_tree_add_24_21_groupi_n_1163, csa_tree_add_24_21_groupi_n_1164, csa_tree_add_24_21_groupi_n_1165, csa_tree_add_24_21_groupi_n_1166, csa_tree_add_24_21_groupi_n_1167;
  wire csa_tree_add_24_21_groupi_n_1168, csa_tree_add_24_21_groupi_n_1169, csa_tree_add_24_21_groupi_n_1170, csa_tree_add_24_21_groupi_n_1171, csa_tree_add_24_21_groupi_n_1172, csa_tree_add_24_21_groupi_n_1173, csa_tree_add_24_21_groupi_n_1174, csa_tree_add_24_21_groupi_n_1175;
  wire csa_tree_add_24_21_groupi_n_1176, csa_tree_add_24_21_groupi_n_1177, csa_tree_add_24_21_groupi_n_1178, csa_tree_add_24_21_groupi_n_1179, csa_tree_add_24_21_groupi_n_1180, csa_tree_add_24_21_groupi_n_1181, csa_tree_add_24_21_groupi_n_1182, csa_tree_add_24_21_groupi_n_1183;
  wire csa_tree_add_24_21_groupi_n_1184, csa_tree_add_24_21_groupi_n_1185, csa_tree_add_24_21_groupi_n_1186, csa_tree_add_24_21_groupi_n_1187, csa_tree_add_24_21_groupi_n_1188, csa_tree_add_24_21_groupi_n_1189, csa_tree_add_24_21_groupi_n_1190, csa_tree_add_24_21_groupi_n_1191;
  wire csa_tree_add_24_21_groupi_n_1192, csa_tree_add_24_21_groupi_n_1193, csa_tree_add_24_21_groupi_n_1194, csa_tree_add_24_21_groupi_n_1195, csa_tree_add_24_21_groupi_n_1196, csa_tree_add_24_21_groupi_n_1197, csa_tree_add_24_21_groupi_n_1198, csa_tree_add_24_21_groupi_n_1199;
  wire csa_tree_add_24_21_groupi_n_1200, csa_tree_add_24_21_groupi_n_1201, csa_tree_add_24_21_groupi_n_1202, csa_tree_add_24_21_groupi_n_1203, csa_tree_add_24_21_groupi_n_1204, csa_tree_add_24_21_groupi_n_1205, csa_tree_add_24_21_groupi_n_1206, csa_tree_add_24_21_groupi_n_1207;
  wire csa_tree_add_24_21_groupi_n_1208, csa_tree_add_24_21_groupi_n_1209, csa_tree_add_24_21_groupi_n_1210, csa_tree_add_24_21_groupi_n_1211, csa_tree_add_24_21_groupi_n_1212, csa_tree_add_24_21_groupi_n_1213, csa_tree_add_24_21_groupi_n_1214, csa_tree_add_24_21_groupi_n_1215;
  wire csa_tree_add_24_21_groupi_n_1216, csa_tree_add_24_21_groupi_n_1217, csa_tree_add_24_21_groupi_n_1218, csa_tree_add_24_21_groupi_n_1219, csa_tree_add_24_21_groupi_n_1220, csa_tree_add_24_21_groupi_n_1221, csa_tree_add_24_21_groupi_n_1222, csa_tree_add_24_21_groupi_n_1223;
  wire csa_tree_add_24_21_groupi_n_1224, csa_tree_add_24_21_groupi_n_1225, csa_tree_add_24_21_groupi_n_1226, csa_tree_add_24_21_groupi_n_1227, csa_tree_add_24_21_groupi_n_1228, csa_tree_add_24_21_groupi_n_1229, csa_tree_add_24_21_groupi_n_1230, csa_tree_add_24_21_groupi_n_1231;
  wire csa_tree_add_24_21_groupi_n_1232, csa_tree_add_24_21_groupi_n_1233, csa_tree_add_24_21_groupi_n_1234, csa_tree_add_24_21_groupi_n_1235, csa_tree_add_24_21_groupi_n_1236, csa_tree_add_24_21_groupi_n_1237, csa_tree_add_24_21_groupi_n_1238, csa_tree_add_24_21_groupi_n_1239;
  wire csa_tree_add_24_21_groupi_n_1240, csa_tree_add_24_21_groupi_n_1241, csa_tree_add_24_21_groupi_n_1242, csa_tree_add_24_21_groupi_n_1243, csa_tree_add_24_21_groupi_n_1244, csa_tree_add_24_21_groupi_n_1245, csa_tree_add_24_21_groupi_n_1246, csa_tree_add_24_21_groupi_n_1247;
  wire csa_tree_add_24_21_groupi_n_1248, csa_tree_add_24_21_groupi_n_1249, csa_tree_add_24_21_groupi_n_1250, csa_tree_add_24_21_groupi_n_1251, csa_tree_add_24_21_groupi_n_1252, csa_tree_add_24_21_groupi_n_1253, csa_tree_add_24_21_groupi_n_1254, csa_tree_add_24_21_groupi_n_1255;
  wire csa_tree_add_24_21_groupi_n_1256, csa_tree_add_24_21_groupi_n_1257, csa_tree_add_24_21_groupi_n_1258, csa_tree_add_24_21_groupi_n_1259, csa_tree_add_24_21_groupi_n_1260, csa_tree_add_24_21_groupi_n_1261, csa_tree_add_24_21_groupi_n_1262, csa_tree_add_24_21_groupi_n_1263;
  wire csa_tree_add_24_21_groupi_n_1264, csa_tree_add_24_21_groupi_n_1265, csa_tree_add_24_21_groupi_n_1266, csa_tree_add_24_21_groupi_n_1267, csa_tree_add_24_21_groupi_n_1268, csa_tree_add_24_21_groupi_n_1269, csa_tree_add_24_21_groupi_n_1270, csa_tree_add_24_21_groupi_n_1271;
  wire csa_tree_add_24_21_groupi_n_1272, csa_tree_add_24_21_groupi_n_1273, csa_tree_add_24_21_groupi_n_1274, csa_tree_add_24_21_groupi_n_1275, csa_tree_add_24_21_groupi_n_1276, csa_tree_add_24_21_groupi_n_1277, csa_tree_add_24_21_groupi_n_1278, csa_tree_add_24_21_groupi_n_1279;
  wire csa_tree_add_24_21_groupi_n_1280, csa_tree_add_24_21_groupi_n_1281, csa_tree_add_24_21_groupi_n_1282, csa_tree_add_24_21_groupi_n_1283, csa_tree_add_24_21_groupi_n_1284, csa_tree_add_24_21_groupi_n_1285, csa_tree_add_24_21_groupi_n_1286, csa_tree_add_24_21_groupi_n_1287;
  wire csa_tree_add_24_21_groupi_n_1288, csa_tree_add_24_21_groupi_n_1289, csa_tree_add_24_21_groupi_n_1290, csa_tree_add_24_21_groupi_n_1291, csa_tree_add_24_21_groupi_n_1292, csa_tree_add_24_21_groupi_n_1293, csa_tree_add_24_21_groupi_n_1294, csa_tree_add_24_21_groupi_n_1295;
  wire csa_tree_add_24_21_groupi_n_1296, csa_tree_add_24_21_groupi_n_1297, csa_tree_add_24_21_groupi_n_1298, csa_tree_add_24_21_groupi_n_1299, csa_tree_add_24_21_groupi_n_1300, csa_tree_add_24_21_groupi_n_1301, csa_tree_add_24_21_groupi_n_1302, csa_tree_add_24_21_groupi_n_1303;
  wire csa_tree_add_24_21_groupi_n_1304, csa_tree_add_24_21_groupi_n_1305, csa_tree_add_24_21_groupi_n_1306, csa_tree_add_24_21_groupi_n_1307, csa_tree_add_24_21_groupi_n_1308, csa_tree_add_24_21_groupi_n_1309, csa_tree_add_24_21_groupi_n_1310, csa_tree_add_24_21_groupi_n_1311;
  wire csa_tree_add_24_21_groupi_n_1312, csa_tree_add_24_21_groupi_n_1313, csa_tree_add_24_21_groupi_n_1314, csa_tree_add_24_21_groupi_n_1315, csa_tree_add_24_21_groupi_n_1316, csa_tree_add_24_21_groupi_n_1317, csa_tree_add_24_21_groupi_n_1318, csa_tree_add_24_21_groupi_n_1319;
  wire csa_tree_add_24_21_groupi_n_1320, csa_tree_add_24_21_groupi_n_1321, csa_tree_add_24_21_groupi_n_1322, csa_tree_add_24_21_groupi_n_1323, csa_tree_add_24_21_groupi_n_1324, csa_tree_add_24_21_groupi_n_1325, csa_tree_add_24_21_groupi_n_1326, csa_tree_add_24_21_groupi_n_1327;
  wire csa_tree_add_24_21_groupi_n_1328, csa_tree_add_24_21_groupi_n_1329, csa_tree_add_24_21_groupi_n_1330, csa_tree_add_24_21_groupi_n_1331, csa_tree_add_24_21_groupi_n_1332, csa_tree_add_24_21_groupi_n_1333, csa_tree_add_24_21_groupi_n_1334, csa_tree_add_24_21_groupi_n_1335;
  wire csa_tree_add_24_21_groupi_n_1336, csa_tree_add_24_21_groupi_n_1337, csa_tree_add_24_21_groupi_n_1338, csa_tree_add_24_21_groupi_n_1339, csa_tree_add_24_21_groupi_n_1340, csa_tree_add_24_21_groupi_n_1341, csa_tree_add_24_21_groupi_n_1342, csa_tree_add_24_21_groupi_n_1343;
  wire csa_tree_add_24_21_groupi_n_1344, csa_tree_add_24_21_groupi_n_1345, csa_tree_add_24_21_groupi_n_1346, csa_tree_add_24_21_groupi_n_1347, csa_tree_add_24_21_groupi_n_1348, csa_tree_add_24_21_groupi_n_1349, csa_tree_add_24_21_groupi_n_1350, csa_tree_add_24_21_groupi_n_1351;
  wire csa_tree_add_24_21_groupi_n_1352, csa_tree_add_24_21_groupi_n_1353, csa_tree_add_24_21_groupi_n_1354, csa_tree_add_24_21_groupi_n_1355, csa_tree_add_24_21_groupi_n_1356, csa_tree_add_24_21_groupi_n_1357, csa_tree_add_24_21_groupi_n_1358, csa_tree_add_24_21_groupi_n_1359;
  wire csa_tree_add_24_21_groupi_n_1360, csa_tree_add_24_21_groupi_n_1361, csa_tree_add_24_21_groupi_n_1362, csa_tree_add_24_21_groupi_n_1363, csa_tree_add_24_21_groupi_n_1364, csa_tree_add_24_21_groupi_n_1365, csa_tree_add_24_21_groupi_n_1366, csa_tree_add_24_21_groupi_n_1367;
  wire csa_tree_add_24_21_groupi_n_1368, csa_tree_add_24_21_groupi_n_1369, csa_tree_add_24_21_groupi_n_1370, csa_tree_add_24_21_groupi_n_1371, csa_tree_add_24_21_groupi_n_1372, csa_tree_add_24_21_groupi_n_1373, csa_tree_add_24_21_groupi_n_1374, csa_tree_add_24_21_groupi_n_1375;
  wire csa_tree_add_24_21_groupi_n_1376, csa_tree_add_24_21_groupi_n_1377, csa_tree_add_24_21_groupi_n_1378, csa_tree_add_24_21_groupi_n_1379, csa_tree_add_24_21_groupi_n_1380, csa_tree_add_24_21_groupi_n_1381, csa_tree_add_24_21_groupi_n_1382, csa_tree_add_24_21_groupi_n_1383;
  wire csa_tree_add_24_21_groupi_n_1384, csa_tree_add_24_21_groupi_n_1385, csa_tree_add_24_21_groupi_n_1386, csa_tree_add_24_21_groupi_n_1387, csa_tree_add_24_21_groupi_n_1388, csa_tree_add_24_21_groupi_n_1389, csa_tree_add_24_21_groupi_n_1390, csa_tree_add_24_21_groupi_n_1391;
  wire csa_tree_add_24_21_groupi_n_1392, csa_tree_add_24_21_groupi_n_1393, csa_tree_add_24_21_groupi_n_1394, csa_tree_add_24_21_groupi_n_1395, csa_tree_add_24_21_groupi_n_1396, csa_tree_add_24_21_groupi_n_1397, csa_tree_add_24_21_groupi_n_1398, csa_tree_add_24_21_groupi_n_1399;
  wire csa_tree_add_24_21_groupi_n_1400, csa_tree_add_24_21_groupi_n_1401, csa_tree_add_24_21_groupi_n_1402, csa_tree_add_24_21_groupi_n_1403, csa_tree_add_24_21_groupi_n_1404, csa_tree_add_24_21_groupi_n_1405, csa_tree_add_24_21_groupi_n_1406, csa_tree_add_24_21_groupi_n_1407;
  wire csa_tree_add_24_21_groupi_n_1408, csa_tree_add_24_21_groupi_n_1409, csa_tree_add_24_21_groupi_n_1410, csa_tree_add_24_21_groupi_n_1411, csa_tree_add_24_21_groupi_n_1412, csa_tree_add_24_21_groupi_n_1413, csa_tree_add_24_21_groupi_n_1414, csa_tree_add_24_21_groupi_n_1415;
  wire csa_tree_add_24_21_groupi_n_1416, csa_tree_add_24_21_groupi_n_1417, csa_tree_add_24_21_groupi_n_1418, csa_tree_add_24_21_groupi_n_1419, csa_tree_add_24_21_groupi_n_1420, csa_tree_add_24_21_groupi_n_1421, csa_tree_add_24_21_groupi_n_1422, csa_tree_add_24_21_groupi_n_1423;
  wire csa_tree_add_24_21_groupi_n_1424, csa_tree_add_24_21_groupi_n_1425, csa_tree_add_24_21_groupi_n_1426, csa_tree_add_24_21_groupi_n_1427, csa_tree_add_24_21_groupi_n_1428, csa_tree_add_24_21_groupi_n_1429, csa_tree_add_24_21_groupi_n_1430, csa_tree_add_24_21_groupi_n_1431;
  wire csa_tree_add_24_21_groupi_n_1432, csa_tree_add_24_21_groupi_n_1433, csa_tree_add_24_21_groupi_n_1434, csa_tree_add_24_21_groupi_n_1435, csa_tree_add_24_21_groupi_n_1436, csa_tree_add_24_21_groupi_n_1437, csa_tree_add_24_21_groupi_n_1438, csa_tree_add_24_21_groupi_n_1439;
  wire csa_tree_add_24_21_groupi_n_1440, csa_tree_add_24_21_groupi_n_1441, csa_tree_add_24_21_groupi_n_1442, csa_tree_add_24_21_groupi_n_1443, csa_tree_add_24_21_groupi_n_1444, csa_tree_add_24_21_groupi_n_1445, csa_tree_add_24_21_groupi_n_1446, csa_tree_add_24_21_groupi_n_1447;
  wire csa_tree_add_24_21_groupi_n_1448, csa_tree_add_24_21_groupi_n_1449, csa_tree_add_24_21_groupi_n_1450, csa_tree_add_24_21_groupi_n_1451, csa_tree_add_24_21_groupi_n_1452, csa_tree_add_24_21_groupi_n_1453, csa_tree_add_24_21_groupi_n_1454, csa_tree_add_24_21_groupi_n_1455;
  wire csa_tree_add_24_21_groupi_n_1456, csa_tree_add_24_21_groupi_n_1457, csa_tree_add_24_21_groupi_n_1458, csa_tree_add_24_21_groupi_n_1459, csa_tree_add_24_21_groupi_n_1460, csa_tree_add_24_21_groupi_n_1461, csa_tree_add_24_21_groupi_n_1462, csa_tree_add_24_21_groupi_n_1463;
  wire csa_tree_add_24_21_groupi_n_1464, csa_tree_add_24_21_groupi_n_1465, csa_tree_add_24_21_groupi_n_1466, csa_tree_add_24_21_groupi_n_1467, csa_tree_add_24_21_groupi_n_1468, csa_tree_add_24_21_groupi_n_1469, csa_tree_add_24_21_groupi_n_1470, csa_tree_add_24_21_groupi_n_1471;
  wire csa_tree_add_24_21_groupi_n_1472, csa_tree_add_24_21_groupi_n_1473, csa_tree_add_24_21_groupi_n_1474, csa_tree_add_24_21_groupi_n_1475, csa_tree_add_24_21_groupi_n_1476, csa_tree_add_24_21_groupi_n_1477, csa_tree_add_24_21_groupi_n_1478, csa_tree_add_24_21_groupi_n_1479;
  wire csa_tree_add_24_21_groupi_n_1480, csa_tree_add_24_21_groupi_n_1481, csa_tree_add_24_21_groupi_n_1482, csa_tree_add_24_21_groupi_n_1483, csa_tree_add_24_21_groupi_n_1484, csa_tree_add_24_21_groupi_n_1485, csa_tree_add_24_21_groupi_n_1486, csa_tree_add_24_21_groupi_n_1487;
  wire csa_tree_add_24_21_groupi_n_1488, csa_tree_add_24_21_groupi_n_1489, csa_tree_add_24_21_groupi_n_1490, csa_tree_add_24_21_groupi_n_1491, csa_tree_add_24_21_groupi_n_1492, csa_tree_add_24_21_groupi_n_1493, csa_tree_add_24_21_groupi_n_1494, csa_tree_add_24_21_groupi_n_1495;
  wire csa_tree_add_24_21_groupi_n_1496, csa_tree_add_24_21_groupi_n_1497, csa_tree_add_24_21_groupi_n_1498, csa_tree_add_24_21_groupi_n_1499, csa_tree_add_24_21_groupi_n_1500, csa_tree_add_24_21_groupi_n_1501, csa_tree_add_24_21_groupi_n_1502, csa_tree_add_24_21_groupi_n_1503;
  wire csa_tree_add_24_21_groupi_n_1504, csa_tree_add_24_21_groupi_n_1505, csa_tree_add_24_21_groupi_n_1506, csa_tree_add_24_21_groupi_n_1507, csa_tree_add_24_21_groupi_n_1508, csa_tree_add_24_21_groupi_n_1509, csa_tree_add_24_21_groupi_n_1510, csa_tree_add_24_21_groupi_n_1511;
  wire csa_tree_add_24_21_groupi_n_1512, csa_tree_add_24_21_groupi_n_1513, csa_tree_add_24_21_groupi_n_1514, csa_tree_add_24_21_groupi_n_1515, csa_tree_add_24_21_groupi_n_1516, csa_tree_add_24_21_groupi_n_1517, csa_tree_add_24_21_groupi_n_1518, csa_tree_add_24_21_groupi_n_1519;
  wire csa_tree_add_24_21_groupi_n_1520, csa_tree_add_24_21_groupi_n_1521, csa_tree_add_24_21_groupi_n_1522, csa_tree_add_24_21_groupi_n_1523, csa_tree_add_24_21_groupi_n_1524, csa_tree_add_24_21_groupi_n_1525, csa_tree_add_24_21_groupi_n_1526, csa_tree_add_24_21_groupi_n_1527;
  wire csa_tree_add_24_21_groupi_n_1528, csa_tree_add_24_21_groupi_n_1529, csa_tree_add_24_21_groupi_n_1530, csa_tree_add_24_21_groupi_n_1531, csa_tree_add_24_21_groupi_n_1532, csa_tree_add_24_21_groupi_n_1533, csa_tree_add_24_21_groupi_n_1534, csa_tree_add_24_21_groupi_n_1535;
  wire csa_tree_add_24_21_groupi_n_1536, csa_tree_add_24_21_groupi_n_1537, csa_tree_add_24_21_groupi_n_1538, csa_tree_add_24_21_groupi_n_1539, csa_tree_add_24_21_groupi_n_1540, csa_tree_add_24_21_groupi_n_1541, csa_tree_add_24_21_groupi_n_1542, csa_tree_add_24_21_groupi_n_1543;
  wire csa_tree_add_24_21_groupi_n_1544, csa_tree_add_24_21_groupi_n_1545, csa_tree_add_24_21_groupi_n_1546, csa_tree_add_24_21_groupi_n_1547, csa_tree_add_24_21_groupi_n_1548, csa_tree_add_24_21_groupi_n_1549, csa_tree_add_24_21_groupi_n_1550, csa_tree_add_24_21_groupi_n_1551;
  wire csa_tree_add_24_21_groupi_n_1552, csa_tree_add_24_21_groupi_n_1553, csa_tree_add_24_21_groupi_n_1554, csa_tree_add_24_21_groupi_n_1555, csa_tree_add_24_21_groupi_n_1556, csa_tree_add_24_21_groupi_n_1557, csa_tree_add_24_21_groupi_n_1558, csa_tree_add_24_21_groupi_n_1559;
  wire csa_tree_add_24_21_groupi_n_1560, csa_tree_add_24_21_groupi_n_1561, csa_tree_add_24_21_groupi_n_1562, csa_tree_add_24_21_groupi_n_1563, csa_tree_add_24_21_groupi_n_1564, csa_tree_add_24_21_groupi_n_1565, csa_tree_add_24_21_groupi_n_1566, csa_tree_add_24_21_groupi_n_1567;
  wire csa_tree_add_24_21_groupi_n_1568, csa_tree_add_24_21_groupi_n_1569, csa_tree_add_24_21_groupi_n_1570, csa_tree_add_24_21_groupi_n_1571, csa_tree_add_24_21_groupi_n_1572, csa_tree_add_24_21_groupi_n_1573, csa_tree_add_24_21_groupi_n_1574, csa_tree_add_24_21_groupi_n_1575;
  wire csa_tree_add_24_21_groupi_n_1576, csa_tree_add_24_21_groupi_n_1577, csa_tree_add_24_21_groupi_n_1578, csa_tree_add_24_21_groupi_n_1579, csa_tree_add_24_21_groupi_n_1580, csa_tree_add_24_21_groupi_n_1581, csa_tree_add_24_21_groupi_n_1582, csa_tree_add_24_21_groupi_n_1583;
  wire csa_tree_add_24_21_groupi_n_1584, csa_tree_add_24_21_groupi_n_1585, csa_tree_add_24_21_groupi_n_1586, csa_tree_add_24_21_groupi_n_1587, csa_tree_add_24_21_groupi_n_1588, csa_tree_add_24_21_groupi_n_1589, csa_tree_add_24_21_groupi_n_1590, csa_tree_add_24_21_groupi_n_1591;
  wire csa_tree_add_24_21_groupi_n_1592, csa_tree_add_24_21_groupi_n_1593, csa_tree_add_24_21_groupi_n_1594, csa_tree_add_24_21_groupi_n_1595, csa_tree_add_24_21_groupi_n_1596, csa_tree_add_24_21_groupi_n_1597, csa_tree_add_24_21_groupi_n_1598, csa_tree_add_24_21_groupi_n_1599;
  wire csa_tree_add_24_21_groupi_n_1600, csa_tree_add_24_21_groupi_n_1601, csa_tree_add_24_21_groupi_n_1602, csa_tree_add_24_21_groupi_n_1603, csa_tree_add_24_21_groupi_n_1604, csa_tree_add_24_21_groupi_n_1605, csa_tree_add_24_21_groupi_n_1606, csa_tree_add_24_21_groupi_n_1607;
  wire csa_tree_add_24_21_groupi_n_1608, csa_tree_add_24_21_groupi_n_1609, csa_tree_add_24_21_groupi_n_1610, csa_tree_add_24_21_groupi_n_1611, csa_tree_add_24_21_groupi_n_1612, csa_tree_add_24_21_groupi_n_1613, csa_tree_add_24_21_groupi_n_1614, csa_tree_add_24_21_groupi_n_1615;
  wire csa_tree_add_24_21_groupi_n_1616, csa_tree_add_24_21_groupi_n_1617, csa_tree_add_24_21_groupi_n_1618, csa_tree_add_24_21_groupi_n_1619, csa_tree_add_24_21_groupi_n_1620, csa_tree_add_24_21_groupi_n_1621, csa_tree_add_24_21_groupi_n_1622, csa_tree_add_24_21_groupi_n_1623;
  wire csa_tree_add_24_21_groupi_n_1624, csa_tree_add_24_21_groupi_n_1625, csa_tree_add_24_21_groupi_n_1626, csa_tree_add_24_21_groupi_n_1627, csa_tree_add_24_21_groupi_n_1628, csa_tree_add_24_21_groupi_n_1629, csa_tree_add_24_21_groupi_n_1630, csa_tree_add_24_21_groupi_n_1631;
  wire csa_tree_add_24_21_groupi_n_1632, csa_tree_add_24_21_groupi_n_1633, csa_tree_add_24_21_groupi_n_1634, csa_tree_add_24_21_groupi_n_1635, csa_tree_add_24_21_groupi_n_1636, csa_tree_add_24_21_groupi_n_1637, csa_tree_add_24_21_groupi_n_1638, csa_tree_add_24_21_groupi_n_1639;
  wire csa_tree_add_24_21_groupi_n_1640, csa_tree_add_24_21_groupi_n_1641, csa_tree_add_24_21_groupi_n_1642, csa_tree_add_24_21_groupi_n_1643, csa_tree_add_24_21_groupi_n_1644, csa_tree_add_24_21_groupi_n_1645, csa_tree_add_24_21_groupi_n_1646, csa_tree_add_24_21_groupi_n_1647;
  wire csa_tree_add_24_21_groupi_n_1648, csa_tree_add_24_21_groupi_n_1649, csa_tree_add_24_21_groupi_n_1650, csa_tree_add_24_21_groupi_n_1651, csa_tree_add_24_21_groupi_n_1652, csa_tree_add_24_21_groupi_n_1653, csa_tree_add_24_21_groupi_n_1654, csa_tree_add_24_21_groupi_n_1655;
  wire csa_tree_add_24_21_groupi_n_1656, csa_tree_add_24_21_groupi_n_1657, csa_tree_add_24_21_groupi_n_1658, csa_tree_add_24_21_groupi_n_1659, csa_tree_add_24_21_groupi_n_1660, csa_tree_add_24_21_groupi_n_1661, csa_tree_add_24_21_groupi_n_1662, csa_tree_add_24_21_groupi_n_1663;
  wire csa_tree_add_24_21_groupi_n_1664, csa_tree_add_24_21_groupi_n_1665, csa_tree_add_24_21_groupi_n_1666, csa_tree_add_24_21_groupi_n_1667, csa_tree_add_24_21_groupi_n_1668, csa_tree_add_24_21_groupi_n_1669, csa_tree_add_24_21_groupi_n_1670, csa_tree_add_24_21_groupi_n_1671;
  wire csa_tree_add_24_21_groupi_n_1672, csa_tree_add_24_21_groupi_n_1673, csa_tree_add_24_21_groupi_n_1674, csa_tree_add_24_21_groupi_n_1675, csa_tree_add_24_21_groupi_n_1676, csa_tree_add_24_21_groupi_n_1677, csa_tree_add_24_21_groupi_n_1678, csa_tree_add_24_21_groupi_n_1679;
  wire csa_tree_add_24_21_groupi_n_1680, csa_tree_add_24_21_groupi_n_1681, csa_tree_add_24_21_groupi_n_1682, csa_tree_add_24_21_groupi_n_1683, csa_tree_add_24_21_groupi_n_1684, csa_tree_add_24_21_groupi_n_1685, csa_tree_add_24_21_groupi_n_1686, csa_tree_add_24_21_groupi_n_1687;
  wire csa_tree_add_24_21_groupi_n_1688, csa_tree_add_24_21_groupi_n_1689, csa_tree_add_24_21_groupi_n_1690, csa_tree_add_24_21_groupi_n_1691, csa_tree_add_24_21_groupi_n_1692, csa_tree_add_24_21_groupi_n_1693, csa_tree_add_24_21_groupi_n_1694, csa_tree_add_24_21_groupi_n_1695;
  wire csa_tree_add_24_21_groupi_n_1696, csa_tree_add_24_21_groupi_n_1697, csa_tree_add_24_21_groupi_n_1698, csa_tree_add_24_21_groupi_n_1699, csa_tree_add_24_21_groupi_n_1700, csa_tree_add_24_21_groupi_n_1701, csa_tree_add_24_21_groupi_n_1702, csa_tree_add_24_21_groupi_n_1703;
  wire csa_tree_add_24_21_groupi_n_1704, csa_tree_add_24_21_groupi_n_1705, csa_tree_add_24_21_groupi_n_1706, csa_tree_add_24_21_groupi_n_1707, csa_tree_add_24_21_groupi_n_1708, csa_tree_add_24_21_groupi_n_1709, csa_tree_add_24_21_groupi_n_1710, csa_tree_add_24_21_groupi_n_1711;
  wire csa_tree_add_24_21_groupi_n_1712, csa_tree_add_24_21_groupi_n_1713, csa_tree_add_24_21_groupi_n_1714, csa_tree_add_24_21_groupi_n_1715, csa_tree_add_24_21_groupi_n_1716, csa_tree_add_24_21_groupi_n_1717, csa_tree_add_24_21_groupi_n_1718, csa_tree_add_24_21_groupi_n_1719;
  wire csa_tree_add_24_21_groupi_n_1720, csa_tree_add_24_21_groupi_n_1721, csa_tree_add_24_21_groupi_n_1722, csa_tree_add_24_21_groupi_n_1723, csa_tree_add_24_21_groupi_n_1724, csa_tree_add_24_21_groupi_n_1725, csa_tree_add_24_21_groupi_n_1726, csa_tree_add_24_21_groupi_n_1727;
  wire csa_tree_add_24_21_groupi_n_1728, csa_tree_add_24_21_groupi_n_1729, csa_tree_add_24_21_groupi_n_1730, csa_tree_add_24_21_groupi_n_1731, csa_tree_add_24_21_groupi_n_1732, csa_tree_add_24_21_groupi_n_1733, csa_tree_add_24_21_groupi_n_1734, csa_tree_add_24_21_groupi_n_1735;
  wire csa_tree_add_24_21_groupi_n_1736, csa_tree_add_24_21_groupi_n_1737, csa_tree_add_24_21_groupi_n_1738, csa_tree_add_24_21_groupi_n_1739, csa_tree_add_24_21_groupi_n_1740, csa_tree_add_24_21_groupi_n_1741, csa_tree_add_24_21_groupi_n_1742, csa_tree_add_24_21_groupi_n_1743;
  wire csa_tree_add_24_21_groupi_n_1744, csa_tree_add_24_21_groupi_n_1745, csa_tree_add_24_21_groupi_n_1746, csa_tree_add_24_21_groupi_n_1747, csa_tree_add_24_21_groupi_n_1748, csa_tree_add_24_21_groupi_n_1749, csa_tree_add_24_21_groupi_n_1750, csa_tree_add_24_21_groupi_n_1751;
  wire csa_tree_add_24_21_groupi_n_1752, csa_tree_add_24_21_groupi_n_1753, csa_tree_add_24_21_groupi_n_1754, csa_tree_add_24_21_groupi_n_1755, csa_tree_add_24_21_groupi_n_1756, csa_tree_add_24_21_groupi_n_1757, csa_tree_add_24_21_groupi_n_1758, csa_tree_add_24_21_groupi_n_1759;
  wire csa_tree_add_24_21_groupi_n_1760, csa_tree_add_24_21_groupi_n_1761, csa_tree_add_24_21_groupi_n_1762, csa_tree_add_24_21_groupi_n_1763, csa_tree_add_24_21_groupi_n_1764, csa_tree_add_24_21_groupi_n_1765, csa_tree_add_24_21_groupi_n_1766, csa_tree_add_24_21_groupi_n_1767;
  wire csa_tree_add_24_21_groupi_n_1768, csa_tree_add_24_21_groupi_n_1769, csa_tree_add_24_21_groupi_n_1770, csa_tree_add_24_21_groupi_n_1771, csa_tree_add_24_21_groupi_n_1772, csa_tree_add_24_21_groupi_n_1773, csa_tree_add_24_21_groupi_n_1774, csa_tree_add_24_21_groupi_n_1775;
  wire csa_tree_add_24_21_groupi_n_1776, csa_tree_add_24_21_groupi_n_1777, csa_tree_add_24_21_groupi_n_1778, csa_tree_add_24_21_groupi_n_1779, csa_tree_add_24_21_groupi_n_1780, csa_tree_add_24_21_groupi_n_1781, csa_tree_add_24_21_groupi_n_1782, csa_tree_add_24_21_groupi_n_1783;
  wire csa_tree_add_24_21_groupi_n_1784, csa_tree_add_24_21_groupi_n_1785, csa_tree_add_24_21_groupi_n_1786, csa_tree_add_24_21_groupi_n_1787, csa_tree_add_24_21_groupi_n_1788, csa_tree_add_24_21_groupi_n_1789, csa_tree_add_24_21_groupi_n_1790, csa_tree_add_24_21_groupi_n_1791;
  wire csa_tree_add_24_21_groupi_n_1792, csa_tree_add_24_21_groupi_n_1793, csa_tree_add_24_21_groupi_n_1794, csa_tree_add_24_21_groupi_n_1795, csa_tree_add_24_21_groupi_n_1796, csa_tree_add_24_21_groupi_n_1797, csa_tree_add_24_21_groupi_n_1798, csa_tree_add_24_21_groupi_n_1799;
  wire csa_tree_add_24_21_groupi_n_1800, csa_tree_add_24_21_groupi_n_1801, csa_tree_add_24_21_groupi_n_1802, csa_tree_add_24_21_groupi_n_1803, csa_tree_add_24_21_groupi_n_1804, csa_tree_add_24_21_groupi_n_1805, csa_tree_add_24_21_groupi_n_1806, csa_tree_add_24_21_groupi_n_1807;
  wire csa_tree_add_24_21_groupi_n_1808, csa_tree_add_24_21_groupi_n_1809, csa_tree_add_24_21_groupi_n_1810, csa_tree_add_24_21_groupi_n_1811, csa_tree_add_24_21_groupi_n_1812, csa_tree_add_24_21_groupi_n_1813, csa_tree_add_24_21_groupi_n_1814, csa_tree_add_24_21_groupi_n_1815;
  wire csa_tree_add_24_21_groupi_n_1816, csa_tree_add_24_21_groupi_n_1817, csa_tree_add_24_21_groupi_n_1818, csa_tree_add_24_21_groupi_n_1819, csa_tree_add_24_21_groupi_n_1820, csa_tree_add_24_21_groupi_n_1821, csa_tree_add_24_21_groupi_n_1822, csa_tree_add_24_21_groupi_n_1823;
  wire csa_tree_add_24_21_groupi_n_1824, csa_tree_add_24_21_groupi_n_1825, csa_tree_add_24_21_groupi_n_1826, csa_tree_add_24_21_groupi_n_1827, csa_tree_add_24_21_groupi_n_1828, csa_tree_add_24_21_groupi_n_1829, csa_tree_add_24_21_groupi_n_1830, csa_tree_add_24_21_groupi_n_1831;
  wire csa_tree_add_24_21_groupi_n_1832, csa_tree_add_24_21_groupi_n_1833, csa_tree_add_24_21_groupi_n_1834, csa_tree_add_24_21_groupi_n_1835, csa_tree_add_24_21_groupi_n_1836, csa_tree_add_24_21_groupi_n_1837, csa_tree_add_24_21_groupi_n_1838, csa_tree_add_24_21_groupi_n_1839;
  wire csa_tree_add_24_21_groupi_n_1840, csa_tree_add_24_21_groupi_n_1841, csa_tree_add_24_21_groupi_n_1842, csa_tree_add_24_21_groupi_n_1843, csa_tree_add_24_21_groupi_n_1844, csa_tree_add_24_21_groupi_n_1845, csa_tree_add_24_21_groupi_n_1846, csa_tree_add_24_21_groupi_n_1847;
  wire csa_tree_add_24_21_groupi_n_1848, csa_tree_add_24_21_groupi_n_1849, csa_tree_add_24_21_groupi_n_1850, csa_tree_add_24_21_groupi_n_1851, csa_tree_add_24_21_groupi_n_1852, csa_tree_add_24_21_groupi_n_1853, csa_tree_add_24_21_groupi_n_1854, csa_tree_add_24_21_groupi_n_1855;
  wire csa_tree_add_24_21_groupi_n_1856, csa_tree_add_24_21_groupi_n_1857, csa_tree_add_24_21_groupi_n_1858, csa_tree_add_24_21_groupi_n_1859, csa_tree_add_24_21_groupi_n_1860, csa_tree_add_24_21_groupi_n_1861, csa_tree_add_24_21_groupi_n_1862, csa_tree_add_24_21_groupi_n_1863;
  wire csa_tree_add_24_21_groupi_n_1864, csa_tree_add_24_21_groupi_n_1865, csa_tree_add_24_21_groupi_n_1866, csa_tree_add_24_21_groupi_n_1867, csa_tree_add_24_21_groupi_n_1868, csa_tree_add_24_21_groupi_n_1869, csa_tree_add_24_21_groupi_n_1870, csa_tree_add_24_21_groupi_n_1871;
  wire csa_tree_add_24_21_groupi_n_1872, csa_tree_add_24_21_groupi_n_1873, csa_tree_add_24_21_groupi_n_1874, csa_tree_add_24_21_groupi_n_1875, csa_tree_add_24_21_groupi_n_1876, csa_tree_add_24_21_groupi_n_1877, csa_tree_add_24_21_groupi_n_1878, csa_tree_add_24_21_groupi_n_1879;
  wire csa_tree_add_24_21_groupi_n_1880, csa_tree_add_24_21_groupi_n_1881, csa_tree_add_24_21_groupi_n_1882, csa_tree_add_24_21_groupi_n_1883, csa_tree_add_24_21_groupi_n_1884, csa_tree_add_24_21_groupi_n_1885, csa_tree_add_24_21_groupi_n_1886, csa_tree_add_24_21_groupi_n_1887;
  wire csa_tree_add_24_21_groupi_n_1888, csa_tree_add_24_21_groupi_n_1889, csa_tree_add_24_21_groupi_n_1890, csa_tree_add_24_21_groupi_n_1891, csa_tree_add_24_21_groupi_n_1892, csa_tree_add_24_21_groupi_n_1893, csa_tree_add_24_21_groupi_n_1894, csa_tree_add_24_21_groupi_n_1895;
  wire csa_tree_add_24_21_groupi_n_1896, csa_tree_add_24_21_groupi_n_1897, csa_tree_add_24_21_groupi_n_1898, csa_tree_add_24_21_groupi_n_1899, csa_tree_add_24_21_groupi_n_1900, csa_tree_add_24_21_groupi_n_1901, csa_tree_add_24_21_groupi_n_1902, csa_tree_add_24_21_groupi_n_1903;
  wire csa_tree_add_24_21_groupi_n_1904, csa_tree_add_24_21_groupi_n_1905, csa_tree_add_24_21_groupi_n_1906, csa_tree_add_24_21_groupi_n_1907, csa_tree_add_24_21_groupi_n_1908, csa_tree_add_24_21_groupi_n_1909, csa_tree_add_24_21_groupi_n_1910, csa_tree_add_24_21_groupi_n_1911;
  wire csa_tree_add_24_21_groupi_n_1912, csa_tree_add_24_21_groupi_n_1913, csa_tree_add_24_21_groupi_n_1914, csa_tree_add_24_21_groupi_n_1915, csa_tree_add_24_21_groupi_n_1916, csa_tree_add_24_21_groupi_n_1917, csa_tree_add_24_21_groupi_n_1918, csa_tree_add_24_21_groupi_n_1919;
  wire csa_tree_add_24_21_groupi_n_1920, csa_tree_add_24_21_groupi_n_1921, csa_tree_add_24_21_groupi_n_1922, csa_tree_add_24_21_groupi_n_1923, csa_tree_add_24_21_groupi_n_1924, csa_tree_add_24_21_groupi_n_1925, csa_tree_add_24_21_groupi_n_1926, csa_tree_add_24_21_groupi_n_1927;
  wire csa_tree_add_24_21_groupi_n_1928, csa_tree_add_24_21_groupi_n_1929, csa_tree_add_24_21_groupi_n_1930, csa_tree_add_24_21_groupi_n_1931, csa_tree_add_24_21_groupi_n_1932, csa_tree_add_24_21_groupi_n_1933, csa_tree_add_24_21_groupi_n_1934, csa_tree_add_24_21_groupi_n_1935;
  wire csa_tree_add_24_21_groupi_n_1936, csa_tree_add_24_21_groupi_n_1937, csa_tree_add_24_21_groupi_n_1938, csa_tree_add_24_21_groupi_n_1939, csa_tree_add_24_21_groupi_n_1940, csa_tree_add_24_21_groupi_n_1941, csa_tree_add_24_21_groupi_n_1942, csa_tree_add_24_21_groupi_n_1943;
  wire csa_tree_add_24_21_groupi_n_1944, csa_tree_add_24_21_groupi_n_1945, csa_tree_add_24_21_groupi_n_1946, csa_tree_add_24_21_groupi_n_1947, csa_tree_add_24_21_groupi_n_1948, csa_tree_add_24_21_groupi_n_1949, csa_tree_add_24_21_groupi_n_1950, csa_tree_add_24_21_groupi_n_1951;
  wire csa_tree_add_24_21_groupi_n_1952, csa_tree_add_24_21_groupi_n_1953, csa_tree_add_24_21_groupi_n_1954, csa_tree_add_24_21_groupi_n_1955, csa_tree_add_24_21_groupi_n_1956, csa_tree_add_24_21_groupi_n_1957, csa_tree_add_24_21_groupi_n_1958, csa_tree_add_24_21_groupi_n_1959;
  wire csa_tree_add_24_21_groupi_n_1960, csa_tree_add_24_21_groupi_n_1961, csa_tree_add_24_21_groupi_n_1962, csa_tree_add_24_21_groupi_n_1963, csa_tree_add_24_21_groupi_n_1964, csa_tree_add_24_21_groupi_n_1965, csa_tree_add_24_21_groupi_n_1966, csa_tree_add_24_21_groupi_n_1967;
  wire csa_tree_add_24_21_groupi_n_1968, csa_tree_add_24_21_groupi_n_1969, csa_tree_add_24_21_groupi_n_1970, csa_tree_add_24_21_groupi_n_1971, csa_tree_add_24_21_groupi_n_1972, csa_tree_add_24_21_groupi_n_1973, csa_tree_add_24_21_groupi_n_1974, csa_tree_add_24_21_groupi_n_1975;
  wire csa_tree_add_24_21_groupi_n_1976, csa_tree_add_24_21_groupi_n_1977, csa_tree_add_24_21_groupi_n_1978, csa_tree_add_24_21_groupi_n_1979, csa_tree_add_24_21_groupi_n_1980, csa_tree_add_24_21_groupi_n_1981, csa_tree_add_24_21_groupi_n_1982, csa_tree_add_24_21_groupi_n_1983;
  wire csa_tree_add_24_21_groupi_n_1984, csa_tree_add_24_21_groupi_n_1985, csa_tree_add_24_21_groupi_n_1986, csa_tree_add_24_21_groupi_n_1987, csa_tree_add_24_21_groupi_n_1988, csa_tree_add_24_21_groupi_n_1989, csa_tree_add_24_21_groupi_n_1990, csa_tree_add_24_21_groupi_n_1991;
  wire csa_tree_add_24_21_groupi_n_1992, csa_tree_add_24_21_groupi_n_1993, csa_tree_add_24_21_groupi_n_1994, csa_tree_add_24_21_groupi_n_1995, csa_tree_add_24_21_groupi_n_1996, csa_tree_add_24_21_groupi_n_1997, csa_tree_add_24_21_groupi_n_1998, csa_tree_add_24_21_groupi_n_1999;
  wire csa_tree_add_24_21_groupi_n_2000, csa_tree_add_24_21_groupi_n_2001, csa_tree_add_24_21_groupi_n_2002, csa_tree_add_24_21_groupi_n_2003, csa_tree_add_24_21_groupi_n_2004, csa_tree_add_24_21_groupi_n_2005, csa_tree_add_24_21_groupi_n_2006, csa_tree_add_24_21_groupi_n_2007;
  wire csa_tree_add_24_21_groupi_n_2008, csa_tree_add_24_21_groupi_n_2009, csa_tree_add_24_21_groupi_n_2010, csa_tree_add_24_21_groupi_n_2011, csa_tree_add_24_21_groupi_n_2012, csa_tree_add_24_21_groupi_n_2013, csa_tree_add_24_21_groupi_n_2014, csa_tree_add_24_21_groupi_n_2015;
  wire csa_tree_add_24_21_groupi_n_2016, csa_tree_add_24_21_groupi_n_2017, csa_tree_add_24_21_groupi_n_2018, csa_tree_add_24_21_groupi_n_2019, csa_tree_add_24_21_groupi_n_2020, csa_tree_add_24_21_groupi_n_2021, csa_tree_add_24_21_groupi_n_2022, csa_tree_add_24_21_groupi_n_2023;
  wire csa_tree_add_24_21_groupi_n_2024, csa_tree_add_24_21_groupi_n_2025, csa_tree_add_24_21_groupi_n_2026, csa_tree_add_24_21_groupi_n_2027, csa_tree_add_26_22_groupi_n_0, csa_tree_add_26_22_groupi_n_1, csa_tree_add_26_22_groupi_n_2, csa_tree_add_26_22_groupi_n_3;
  wire csa_tree_add_26_22_groupi_n_4, csa_tree_add_26_22_groupi_n_5, csa_tree_add_26_22_groupi_n_6, csa_tree_add_26_22_groupi_n_7, csa_tree_add_26_22_groupi_n_8, csa_tree_add_26_22_groupi_n_9, csa_tree_add_26_22_groupi_n_10, csa_tree_add_26_22_groupi_n_11;
  wire csa_tree_add_26_22_groupi_n_12, csa_tree_add_26_22_groupi_n_13, csa_tree_add_26_22_groupi_n_14, csa_tree_add_26_22_groupi_n_15, csa_tree_add_26_22_groupi_n_16, csa_tree_add_26_22_groupi_n_17, csa_tree_add_26_22_groupi_n_18, csa_tree_add_26_22_groupi_n_19;
  wire csa_tree_add_26_22_groupi_n_20, csa_tree_add_26_22_groupi_n_21, csa_tree_add_26_22_groupi_n_22, csa_tree_add_26_22_groupi_n_29, csa_tree_add_26_22_groupi_n_30, csa_tree_add_26_22_groupi_n_31, csa_tree_add_26_22_groupi_n_32, csa_tree_add_26_22_groupi_n_37;
  wire csa_tree_add_26_22_groupi_n_39, csa_tree_add_26_22_groupi_n_40, csa_tree_add_26_22_groupi_n_41, csa_tree_add_26_22_groupi_n_42, csa_tree_add_26_22_groupi_n_43, csa_tree_add_26_22_groupi_n_44, csa_tree_add_26_22_groupi_n_45, csa_tree_add_26_22_groupi_n_46;
  wire csa_tree_add_26_22_groupi_n_47, csa_tree_add_26_22_groupi_n_48, csa_tree_add_26_22_groupi_n_49, csa_tree_add_26_22_groupi_n_50, csa_tree_add_26_22_groupi_n_51, csa_tree_add_26_22_groupi_n_52, csa_tree_add_26_22_groupi_n_53, csa_tree_add_26_22_groupi_n_68;
  wire csa_tree_add_26_22_groupi_n_69, csa_tree_add_26_22_groupi_n_70, csa_tree_add_26_22_groupi_n_71, csa_tree_add_26_22_groupi_n_72, csa_tree_add_26_22_groupi_n_73, csa_tree_add_26_22_groupi_n_74, csa_tree_add_26_22_groupi_n_75, csa_tree_add_26_22_groupi_n_76;
  wire csa_tree_add_26_22_groupi_n_77, csa_tree_add_26_22_groupi_n_78, csa_tree_add_26_22_groupi_n_80, csa_tree_add_26_22_groupi_n_81, csa_tree_add_26_22_groupi_n_83, csa_tree_add_26_22_groupi_n_84, csa_tree_add_26_22_groupi_n_85, csa_tree_add_26_22_groupi_n_87;
  wire csa_tree_add_26_22_groupi_n_88, csa_tree_add_26_22_groupi_n_89, csa_tree_add_26_22_groupi_n_91, csa_tree_add_26_22_groupi_n_93, csa_tree_add_26_22_groupi_n_94, csa_tree_add_26_22_groupi_n_95, csa_tree_add_26_22_groupi_n_96, csa_tree_add_26_22_groupi_n_97;
  wire csa_tree_add_26_22_groupi_n_99, csa_tree_add_26_22_groupi_n_101, csa_tree_add_26_22_groupi_n_102, csa_tree_add_26_22_groupi_n_103, csa_tree_add_26_22_groupi_n_104, csa_tree_add_26_22_groupi_n_105, csa_tree_add_26_22_groupi_n_106, csa_tree_add_26_22_groupi_n_107;
  wire csa_tree_add_26_22_groupi_n_108, csa_tree_add_26_22_groupi_n_109, csa_tree_add_26_22_groupi_n_110, csa_tree_add_26_22_groupi_n_111, csa_tree_add_26_22_groupi_n_112, csa_tree_add_26_22_groupi_n_113, csa_tree_add_26_22_groupi_n_114, csa_tree_add_26_22_groupi_n_115;
  wire csa_tree_add_26_22_groupi_n_116, csa_tree_add_26_22_groupi_n_117, csa_tree_add_26_22_groupi_n_118, csa_tree_add_26_22_groupi_n_120, csa_tree_add_26_22_groupi_n_122, csa_tree_add_26_22_groupi_n_124, csa_tree_add_26_22_groupi_n_126, csa_tree_add_26_22_groupi_n_128;
  wire csa_tree_add_26_22_groupi_n_130, csa_tree_add_26_22_groupi_n_132, csa_tree_add_26_22_groupi_n_133, csa_tree_add_26_22_groupi_n_137, csa_tree_add_26_22_groupi_n_139, csa_tree_add_26_22_groupi_n_141, csa_tree_add_26_22_groupi_n_143, csa_tree_add_26_22_groupi_n_145;
  wire csa_tree_add_26_22_groupi_n_146, csa_tree_add_26_22_groupi_n_147, csa_tree_add_26_22_groupi_n_148, csa_tree_add_26_22_groupi_n_149, csa_tree_add_26_22_groupi_n_150, csa_tree_add_26_22_groupi_n_151, csa_tree_add_26_22_groupi_n_152, csa_tree_add_26_22_groupi_n_153;
  wire csa_tree_add_26_22_groupi_n_154, csa_tree_add_26_22_groupi_n_155, csa_tree_add_26_22_groupi_n_156, csa_tree_add_26_22_groupi_n_157, csa_tree_add_26_22_groupi_n_158, csa_tree_add_26_22_groupi_n_160, csa_tree_add_26_22_groupi_n_161, csa_tree_add_26_22_groupi_n_163;
  wire csa_tree_add_26_22_groupi_n_164, csa_tree_add_26_22_groupi_n_166, csa_tree_add_26_22_groupi_n_167, csa_tree_add_26_22_groupi_n_168, csa_tree_add_26_22_groupi_n_170, csa_tree_add_26_22_groupi_n_171, csa_tree_add_26_22_groupi_n_172, csa_tree_add_26_22_groupi_n_173;
  wire csa_tree_add_26_22_groupi_n_174, csa_tree_add_26_22_groupi_n_175, csa_tree_add_26_22_groupi_n_176, csa_tree_add_26_22_groupi_n_177, csa_tree_add_26_22_groupi_n_178, csa_tree_add_26_22_groupi_n_179, csa_tree_add_26_22_groupi_n_126, csa_tree_add_26_22_groupi_n_93;
  wire csa_tree_add_26_22_groupi_n_122, csa_tree_add_26_22_groupi_n_101, csa_tree_add_26_22_groupi_n_124, csa_tree_add_26_22_groupi_n_87, csa_tree_add_26_22_groupi_n_128, csa_tree_add_26_22_groupi_n_120, csa_tree_add_26_22_groupi_n_99, csa_tree_add_26_22_groupi_n_83;
  wire csa_tree_add_26_22_groupi_n_130, csa_tree_add_26_22_groupi_n_91, csa_tree_add_26_22_groupi_n_192, csa_tree_add_26_22_groupi_n_193, csa_tree_add_26_22_groupi_n_194, csa_tree_add_26_22_groupi_n_195, csa_tree_add_26_22_groupi_n_197, csa_tree_add_26_22_groupi_n_198;
  wire csa_tree_add_26_22_groupi_n_199, csa_tree_add_26_22_groupi_n_200, csa_tree_add_26_22_groupi_n_201, csa_tree_add_26_22_groupi_n_202, csa_tree_add_26_22_groupi_n_203, csa_tree_add_26_22_groupi_n_204, csa_tree_add_26_22_groupi_n_205, csa_tree_add_26_22_groupi_n_206;
  wire csa_tree_add_26_22_groupi_n_207, csa_tree_add_26_22_groupi_n_208, csa_tree_add_26_22_groupi_n_209, csa_tree_add_26_22_groupi_n_210, csa_tree_add_26_22_groupi_n_211, csa_tree_add_26_22_groupi_n_212, csa_tree_add_26_22_groupi_n_213, csa_tree_add_26_22_groupi_n_214;
  wire csa_tree_add_26_22_groupi_n_215, csa_tree_add_26_22_groupi_n_216, csa_tree_add_26_22_groupi_n_217, csa_tree_add_26_22_groupi_n_218, csa_tree_add_26_22_groupi_n_219, csa_tree_add_26_22_groupi_n_220, csa_tree_add_26_22_groupi_n_221, csa_tree_add_26_22_groupi_n_222;
  wire csa_tree_add_26_22_groupi_n_223, csa_tree_add_26_22_groupi_n_224, csa_tree_add_26_22_groupi_n_225, csa_tree_add_26_22_groupi_n_226, csa_tree_add_26_22_groupi_n_227, csa_tree_add_26_22_groupi_n_228, csa_tree_add_26_22_groupi_n_229, csa_tree_add_26_22_groupi_n_230;
  wire csa_tree_add_26_22_groupi_n_231, csa_tree_add_26_22_groupi_n_232, csa_tree_add_26_22_groupi_n_233, csa_tree_add_26_22_groupi_n_234, csa_tree_add_26_22_groupi_n_235, csa_tree_add_26_22_groupi_n_236, csa_tree_add_26_22_groupi_n_237, csa_tree_add_26_22_groupi_n_238;
  wire csa_tree_add_26_22_groupi_n_239, csa_tree_add_26_22_groupi_n_240, csa_tree_add_26_22_groupi_n_241, csa_tree_add_26_22_groupi_n_242, csa_tree_add_26_22_groupi_n_243, csa_tree_add_26_22_groupi_n_244, csa_tree_add_26_22_groupi_n_245, csa_tree_add_26_22_groupi_n_246;
  wire csa_tree_add_26_22_groupi_n_247, csa_tree_add_26_22_groupi_n_248, csa_tree_add_26_22_groupi_n_250, csa_tree_add_26_22_groupi_n_251, csa_tree_add_26_22_groupi_n_252, csa_tree_add_26_22_groupi_n_253, csa_tree_add_26_22_groupi_n_254, csa_tree_add_26_22_groupi_n_255;
  wire csa_tree_add_26_22_groupi_n_256, csa_tree_add_26_22_groupi_n_257, csa_tree_add_26_22_groupi_n_258, csa_tree_add_26_22_groupi_n_260, csa_tree_add_26_22_groupi_n_262, csa_tree_add_26_22_groupi_n_263, csa_tree_add_26_22_groupi_n_265, csa_tree_add_26_22_groupi_n_266;
  wire csa_tree_add_26_22_groupi_n_268, csa_tree_add_26_22_groupi_n_269, csa_tree_add_26_22_groupi_n_271, csa_tree_add_26_22_groupi_n_272, csa_tree_add_26_22_groupi_n_274, csa_tree_add_26_22_groupi_n_275, csa_tree_add_26_22_groupi_n_277, csa_tree_add_26_22_groupi_n_278;
  wire csa_tree_add_26_22_groupi_n_280, csa_tree_add_26_22_groupi_n_281, csa_tree_add_26_22_groupi_n_283, csa_tree_add_26_22_groupi_n_284, csa_tree_add_26_22_groupi_n_286, csa_tree_add_26_22_groupi_n_287, csa_tree_add_26_22_groupi_n_289, csa_tree_add_26_22_groupi_n_290;
  wire csa_tree_add_26_22_groupi_n_292, csa_tree_add_26_22_groupi_n_293, csa_tree_add_26_22_groupi_n_295, csa_tree_add_26_22_groupi_n_296, csa_tree_add_26_22_groupi_n_298, csa_tree_add_26_22_groupi_n_299, csa_tree_add_26_22_groupi_n_301, csa_tree_add_26_22_groupi_n_302;
  wire csa_tree_add_26_22_groupi_n_304, csa_tree_add_26_22_groupi_n_305, csa_tree_add_26_22_groupi_n_307, csa_tree_add_26_22_groupi_n_308, csa_tree_add_26_22_groupi_n_310, csa_tree_add_26_22_groupi_n_311, csa_tree_add_26_22_groupi_n_313, csa_tree_add_26_22_groupi_n_314;
  wire csa_tree_add_26_22_groupi_n_316, csa_tree_add_26_22_groupi_n_317, csa_tree_add_26_22_groupi_n_319, csa_tree_add_26_22_groupi_n_320, csa_tree_add_26_22_groupi_n_322, csa_tree_add_26_22_groupi_n_323, csa_tree_add_26_22_groupi_n_325, csa_tree_add_26_22_groupi_n_326;
  wire csa_tree_add_26_22_groupi_n_328, csa_tree_add_26_22_groupi_n_329, csa_tree_add_26_22_groupi_n_331, csa_tree_add_26_22_groupi_n_332, csa_tree_add_26_22_groupi_n_334, csa_tree_add_26_22_groupi_n_335, csa_tree_add_26_22_groupi_n_337, csa_tree_add_26_22_groupi_n_338;
  wire csa_tree_add_26_22_groupi_n_340, csa_tree_add_26_22_groupi_n_341, csa_tree_add_26_22_groupi_n_343, n_2, n_3, n_4, n_5, n_6;
  wire n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14;
  wire n_15, n_16, n_17, n_18, n_19, n_34, n_35, n_36;
  wire n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44;
  wire n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52;
  wire n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60;
  wire n_61, n_62, n_63, n_64, n_65, n_307, n_308, n_309;
  wire n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317;
  wire n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
  wire n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381;
  wire n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389;
  wire n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397;
  wire n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405;
  wire n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413;
  wire n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421;
  wire n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429;
  wire n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437;
  wire n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445;
  wire n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453;
  wire n_454, n_470, n_471, n_472, n_473, n_474, n_475, n_476;
  wire n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484;
  wire n_485, n_487, n_488, n_489, n_490, n_491, n_492, n_493;
  wire n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501;
  wire n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509;
  wire n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517;
  wire n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_530, n_531, n_532, n_533;
  wire n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541;
  wire n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581;
  wire n_582, n_597, n_598, n_599, n_600, n_601, n_602, n_603;
  wire n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611;
  wire n_612, n_613, n_614, n_615, n_616, n_617, n_618, n_619;
  wire n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627;
  wire n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635;
  wire n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643;
  wire n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651;
  wire n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659;
  wire n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667;
  wire n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675;
  wire n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683;
  wire n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691;
  wire n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699;
  wire n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707;
  wire n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715;
  wire n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723;
  wire n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731;
  wire n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739;
  wire n_740, n_741, n_742, n_747, n_748, n_749, n_750, n_751;
  wire n_752, n_753, n_754, n_755, n_756, n_757, n_758, n_759;
  wire n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767;
  wire n_768, n_769, n_770, n_771, n_772, n_776, n_777, n_778;
  wire n_779, n_780, n_781, n_782, n_783, n_785, n_786, n_788;
  wire n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796;
  wire n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810;
  wire n_811, n_812, n_814, n_815, n_816, n_817, n_818, n_819;
  wire n_820, n_821, n_823, n_825, n_827, n_829, n_830, n_832;
  wire n_833, n_835, n_836, n_840, n_842, n_843, n_847, n_848;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865;
  wire n_866, n_867, n_868, n_869, n_870, n_871, n_874, n_875;
  wire n_877, n_878, n_881, n_882, n_884, n_885, n_888, n_889;
  wire n_892, n_893, n_897;
  buf constbuf_n1(out2[0] ,out1[0]);
  buf constbuf_n2(out2[1] ,out1[1]);
  buf constbuf_n3(out2[2] ,out1[2]);
  buf constbuf_n4(out2[3] ,out1[3]);
  buf constbuf_n5(out2[4] ,out1[4]);
  buf constbuf_n6(out2[5] ,out1[5]);
  not g63(out2[6] ,out1[6]);
  buf g646(n_766 ,in9[29]);
  buf g645(n_765 ,in9[30]);
  buf g644(n_764 ,in9[31]);
  buf g647(n_763 ,in9[28]);
  buf g648(n_762 ,in9[27]);
  buf g649(n_761 ,in9[26]);
  buf g651(n_760 ,in9[24]);
  buf g652(n_759 ,in9[23]);
  buf g653(n_758 ,in9[22]);
  buf g654(n_757 ,in9[21]);
  buf g655(n_756 ,in9[20]);
  buf g656(n_755 ,in9[19]);
  buf g657(n_754 ,in9[18]);
  buf g658(n_753 ,in9[17]);
  buf g659(n_752 ,n_470);
  buf g660(n_751 ,n_471);
  buf g661(n_750 ,n_472);
  buf g662(n_749 ,n_473);
  buf g663(n_748 ,n_474);
  buf g664(n_747 ,n_475);
  buf g665(n_742 ,n_476);
  buf g667(n_741 ,n_478);
  buf g668(n_740 ,n_479);
  buf g669(n_739 ,n_480);
  buf g670(n_738 ,n_481);
  buf g671(n_737 ,n_482);
  buf g672(n_736 ,n_483);
  buf g673(n_735 ,n_484);
  buf g650(n_734 ,in9[25]);
  buf g675(n_733 ,in9[0]);
  buf g666(n_732 ,n_477);
  buf g674(n_731 ,n_485);
  or g1316__2398(n_51 ,n_656 ,n_703);
  or g1317__5107(n_64 ,n_651 ,n_708);
  or g1318__6260(n_60 ,n_655 ,n_718);
  or g1319__4319(n_54 ,n_653 ,n_715);
  or g1320__8428(n_44 ,n_640 ,n_719);
  or g1321__5526(n_43 ,n_654 ,n_717);
  or g1322__6783(n_42 ,n_652 ,n_714);
  or g1323__3680(n_59 ,n_647 ,n_710);
  or g1324__1617(n_53 ,n_649 ,n_712);
  or g1325__2802(n_730 ,n_650 ,n_713);
  or g1326__1705(n_729 ,n_648 ,n_711);
  or g1327__5122(n_728 ,n_646 ,n_709);
  or g1328__8246(n_62 ,n_641 ,n_689);
  or g1329__7098(n_52 ,n_645 ,n_707);
  or g1330__6131(n_727 ,n_644 ,n_706);
  or g1331__1881(n_65 ,n_643 ,n_692);
  or g1332__5115(n_45 ,n_626 ,n_704);
  or g1333__7482(n_58 ,n_638 ,n_701);
  or g1334__4733(n_726 ,n_639 ,n_702);
  or g1335__6161(n_725 ,n_637 ,n_700);
  or g1336__9315(n_50 ,n_636 ,n_699);
  or g1337__9945(n_724 ,n_635 ,n_698);
  or g1338__2883(n_63 ,n_627 ,n_716);
  or g1339__2346(n_61 ,n_631 ,n_694);
  or g1340__1666(n_57 ,n_633 ,n_696);
  or g1341__7410(n_723 ,n_634 ,n_697);
  or g1342__6417(n_48 ,n_632 ,n_695);
  or g1343__5477(n_722 ,n_630 ,n_693);
  or g1344__2398(n_56 ,n_629 ,n_691);
  or g1345__5107(n_721 ,n_628 ,n_690);
  or g1346__6260(n_55 ,n_625 ,n_705);
  or g1347__4319(n_37 ,n_642 ,n_720);
  or g1348__8428(n_720 ,n_454 ,n_688);
  or g1349__5526(n_719 ,n_513 ,n_687);
  or g1350__6783(n_718 ,n_504 ,n_682);
  or g1351__3680(n_717 ,n_508 ,n_685);
  or g1352__1617(n_716 ,n_507 ,n_680);
  or g1353__2802(n_715 ,n_506 ,n_683);
  or g1354__1705(n_714 ,n_550 ,n_684);
  or g1355__5122(n_713 ,n_501 ,n_681);
  or g1356__8246(n_712 ,n_498 ,n_678);
  or g1357__7098(n_711 ,n_497 ,n_679);
  or g1358__6131(n_710 ,n_491 ,n_674);
  or g1359__1881(n_709 ,n_494 ,n_677);
  or g1360__5115(n_708 ,n_437 ,n_664);
  or g1361__7482(n_707 ,n_490 ,n_675);
  or g1362__4733(n_706 ,n_489 ,n_676);
  or g1363__6161(n_705 ,n_514 ,n_686);
  or g1364__9315(n_704 ,n_503 ,n_672);
  or g1365__9945(n_703 ,n_451 ,n_671);
  or g1366__2883(n_702 ,n_450 ,n_657);
  or g1367__2346(n_701 ,n_517 ,n_667);
  or g1368__1666(n_700 ,n_447 ,n_670);
  or g1369__7410(n_699 ,n_445 ,n_669);
  or g1370__6417(n_698 ,n_510 ,n_668);
  or g1371__5477(n_697 ,n_440 ,n_665);
  or g1372__2398(n_696 ,n_436 ,n_662);
  or g1373__5107(n_695 ,n_435 ,n_663);
  or g1374__6260(n_694 ,n_428 ,n_658);
  or g1375__4319(n_693 ,n_431 ,n_661);
  or g1376__8428(n_692 ,n_511 ,n_673);
  or g1377__5526(n_691 ,n_427 ,n_659);
  or g1378__6783(n_690 ,n_426 ,n_660);
  or g1379__3680(n_689 ,n_452 ,n_666);
  nor g1380__1617(n_688 ,n_538 ,n_576);
  nor g1381__2802(n_687 ,n_548 ,n_623);
  nor g1382__1705(n_686 ,n_547 ,n_622);
  nor g1383__5122(n_685 ,n_546 ,n_621);
  nor g1384__8246(n_684 ,n_545 ,n_619);
  nor g1385__7098(n_683 ,n_544 ,n_618);
  nor g1386__6131(n_682 ,n_543 ,n_617);
  nor g1387__1881(n_681 ,n_520 ,n_616);
  nor g1388__5115(n_680 ,n_541 ,n_620);
  nor g1389__7482(n_679 ,n_536 ,n_615);
  nor g1390__4733(n_678 ,n_540 ,n_582);
  nor g1391__6161(n_677 ,n_539 ,n_580);
  nor g1392__9315(n_676 ,n_537 ,n_579);
  nor g1393__9945(n_675 ,n_534 ,n_578);
  nor g1394__2883(n_674 ,n_532 ,n_581);
  nor g1395__2346(n_673 ,n_527 ,n_562);
  nor g1396__1666(n_672 ,n_518 ,n_561);
  nor g1397__7410(n_671 ,n_522 ,n_570);
  nor g1398__6417(n_670 ,n_533 ,n_624);
  nor g1399__5477(n_669 ,n_549 ,n_574);
  nor g1400__2398(n_668 ,n_542 ,n_575);
  nor g1401__5107(n_667 ,n_530 ,n_573);
  nor g1402__6260(n_666 ,n_529 ,n_572);
  nor g1403__4319(n_665 ,n_528 ,n_571);
  nor g1404__8428(n_664 ,n_531 ,n_567);
  nor g1405__5526(n_663 ,n_526 ,n_569);
  nor g1406__6783(n_662 ,n_525 ,n_568);
  nor g1407__3680(n_661 ,n_523 ,n_566);
  nor g1408__1617(n_660 ,n_521 ,n_565);
  nor g1409__2802(n_659 ,n_524 ,n_564);
  nor g1410__1705(n_658 ,n_519 ,n_563);
  nor g1411__5122(n_657 ,n_535 ,n_577);
  and g1412__8246(n_656 ,out1[17] ,n_309);
  and g1413__7098(n_655 ,out1[26] ,n_333);
  and g1414__6131(n_654 ,out1[9] ,n_342);
  and g1415__1881(n_653 ,out1[20] ,n_350);
  and g1416__5115(n_652 ,out1[8] ,n_344);
  and g1417__7482(n_651 ,out1[30] ,n_338);
  and g1418__4733(n_650 ,out1[7] ,n_348);
  and g1419__6161(n_649 ,out1[19] ,n_344);
  and g1420__9315(n_648 ,out1[6] ,n_348);
  and g1421__9945(n_647 ,out1[25] ,n_338);
  and g1422__2883(n_646 ,out1[5] ,n_350);
  and g1423__2346(n_645 ,out1[18] ,n_339);
  and g1424__1666(n_644 ,out1[4] ,n_336);
  and g1425__7410(n_643 ,out1[31] ,n_351);
  and g1426__6417(n_642 ,out1[3] ,n_341);
  and g1427__5477(n_641 ,out1[28] ,n_335);
  and g1428__2398(n_640 ,out1[10] ,n_341);
  and g1429__5107(n_639 ,out1[2] ,n_308);
  and g1430__6260(n_638 ,out1[24] ,n_332);
  and g1431__4319(n_637 ,out1[1] ,n_336);
  and g1432__8428(n_636 ,out1[16] ,n_345);
  and g1433__5526(n_635 ,out1[0] ,n_332);
  and g1434__6783(n_634 ,out1[15] ,n_347);
  and g1435__3680(n_633 ,out1[23] ,n_351);
  and g1436__1617(n_632 ,out1[14] ,n_347);
  and g1437__2802(n_631 ,out1[27] ,n_339);
  and g1438__1705(n_630 ,out1[13] ,n_342);
  and g1439__5122(n_629 ,out1[22] ,n_335);
  and g1440__8246(n_628 ,out1[12] ,n_345);
  and g1441__7098(n_627 ,out1[29] ,n_308);
  and g1442__6131(n_626 ,out1[11] ,n_333);
  and g1443__1881(n_625 ,out1[21] ,n_309);
  or g1444__5115(n_624 ,n_446 ,n_315);
  or g1445__7482(n_623 ,n_512 ,n_330);
  or g1446__4733(n_622 ,n_509 ,n_324);
  or g1447__6161(n_621 ,n_505 ,n_320);
  or g1448__9315(n_620 ,n_493 ,n_353);
  or g1449__9945(n_619 ,n_423 ,n_326);
  or g1450__2883(n_618 ,n_502 ,n_318);
  or g1451__2346(n_617 ,n_499 ,n_353);
  or g1452__1666(n_616 ,n_500 ,n_318);
  or g1453__7410(n_615 ,n_496 ,n_326);
  or g1454__6417(n_582 ,n_495 ,n_320);
  or g1455__5477(n_581 ,n_434 ,n_327);
  or g1456__2398(n_580 ,n_492 ,n_312);
  or g1457__5107(n_579 ,n_488 ,n_321);
  or g1458__6260(n_578 ,n_487 ,n_323);
  or g1459__4319(n_577 ,n_449 ,n_311);
  or g1460__8428(n_576 ,n_453 ,n_323);
  or g1461__5526(n_575 ,n_443 ,n_314);
  or g1462__6783(n_574 ,n_442 ,n_329);
  or g1463__3680(n_573 ,n_441 ,n_312);
  or g1464__1617(n_572 ,n_444 ,n_354);
  or g1465__2802(n_571 ,n_438 ,n_329);
  or g1466__1705(n_570 ,n_448 ,n_317);
  or g1467__5122(n_569 ,n_433 ,n_321);
  or g1468__8246(n_568 ,n_432 ,n_317);
  or g1469__7098(n_567 ,n_430 ,n_327);
  or g1470__6131(n_566 ,n_429 ,n_324);
  or g1471__1881(n_565 ,n_425 ,n_311);
  or g1472__5115(n_564 ,n_424 ,n_354);
  or g1473__7482(n_563 ,n_515 ,n_314);
  or g1474__4733(n_562 ,n_439 ,n_330);
  or g1475__6161(n_561 ,n_516 ,n_315);
  not g1476(n_560 ,n_558);
  not g1477(n_559 ,n_360);
  not g1478(n_557 ,n_360);
  not g1479(n_556 ,n_558);
  not g1480(n_555 ,n_553);
  not g1481(n_554 ,n_358);
  not g1482(n_552 ,n_358);
  not g1483(n_551 ,n_553);
  and g1484__9315(n_550 ,in4 ,out2[8]);
  nor g1485__9945(n_549 ,n_382 ,n_752);
  nor g1486__2883(n_548 ,n_377 ,n_742);
  nor g1487__2346(n_547 ,n_385 ,n_757);
  nor g1488__1666(n_546 ,n_368 ,n_732);
  nor g1489__7410(n_545 ,n_365 ,n_741);
  nor g1490__6417(n_544 ,n_368 ,n_756);
  nor g1491__5477(n_543 ,n_370 ,n_761);
  nor g1492__2398(n_542 ,n_379 ,n_733);
  nor g1493__5107(n_541 ,n_367 ,n_766);
  nor g1494__6260(n_540 ,n_374 ,n_755);
  nor g1495__4319(n_539 ,n_383 ,n_738);
  nor g1496__8428(n_538 ,n_374 ,n_736);
  nor g1497__5526(n_537 ,n_373 ,n_737);
  nor g1498__6783(n_536 ,n_371 ,n_739);
  nor g1499__3680(n_535 ,n_380 ,n_735);
  nor g1500__1617(n_534 ,n_373 ,n_754);
  nor g1501__2802(n_533 ,n_376 ,n_731);
  nor g1502__1705(n_532 ,n_386 ,n_734);
  nor g1503__5122(n_531 ,n_367 ,n_765);
  nor g1504__8246(n_530 ,n_382 ,n_760);
  nor g1505__7098(n_529 ,n_370 ,n_763);
  nor g1506__6131(n_528 ,n_371 ,n_751);
  nor g1507__1881(n_527 ,n_380 ,n_764);
  nor g1508__5115(n_526 ,n_379 ,n_750);
  nor g1509__7482(n_525 ,n_385 ,n_759);
  nor g1510__4733(n_524 ,n_364 ,n_758);
  nor g1511__6161(n_523 ,n_383 ,n_749);
  nor g1512__9315(n_522 ,n_376 ,n_753);
  nor g1513__9945(n_521 ,n_365 ,n_748);
  nor g1514__2883(n_520 ,n_377 ,n_740);
  nor g1515__2346(n_519 ,n_386 ,n_762);
  nor g1516__1666(n_518 ,n_364 ,n_747);
  and g1517__7410(n_517 ,in4 ,out2[24]);
  nor g1518__6417(n_516 ,n_403 ,in7[11]);
  nor g1519__5477(n_515 ,n_398 ,in7[27]);
  and g1520__2398(n_514 ,in4 ,out2[21]);
  and g1521__5107(n_513 ,in4 ,out2[10]);
  nor g1522__6260(n_512 ,n_404 ,in7[10]);
  and g1523__4319(n_511 ,in4 ,out2[31]);
  and g1524__8428(n_510 ,in4 ,out1[0]);
  nor g1525__5526(n_509 ,n_409 ,in7[21]);
  and g1526__6783(n_508 ,in4 ,out2[9]);
  and g1527__3680(n_507 ,in4 ,out2[29]);
  and g1528__1617(n_506 ,in4 ,out2[20]);
  nor g1529__2802(n_505 ,n_389 ,in7[9]);
  and g1530__1705(n_504 ,in4 ,out2[26]);
  or g1531__5122(n_558 ,n_422 ,in4);
  and g1532__8246(n_553 ,n_421 ,n_422);
  and g1533__7098(n_503 ,in4 ,out2[11]);
  nor g1534__6131(n_502 ,n_403 ,in7[20]);
  and g1535__1881(n_501 ,in4 ,out2[7]);
  nor g1536__5115(n_500 ,n_388 ,in7[7]);
  nor g1537__7482(n_499 ,n_407 ,in7[26]);
  and g1538__4733(n_498 ,in4 ,out2[19]);
  and g1539__6161(n_497 ,in4 ,out2[6]);
  nor g1540__9315(n_496 ,n_406 ,in7[6]);
  nor g1541__9945(n_495 ,n_391 ,in7[19]);
  and g1542__2883(n_494 ,in4 ,out1[5]);
  nor g1543__2346(n_493 ,n_409 ,in7[29]);
  nor g1544__1666(n_492 ,n_401 ,in7[5]);
  and g1545__7410(n_491 ,in4 ,out2[25]);
  and g1546__6417(n_490 ,in4 ,out2[18]);
  and g1547__5477(n_489 ,in4 ,out1[4]);
  nor g1548__2398(n_488 ,n_400 ,in7[4]);
  nor g1549__5107(n_487 ,n_394 ,in7[18]);
  and g1550__6260(n_454 ,in4 ,out1[3]);
  nor g1551__4319(n_453 ,n_395 ,in7[3]);
  and g1552__8428(n_452 ,in4 ,out2[28]);
  and g1553__5526(n_451 ,in4 ,out2[17]);
  and g1554__6783(n_450 ,in4 ,out1[2]);
  nor g1555__3680(n_449 ,n_394 ,in7[2]);
  nor g1556__1617(n_448 ,n_397 ,in7[17]);
  and g1557__2802(n_447 ,in4 ,out1[1]);
  nor g1558__1705(n_446 ,n_410 ,in7[1]);
  and g1559__5122(n_445 ,in4 ,out2[16]);
  nor g1560__8246(n_444 ,n_388 ,in7[28]);
  nor g1561__7098(n_443 ,n_389 ,in7[0]);
  nor g1562__6131(n_442 ,n_406 ,in7[16]);
  nor g1563__1881(n_441 ,n_410 ,in7[24]);
  and g1564__5115(n_440 ,in4 ,out2[15]);
  nor g1565__7482(n_439 ,n_391 ,in7[31]);
  nor g1566__4733(n_438 ,n_395 ,in7[15]);
  and g1567__6161(n_437 ,in4 ,out2[30]);
  and g1568__9315(n_436 ,in4 ,out2[23]);
  and g1569__9945(n_435 ,in4 ,out2[14]);
  nor g1570__2883(n_434 ,n_400 ,in7[25]);
  nor g1571__2346(n_433 ,n_404 ,in7[14]);
  nor g1572__1666(n_432 ,n_407 ,in7[23]);
  and g1573__7410(n_431 ,in4 ,out2[13]);
  nor g1574__6417(n_430 ,n_392 ,in7[30]);
  nor g1575__5477(n_429 ,n_401 ,in7[13]);
  and g1576__2398(n_428 ,in4 ,out2[27]);
  and g1577__5107(n_427 ,in4 ,out2[22]);
  and g1578__6260(n_426 ,in4 ,out2[12]);
  nor g1579__4319(n_425 ,n_392 ,in7[12]);
  nor g1580__8428(n_424 ,n_397 ,in7[22]);
  nor g1581__5526(n_423 ,n_398 ,in7[8]);
  not g1582(n_422 ,in5);
  not g1583(n_421 ,in4);
  not g1584(n_420 ,n_362);
  not g1586(n_415 ,n_362);
  not g1588(n_419 ,n_414);
  not g1589(n_418 ,n_419);
  not g1594(n_414 ,in6);
  not g1596(n_417 ,n_355);
  not g1599(n_412 ,n_355);
  not g1600(n_411 ,n_416);
  not g1601(n_413 ,n_416);
  not g1603(n_416 ,in6);
  not drc_bufs1648(n_410 ,n_408);
  not drc_bufs1649(n_409 ,n_408);
  not drc_bufs1650(n_408 ,n_413);
  not drc_bufs1652(n_407 ,n_405);
  not drc_bufs1653(n_406 ,n_405);
  not drc_bufs1654(n_405 ,n_417);
  not drc_bufs1656(n_404 ,n_402);
  not drc_bufs1657(n_403 ,n_402);
  not drc_bufs1658(n_402 ,n_412);
  not drc_bufs1660(n_401 ,n_399);
  not drc_bufs1661(n_400 ,n_399);
  not drc_bufs1662(n_399 ,n_411);
  not drc_bufs1664(n_398 ,n_396);
  not drc_bufs1665(n_397 ,n_396);
  not drc_bufs1666(n_396 ,n_412);
  not drc_bufs1668(n_395 ,n_393);
  not drc_bufs1669(n_394 ,n_393);
  not drc_bufs1670(n_393 ,n_411);
  not drc_bufs1672(n_392 ,n_390);
  not drc_bufs1673(n_391 ,n_390);
  not drc_bufs1674(n_390 ,n_417);
  not drc_bufs1676(n_389 ,n_387);
  not drc_bufs1677(n_388 ,n_387);
  not drc_bufs1678(n_387 ,n_413);
  not drc_bufs1680(n_386 ,n_384);
  not drc_bufs1681(n_385 ,n_384);
  not drc_bufs1682(n_384 ,n_418);
  not drc_bufs1684(n_383 ,n_381);
  not drc_bufs1685(n_382 ,n_381);
  not drc_bufs1686(n_381 ,n_418);
  not drc_bufs1688(n_380 ,n_378);
  not drc_bufs1689(n_379 ,n_378);
  not drc_bufs1690(n_378 ,n_414);
  not drc_bufs1692(n_377 ,n_375);
  not drc_bufs1693(n_376 ,n_375);
  not drc_bufs1694(n_375 ,n_414);
  not drc_bufs1696(n_374 ,n_372);
  not drc_bufs1697(n_373 ,n_372);
  not drc_bufs1698(n_372 ,n_420);
  not drc_bufs1700(n_371 ,n_369);
  not drc_bufs1701(n_370 ,n_369);
  not drc_bufs1702(n_369 ,n_415);
  not drc_bufs1704(n_368 ,n_366);
  not drc_bufs1705(n_367 ,n_366);
  not drc_bufs1706(n_366 ,n_415);
  not drc_bufs1708(n_365 ,n_363);
  not drc_bufs1709(n_364 ,n_363);
  not drc_bufs1710(n_363 ,n_420);
  not drc_bufs1716(n_362 ,n_361);
  not drc_bufs1718(n_361 ,n_419);
  not drc_bufs1721(n_360 ,n_359);
  not drc_bufs1722(n_359 ,n_558);
  not drc_bufs1725(n_358 ,n_357);
  not drc_bufs1726(n_357 ,n_553);
  buf drc_bufs1765(n_36 ,n_726);
  buf drc_bufs1766(n_35 ,n_725);
  buf drc_bufs1767(n_39 ,n_728);
  buf drc_bufs1768(n_38 ,n_727);
  buf drc_bufs1769(n_47 ,n_722);
  buf drc_bufs1770(n_40 ,n_729);
  buf drc_bufs1771(n_49 ,n_723);
  buf drc_bufs1772(n_41 ,n_730);
  buf drc_bufs1773(n_46 ,n_721);
  buf drc_bufs1774(n_34 ,n_724);
  not drc_bufs1777(n_356 ,n_416);
  not drc_bufs1779(n_355 ,n_356);
  not drc_bufs1783(n_354 ,n_352);
  not drc_bufs1784(n_353 ,n_352);
  not drc_bufs1785(n_352 ,n_551);
  not drc_bufs1787(n_351 ,n_349);
  not drc_bufs1788(n_350 ,n_349);
  not drc_bufs1789(n_349 ,n_557);
  not drc_bufs1791(n_348 ,n_346);
  not drc_bufs1792(n_347 ,n_346);
  not drc_bufs1793(n_346 ,n_557);
  not drc_bufs1795(n_345 ,n_343);
  not drc_bufs1796(n_344 ,n_343);
  not drc_bufs1797(n_343 ,n_556);
  not drc_bufs1799(n_342 ,n_340);
  not drc_bufs1800(n_341 ,n_340);
  not drc_bufs1801(n_340 ,n_556);
  not drc_bufs1803(n_339 ,n_337);
  not drc_bufs1804(n_338 ,n_337);
  not drc_bufs1805(n_337 ,n_559);
  not drc_bufs1807(n_336 ,n_334);
  not drc_bufs1808(n_335 ,n_334);
  not drc_bufs1809(n_334 ,n_559);
  not drc_bufs1811(n_333 ,n_331);
  not drc_bufs1812(n_332 ,n_331);
  not drc_bufs1813(n_331 ,n_560);
  not drc_bufs1815(n_330 ,n_328);
  not drc_bufs1816(n_329 ,n_328);
  not drc_bufs1817(n_328 ,n_555);
  not drc_bufs1819(n_327 ,n_325);
  not drc_bufs1820(n_326 ,n_325);
  not drc_bufs1821(n_325 ,n_554);
  not drc_bufs1823(n_324 ,n_322);
  not drc_bufs1824(n_323 ,n_322);
  not drc_bufs1825(n_322 ,n_551);
  not drc_bufs1827(n_321 ,n_319);
  not drc_bufs1828(n_320 ,n_319);
  not drc_bufs1829(n_319 ,n_552);
  not drc_bufs1831(n_318 ,n_316);
  not drc_bufs1832(n_317 ,n_316);
  not drc_bufs1833(n_316 ,n_552);
  not drc_bufs1835(n_315 ,n_313);
  not drc_bufs1836(n_314 ,n_313);
  not drc_bufs1837(n_313 ,n_555);
  not drc_bufs1839(n_312 ,n_310);
  not drc_bufs1840(n_311 ,n_310);
  not drc_bufs1841(n_310 ,n_554);
  not drc_bufs1843(n_309 ,n_307);
  not drc_bufs1844(n_308 ,n_307);
  not drc_bufs1845(n_307 ,n_560);
  buf g577(n_897 ,n_599);
  buf g581(n_893 ,n_598);
  buf g602(n_892 ,n_614);
  buf g585(n_889 ,n_600);
  buf g601(n_888 ,n_601);
  buf g588(n_885 ,n_602);
  buf g598(n_884 ,n_603);
  buf g591(n_882 ,n_604);
  buf g592(n_881 ,n_605);
  buf g582(n_878 ,n_606);
  buf g570(n_877 ,n_607);
  buf g596(n_875 ,n_608);
  buf g597(n_874 ,n_609);
  buf g576(n_871 ,n_610);
  buf g574(n_870 ,n_611);
  buf g575(n_869 ,n_597);
  buf g600(n_868 ,n_612);
  buf g573(n_867 ,n_613);
  not g571(n_866 ,in4);
  not g572(n_865 ,in5);
  and g794__6783(n_7 ,n_874 ,n_853);
  and g798__3680(n_864 ,n_884 ,n_851);
  and g800__1617(n_863 ,n_882 ,n_850);
  and g801__2802(n_862 ,n_881 ,n_847);
  and g803__1705(n_861 ,n_878 ,n_829);
  and g804__5122(n_860 ,n_877 ,n_843);
  and g808__8246(n_859 ,n_875 ,n_840);
  and g810__7098(n_14 ,n_885 ,n_852);
  and g813__6131(n_858 ,n_870 ,n_835);
  and g814__1881(n_19 ,n_869 ,n_832);
  and g815__5115(n_857 ,n_868 ,n_848);
  and g816__7482(n_3 ,n_867 ,n_833);
  and g819__4733(n_18 ,n_893 ,n_836);
  and g820__6161(n_856 ,n_892 ,n_830);
  and g821__9315(n_17 ,n_897 ,n_827);
  and g823__9945(n_855 ,n_889 ,n_825);
  and g824__2883(n_15 ,n_888 ,n_823);
  and g825__2346(n_854 ,n_871 ,n_842);
  nor g826__1666(n_853 ,n_815 ,n_768);
  nor g827__7410(n_852 ,n_816 ,n_789);
  nor g828__6417(n_851 ,n_809 ,n_786);
  nor g829__5477(n_850 ,n_796 ,n_778);
  nor g831__2398(n_848 ,n_814 ,n_772);
  nor g832__5107(n_847 ,n_811 ,n_780);
  nor g836__6260(n_843 ,n_812 ,n_778);
  nor g837__4319(n_842 ,n_814 ,n_771);
  nor g839__8428(n_840 ,n_812 ,n_777);
  nor g843__5526(n_836 ,n_806 ,n_769);
  nor g844__6783(n_835 ,n_816 ,n_790);
  nor g846__3680(n_833 ,n_810 ,n_783);
  nor g847__1617(n_832 ,n_804 ,n_790);
  nor g849__2802(n_830 ,n_796 ,n_777);
  nor g850__1705(n_829 ,n_811 ,n_781);
  nor g852__5122(n_827 ,n_808 ,n_786);
  nor g854__8246(n_825 ,n_794 ,n_783);
  nor g856__7098(n_823 ,n_804 ,n_789);
  not g858(n_821 ,n_792);
  not g859(n_820 ,n_819);
  not g860(n_818 ,n_819);
  not g861(n_817 ,n_792);
  and g862__6131(n_819 ,n_866 ,n_865);
  not g863(n_816 ,in6);
  not g864(n_815 ,in6);
  not g865(n_814 ,in6);
  not g867(n_812 ,in6);
  not g868(n_811 ,in6);
  not g869(n_810 ,in6);
  not g870(n_809 ,in6);
  not drc_bufs891(n_808 ,n_807);
  not drc_bufs892(n_807 ,n_810);
  not drc_bufs895(n_806 ,n_805);
  not drc_bufs896(n_805 ,n_816);
  not drc_bufs899(n_804 ,n_803);
  not drc_bufs900(n_803 ,n_815);
  not drc_bufs915(n_796 ,n_795);
  not drc_bufs916(n_795 ,n_811);
  not drc_bufs919(n_794 ,n_793);
  not drc_bufs920(n_793 ,n_809);
  not drc_bufs923(n_792 ,n_791);
  not drc_bufs924(n_791 ,n_819);
  buf drc_bufs926(n_2 ,n_856);
  buf drc_bufs927(n_4 ,n_857);
  buf drc_bufs928(n_11 ,n_862);
  buf drc_bufs929(n_13 ,n_864);
  buf drc_bufs930(n_5 ,n_858);
  buf drc_bufs931(n_16 ,n_855);
  buf drc_bufs932(n_9 ,n_860);
  buf drc_bufs933(n_10 ,n_861);
  buf drc_bufs934(n_6 ,n_854);
  buf drc_bufs935(n_12 ,n_863);
  buf drc_bufs936(n_8 ,n_859);
  not drc_bufs937(n_790 ,n_788);
  not drc_bufs938(n_789 ,n_788);
  not drc_bufs939(n_788 ,n_821);
  not drc_bufs942(n_786 ,n_785);
  not drc_bufs943(n_785 ,n_817);
  not drc_bufs946(n_783 ,n_782);
  not drc_bufs947(n_782 ,n_817);
  not drc_bufs949(n_781 ,n_779);
  not drc_bufs950(n_780 ,n_779);
  not drc_bufs951(n_779 ,n_818);
  not drc_bufs953(n_778 ,n_776);
  not drc_bufs954(n_777 ,n_776);
  not drc_bufs955(n_776 ,n_818);
  not drc_bufs961(n_772 ,n_770);
  not drc_bufs962(n_771 ,n_770);
  not drc_bufs963(n_770 ,n_820);
  not drc_bufs965(n_769 ,n_767);
  not drc_bufs966(n_768 ,n_767);
  not drc_bufs967(n_767 ,n_821);
  xnor add_25_22_g292__1881(out2[31] ,add_25_22_n_76 ,out1[31]);
  or add_25_22_g294__5115(add_25_22_n_76 ,add_25_22_n_45 ,add_25_22_n_75);
  or add_25_22_g296__7482(add_25_22_n_75 ,add_25_22_n_28 ,add_25_22_n_74);
  or add_25_22_g298__4733(add_25_22_n_74 ,add_25_22_n_27 ,add_25_22_n_73);
  or add_25_22_g300__6161(add_25_22_n_73 ,add_25_22_n_44 ,add_25_22_n_72);
  or add_25_22_g302__9315(add_25_22_n_72 ,add_25_22_n_32 ,add_25_22_n_71);
  or add_25_22_g304__9945(add_25_22_n_71 ,add_25_22_n_29 ,add_25_22_n_70);
  or add_25_22_g306__2883(add_25_22_n_70 ,add_25_22_n_47 ,add_25_22_n_69);
  or add_25_22_g308__2346(add_25_22_n_69 ,add_25_22_n_36 ,add_25_22_n_68);
  or add_25_22_g310__1666(add_25_22_n_68 ,add_25_22_n_34 ,add_25_22_n_67);
  or add_25_22_g312__7410(add_25_22_n_67 ,add_25_22_n_30 ,add_25_22_n_66);
  or add_25_22_g314__6417(add_25_22_n_66 ,add_25_22_n_39 ,add_25_22_n_65);
  or add_25_22_g316__5477(add_25_22_n_65 ,add_25_22_n_41 ,add_25_22_n_64);
  or add_25_22_g318__2398(add_25_22_n_64 ,add_25_22_n_25 ,add_25_22_n_63);
  or add_25_22_g320__5107(add_25_22_n_63 ,add_25_22_n_49 ,add_25_22_n_62);
  or add_25_22_g322__6260(add_25_22_n_62 ,add_25_22_n_26 ,add_25_22_n_61);
  or add_25_22_g324__4319(add_25_22_n_61 ,add_25_22_n_35 ,add_25_22_n_60);
  or add_25_22_g326__8428(add_25_22_n_60 ,add_25_22_n_46 ,add_25_22_n_59);
  or add_25_22_g328__5526(add_25_22_n_59 ,add_25_22_n_33 ,add_25_22_n_58);
  or add_25_22_g330__6783(add_25_22_n_58 ,add_25_22_n_40 ,add_25_22_n_57);
  or add_25_22_g332__3680(add_25_22_n_57 ,add_25_22_n_42 ,add_25_22_n_56);
  or add_25_22_g334__1617(add_25_22_n_56 ,add_25_22_n_48 ,add_25_22_n_55);
  or add_25_22_g336__2802(add_25_22_n_55 ,add_25_22_n_31 ,add_25_22_n_54);
  or add_25_22_g338__1705(add_25_22_n_54 ,add_25_22_n_38 ,add_25_22_n_51);
  and add_25_22_g339__5122(out2[7] ,add_25_22_n_51 ,add_25_22_n_52);
  or add_25_22_g340__8246(add_25_22_n_52 ,add_25_22_n_23 ,add_25_22_n_24);
  or add_25_22_g341__7098(add_25_22_n_51 ,add_25_22_n_43 ,out2[6]);
  not add_25_22_drc_bufs367(add_25_22_n_24 ,out2[6]);
  not add_25_22_drc_bufs372(add_25_22_n_45 ,out1[30]);
  not add_25_22_drc_bufs376(add_25_22_n_28 ,out1[29]);
  not add_25_22_drc_bufs380(add_25_22_n_27 ,out1[28]);
  not add_25_22_drc_bufs384(add_25_22_n_44 ,out1[27]);
  not add_25_22_drc_bufs388(add_25_22_n_32 ,out1[26]);
  not add_25_22_drc_bufs392(add_25_22_n_29 ,out1[25]);
  not add_25_22_drc_bufs396(add_25_22_n_47 ,out1[24]);
  not add_25_22_drc_bufs400(add_25_22_n_36 ,out1[23]);
  not add_25_22_drc_bufs404(add_25_22_n_34 ,out1[22]);
  not add_25_22_drc_bufs408(add_25_22_n_31 ,out1[9]);
  not add_25_22_drc_bufs412(add_25_22_n_39 ,out1[20]);
  not add_25_22_drc_bufs416(add_25_22_n_41 ,out1[19]);
  not add_25_22_drc_bufs420(add_25_22_n_25 ,out1[18]);
  not add_25_22_drc_bufs424(add_25_22_n_49 ,out1[17]);
  not add_25_22_drc_bufs428(add_25_22_n_26 ,out1[16]);
  not add_25_22_drc_bufs432(add_25_22_n_35 ,out1[15]);
  not add_25_22_drc_bufs436(add_25_22_n_46 ,out1[14]);
  not add_25_22_drc_bufs440(add_25_22_n_33 ,out1[13]);
  not add_25_22_drc_bufs444(add_25_22_n_40 ,out1[12]);
  not add_25_22_drc_bufs448(add_25_22_n_42 ,out1[11]);
  not add_25_22_drc_bufs452(add_25_22_n_48 ,out1[10]);
  not add_25_22_drc_bufs456(add_25_22_n_30 ,out1[21]);
  not add_25_22_drc_bufs460(add_25_22_n_38 ,out1[8]);
  not add_25_22_drc_bufs463(add_25_22_n_23 ,add_25_22_n_43);
  not add_25_22_drc_bufs464(add_25_22_n_43 ,out1[7]);
  xor add_25_22_g2__6131(out2[30] ,add_25_22_n_75 ,add_25_22_n_45);
  xor add_25_22_g467__1881(out2[29] ,add_25_22_n_74 ,add_25_22_n_28);
  xor add_25_22_g468__5115(out2[28] ,add_25_22_n_73 ,add_25_22_n_27);
  xor add_25_22_g469__7482(out2[27] ,add_25_22_n_72 ,add_25_22_n_44);
  xor add_25_22_g470__4733(out2[26] ,add_25_22_n_71 ,add_25_22_n_32);
  xor add_25_22_g471__6161(out2[25] ,add_25_22_n_70 ,add_25_22_n_29);
  xor add_25_22_g472__9315(out2[24] ,add_25_22_n_69 ,add_25_22_n_47);
  xor add_25_22_g473__9945(out2[23] ,add_25_22_n_68 ,add_25_22_n_36);
  xor add_25_22_g474__2883(out2[22] ,add_25_22_n_67 ,add_25_22_n_34);
  xor add_25_22_g475__2346(out2[9] ,add_25_22_n_54 ,add_25_22_n_31);
  xor add_25_22_g476__1666(out2[20] ,add_25_22_n_65 ,add_25_22_n_39);
  xor add_25_22_g477__7410(out2[19] ,add_25_22_n_64 ,add_25_22_n_41);
  xor add_25_22_g478__6417(out2[18] ,add_25_22_n_63 ,add_25_22_n_25);
  xor add_25_22_g479__5477(out2[17] ,add_25_22_n_62 ,add_25_22_n_49);
  xor add_25_22_g480__2398(out2[16] ,add_25_22_n_61 ,add_25_22_n_26);
  xor add_25_22_g481__5107(out2[15] ,add_25_22_n_60 ,add_25_22_n_35);
  xor add_25_22_g482__6260(out2[14] ,add_25_22_n_59 ,add_25_22_n_46);
  xor add_25_22_g483__4319(out2[13] ,add_25_22_n_58 ,add_25_22_n_33);
  xor add_25_22_g484__8428(out2[12] ,add_25_22_n_57 ,add_25_22_n_40);
  xor add_25_22_g485__5526(out2[11] ,add_25_22_n_56 ,add_25_22_n_42);
  xor add_25_22_g486__6783(out2[10] ,add_25_22_n_55 ,add_25_22_n_48);
  xor add_25_22_g487__3680(out2[21] ,add_25_22_n_66 ,add_25_22_n_30);
  xor add_25_22_g488__1617(out2[8] ,add_25_22_n_51 ,add_25_22_n_38);
  xnor csa_tree_add_22_22_g3336__2802(n_601 ,csa_tree_add_22_22_n_441 ,csa_tree_add_22_22_n_491);
  xnor csa_tree_add_22_22_g3337__1705(n_602 ,csa_tree_add_22_22_n_443 ,csa_tree_add_22_22_n_492);
  xnor csa_tree_add_22_22_g3338__5122(n_603 ,csa_tree_add_22_22_n_467 ,csa_tree_add_22_22_n_494);
  xnor csa_tree_add_22_22_g3339__8246(n_604 ,csa_tree_add_22_22_n_468 ,csa_tree_add_22_22_n_497);
  xnor csa_tree_add_22_22_g3340__7098(n_605 ,csa_tree_add_22_22_n_466 ,csa_tree_add_22_22_n_496);
  xnor csa_tree_add_22_22_g3341__6131(n_606 ,csa_tree_add_22_22_n_469 ,csa_tree_add_22_22_n_495);
  xnor csa_tree_add_22_22_g3342__1881(n_607 ,csa_tree_add_22_22_n_440 ,csa_tree_add_22_22_n_498);
  xnor csa_tree_add_22_22_g3343__5115(n_608 ,csa_tree_add_22_22_n_442 ,csa_tree_add_22_22_n_493);
  or csa_tree_add_22_22_g3344__7482(n_473 ,csa_tree_add_22_22_n_488 ,csa_tree_add_22_22_n_508);
  or csa_tree_add_22_22_g3345__4733(n_476 ,csa_tree_add_22_22_n_489 ,csa_tree_add_22_22_n_510);
  or csa_tree_add_22_22_g3346__6161(n_472 ,csa_tree_add_22_22_n_479 ,csa_tree_add_22_22_n_504);
  or csa_tree_add_22_22_g3347__9315(n_477 ,csa_tree_add_22_22_n_485 ,csa_tree_add_22_22_n_507);
  or csa_tree_add_22_22_g3348__9945(n_474 ,csa_tree_add_22_22_n_475 ,csa_tree_add_22_22_n_505);
  or csa_tree_add_22_22_g3349__2883(n_478 ,csa_tree_add_22_22_n_481 ,csa_tree_add_22_22_n_506);
  or csa_tree_add_22_22_g3350__2346(n_479 ,csa_tree_add_22_22_n_477 ,csa_tree_add_22_22_n_503);
  or csa_tree_add_22_22_g3351__1666(n_475 ,csa_tree_add_22_22_n_474 ,csa_tree_add_22_22_n_501);
  nor csa_tree_add_22_22_g3352__7410(csa_tree_add_22_22_n_510 ,csa_tree_add_22_22_n_466 ,csa_tree_add_22_22_n_486);
  or csa_tree_add_22_22_g3353__6417(n_471 ,csa_tree_add_22_22_n_462 ,csa_tree_add_22_22_n_484);
  nor csa_tree_add_22_22_g3354__5477(csa_tree_add_22_22_n_508 ,csa_tree_add_22_22_n_443 ,csa_tree_add_22_22_n_483);
  nor csa_tree_add_22_22_g3355__2398(csa_tree_add_22_22_n_507 ,csa_tree_add_22_22_n_469 ,csa_tree_add_22_22_n_482);
  nor csa_tree_add_22_22_g3356__5107(csa_tree_add_22_22_n_506 ,csa_tree_add_22_22_n_440 ,csa_tree_add_22_22_n_478);
  nor csa_tree_add_22_22_g3357__6260(csa_tree_add_22_22_n_505 ,csa_tree_add_22_22_n_467 ,csa_tree_add_22_22_n_480);
  nor csa_tree_add_22_22_g3358__4319(csa_tree_add_22_22_n_504 ,csa_tree_add_22_22_n_441 ,csa_tree_add_22_22_n_487);
  nor csa_tree_add_22_22_g3359__8428(csa_tree_add_22_22_n_503 ,csa_tree_add_22_22_n_442 ,csa_tree_add_22_22_n_476);
  or csa_tree_add_22_22_g3360__5526(n_480 ,csa_tree_add_22_22_n_415 ,csa_tree_add_22_22_n_473);
  nor csa_tree_add_22_22_g3361__6783(csa_tree_add_22_22_n_501 ,csa_tree_add_22_22_n_468 ,csa_tree_add_22_22_n_490);
  xnor csa_tree_add_22_22_g3362__3680(n_600 ,csa_tree_add_22_22_n_439 ,csa_tree_add_22_22_n_461);
  xnor csa_tree_add_22_22_g3363__1617(n_609 ,csa_tree_add_22_22_n_460 ,csa_tree_add_22_22_n_429);
  xnor csa_tree_add_22_22_g3364__2802(csa_tree_add_22_22_n_498 ,csa_tree_add_22_22_n_355 ,csa_tree_add_22_22_n_452);
  xnor csa_tree_add_22_22_g3365__1705(csa_tree_add_22_22_n_497 ,csa_tree_add_22_22_n_349 ,csa_tree_add_22_22_n_444);
  xnor csa_tree_add_22_22_g3366__5122(csa_tree_add_22_22_n_496 ,csa_tree_add_22_22_n_359 ,csa_tree_add_22_22_n_458);
  xnor csa_tree_add_22_22_g3367__8246(csa_tree_add_22_22_n_495 ,csa_tree_add_22_22_n_356 ,csa_tree_add_22_22_n_454);
  xnor csa_tree_add_22_22_g3368__7098(csa_tree_add_22_22_n_494 ,csa_tree_add_22_22_n_354 ,csa_tree_add_22_22_n_450);
  xnor csa_tree_add_22_22_g3369__6131(csa_tree_add_22_22_n_493 ,csa_tree_add_22_22_n_352 ,csa_tree_add_22_22_n_448);
  xnor csa_tree_add_22_22_g3370__1881(csa_tree_add_22_22_n_492 ,csa_tree_add_22_22_n_346 ,csa_tree_add_22_22_n_456);
  xnor csa_tree_add_22_22_g3371__5115(csa_tree_add_22_22_n_491 ,csa_tree_add_22_22_n_353 ,csa_tree_add_22_22_n_446);
  and csa_tree_add_22_22_g3372__7482(csa_tree_add_22_22_n_490 ,csa_tree_add_22_22_n_349 ,csa_tree_add_22_22_n_445);
  nor csa_tree_add_22_22_g3373__4733(csa_tree_add_22_22_n_489 ,csa_tree_add_22_22_n_359 ,csa_tree_add_22_22_n_459);
  nor csa_tree_add_22_22_g3374__6161(csa_tree_add_22_22_n_488 ,csa_tree_add_22_22_n_346 ,csa_tree_add_22_22_n_457);
  and csa_tree_add_22_22_g3375__9315(csa_tree_add_22_22_n_487 ,csa_tree_add_22_22_n_353 ,csa_tree_add_22_22_n_447);
  and csa_tree_add_22_22_g3376__9945(csa_tree_add_22_22_n_486 ,csa_tree_add_22_22_n_359 ,csa_tree_add_22_22_n_459);
  nor csa_tree_add_22_22_g3377__2883(csa_tree_add_22_22_n_485 ,csa_tree_add_22_22_n_356 ,csa_tree_add_22_22_n_455);
  nor csa_tree_add_22_22_g3378__2346(csa_tree_add_22_22_n_484 ,csa_tree_add_22_22_n_411 ,csa_tree_add_22_22_n_463);
  and csa_tree_add_22_22_g3379__1666(csa_tree_add_22_22_n_483 ,csa_tree_add_22_22_n_346 ,csa_tree_add_22_22_n_457);
  and csa_tree_add_22_22_g3380__7410(csa_tree_add_22_22_n_482 ,csa_tree_add_22_22_n_356 ,csa_tree_add_22_22_n_455);
  nor csa_tree_add_22_22_g3381__6417(csa_tree_add_22_22_n_481 ,csa_tree_add_22_22_n_355 ,csa_tree_add_22_22_n_453);
  and csa_tree_add_22_22_g3382__5477(csa_tree_add_22_22_n_480 ,csa_tree_add_22_22_n_354 ,csa_tree_add_22_22_n_451);
  nor csa_tree_add_22_22_g3383__2398(csa_tree_add_22_22_n_479 ,csa_tree_add_22_22_n_353 ,csa_tree_add_22_22_n_447);
  and csa_tree_add_22_22_g3384__5107(csa_tree_add_22_22_n_478 ,csa_tree_add_22_22_n_355 ,csa_tree_add_22_22_n_453);
  nor csa_tree_add_22_22_g3385__6260(csa_tree_add_22_22_n_477 ,csa_tree_add_22_22_n_352 ,csa_tree_add_22_22_n_449);
  and csa_tree_add_22_22_g3386__4319(csa_tree_add_22_22_n_476 ,csa_tree_add_22_22_n_352 ,csa_tree_add_22_22_n_449);
  nor csa_tree_add_22_22_g3387__8428(csa_tree_add_22_22_n_475 ,csa_tree_add_22_22_n_354 ,csa_tree_add_22_22_n_451);
  nor csa_tree_add_22_22_g3388__5526(csa_tree_add_22_22_n_474 ,csa_tree_add_22_22_n_349 ,csa_tree_add_22_22_n_445);
  and csa_tree_add_22_22_g3389__6783(csa_tree_add_22_22_n_473 ,csa_tree_add_22_22_n_413 ,csa_tree_add_22_22_n_460);
  or csa_tree_add_22_22_g3390__3680(n_481 ,csa_tree_add_22_22_n_412 ,csa_tree_add_22_22_n_464);
  xnor csa_tree_add_22_22_g3391__1617(n_610 ,csa_tree_add_22_22_n_435 ,csa_tree_add_22_22_n_428);
  xnor csa_tree_add_22_22_g3392__2802(n_599 ,csa_tree_add_22_22_n_427 ,csa_tree_add_22_22_n_430);
  or csa_tree_add_22_22_g3393__1705(n_598 ,csa_tree_add_22_22_n_405 ,csa_tree_add_22_22_n_436);
  and csa_tree_add_22_22_g3394__5122(csa_tree_add_22_22_n_464 ,csa_tree_add_22_22_n_426 ,csa_tree_add_22_22_n_435);
  and csa_tree_add_22_22_g3395__8246(csa_tree_add_22_22_n_463 ,csa_tree_add_22_22_n_392 ,csa_tree_add_22_22_n_439);
  nor csa_tree_add_22_22_g3396__7098(csa_tree_add_22_22_n_462 ,csa_tree_add_22_22_n_392 ,csa_tree_add_22_22_n_439);
  xnor csa_tree_add_22_22_g3397__6131(csa_tree_add_22_22_n_461 ,csa_tree_add_22_22_n_391 ,csa_tree_add_22_22_n_411);
  and csa_tree_add_22_22_g3398__1881(csa_tree_add_22_22_n_469 ,csa_tree_add_22_22_n_421 ,csa_tree_add_22_22_n_434);
  and csa_tree_add_22_22_g3399__5115(csa_tree_add_22_22_n_468 ,csa_tree_add_22_22_n_409 ,csa_tree_add_22_22_n_432);
  and csa_tree_add_22_22_g3400__7482(csa_tree_add_22_22_n_467 ,csa_tree_add_22_22_n_417 ,csa_tree_add_22_22_n_431);
  and csa_tree_add_22_22_g3401__4733(csa_tree_add_22_22_n_466 ,csa_tree_add_22_22_n_424 ,csa_tree_add_22_22_n_438);
  not csa_tree_add_22_22_g3402(csa_tree_add_22_22_n_459 ,csa_tree_add_22_22_n_458);
  not csa_tree_add_22_22_g3403(csa_tree_add_22_22_n_457 ,csa_tree_add_22_22_n_456);
  not csa_tree_add_22_22_g3404(csa_tree_add_22_22_n_455 ,csa_tree_add_22_22_n_454);
  not csa_tree_add_22_22_g3405(csa_tree_add_22_22_n_453 ,csa_tree_add_22_22_n_452);
  not csa_tree_add_22_22_g3406(csa_tree_add_22_22_n_451 ,csa_tree_add_22_22_n_450);
  not csa_tree_add_22_22_g3407(csa_tree_add_22_22_n_449 ,csa_tree_add_22_22_n_448);
  not csa_tree_add_22_22_g3408(csa_tree_add_22_22_n_447 ,csa_tree_add_22_22_n_446);
  not csa_tree_add_22_22_g3409(csa_tree_add_22_22_n_445 ,csa_tree_add_22_22_n_444);
  xnor csa_tree_add_22_22_g3410__6161(csa_tree_add_22_22_n_460 ,csa_tree_add_22_22_n_364 ,csa_tree_add_22_22_n_395);
  xnor csa_tree_add_22_22_g3411__9315(csa_tree_add_22_22_n_458 ,csa_tree_add_22_22_n_363 ,csa_tree_add_22_22_n_396);
  xnor csa_tree_add_22_22_g3412__9945(csa_tree_add_22_22_n_456 ,csa_tree_add_22_22_n_366 ,csa_tree_add_22_22_n_403);
  xnor csa_tree_add_22_22_g3413__2883(csa_tree_add_22_22_n_454 ,csa_tree_add_22_22_n_390 ,csa_tree_add_22_22_n_402);
  xnor csa_tree_add_22_22_g3414__2346(csa_tree_add_22_22_n_452 ,csa_tree_add_22_22_n_388 ,csa_tree_add_22_22_n_401);
  xnor csa_tree_add_22_22_g3415__1666(csa_tree_add_22_22_n_450 ,csa_tree_add_22_22_n_393 ,csa_tree_add_22_22_n_400);
  xnor csa_tree_add_22_22_g3416__7410(csa_tree_add_22_22_n_448 ,csa_tree_add_22_22_n_368 ,csa_tree_add_22_22_n_399);
  xnor csa_tree_add_22_22_g3417__6417(csa_tree_add_22_22_n_446 ,csa_tree_add_22_22_n_343 ,csa_tree_add_22_22_n_398);
  xnor csa_tree_add_22_22_g3418__5477(csa_tree_add_22_22_n_444 ,csa_tree_add_22_22_n_358 ,csa_tree_add_22_22_n_397);
  or csa_tree_add_22_22_g3419__2398(csa_tree_add_22_22_n_438 ,csa_tree_add_22_22_n_341 ,csa_tree_add_22_22_n_422);
  or csa_tree_add_22_22_g3420__5107(n_482 ,csa_tree_add_22_22_n_315 ,csa_tree_add_22_22_n_408);
  nor csa_tree_add_22_22_g3421__6260(csa_tree_add_22_22_n_436 ,csa_tree_add_22_22_n_427 ,csa_tree_add_22_22_n_425);
  and csa_tree_add_22_22_g3422__4319(csa_tree_add_22_22_n_443 ,csa_tree_add_22_22_n_381 ,csa_tree_add_22_22_n_419);
  and csa_tree_add_22_22_g3423__8428(csa_tree_add_22_22_n_442 ,csa_tree_add_22_22_n_377 ,csa_tree_add_22_22_n_416);
  and csa_tree_add_22_22_g3424__5526(csa_tree_add_22_22_n_441 ,csa_tree_add_22_22_n_373 ,csa_tree_add_22_22_n_410);
  and csa_tree_add_22_22_g3425__6783(csa_tree_add_22_22_n_440 ,csa_tree_add_22_22_n_379 ,csa_tree_add_22_22_n_418);
  and csa_tree_add_22_22_g3426__3680(csa_tree_add_22_22_n_439 ,csa_tree_add_22_22_n_384 ,csa_tree_add_22_22_n_423);
  or csa_tree_add_22_22_g3427__1617(csa_tree_add_22_22_n_434 ,csa_tree_add_22_22_n_340 ,csa_tree_add_22_22_n_420);
  xnor csa_tree_add_22_22_g3428__2802(n_611 ,csa_tree_add_22_22_n_370 ,csa_tree_add_22_22_n_345);
  or csa_tree_add_22_22_g3429__1705(csa_tree_add_22_22_n_432 ,csa_tree_add_22_22_n_327 ,csa_tree_add_22_22_n_407);
  or csa_tree_add_22_22_g3430__5122(csa_tree_add_22_22_n_431 ,csa_tree_add_22_22_n_342 ,csa_tree_add_22_22_n_414);
  xnor csa_tree_add_22_22_g3431__8246(csa_tree_add_22_22_n_430 ,csa_tree_add_22_22_n_322 ,csa_tree_add_22_22_n_360);
  xnor csa_tree_add_22_22_g3432__7098(csa_tree_add_22_22_n_429 ,csa_tree_add_22_22_n_351 ,csa_tree_add_22_22_n_386);
  xnor csa_tree_add_22_22_g3433__6131(csa_tree_add_22_22_n_428 ,csa_tree_add_22_22_n_348 ,csa_tree_add_22_22_n_319);
  xnor csa_tree_add_22_22_g3434__1881(csa_tree_add_22_22_n_435 ,csa_tree_add_22_22_n_255 ,csa_tree_add_22_22_n_344);
  or csa_tree_add_22_22_g3435__5115(csa_tree_add_22_22_n_426 ,csa_tree_add_22_22_n_318 ,csa_tree_add_22_22_n_347);
  and csa_tree_add_22_22_g3436__7482(csa_tree_add_22_22_n_425 ,csa_tree_add_22_22_n_322 ,csa_tree_add_22_22_n_361);
  or csa_tree_add_22_22_g3437__4733(csa_tree_add_22_22_n_424 ,csa_tree_add_22_22_n_329 ,csa_tree_add_22_22_n_389);
  or csa_tree_add_22_22_g3438__6161(csa_tree_add_22_22_n_423 ,csa_tree_add_22_22_n_343 ,csa_tree_add_22_22_n_383);
  nor csa_tree_add_22_22_g3439__9315(csa_tree_add_22_22_n_422 ,csa_tree_add_22_22_n_328 ,csa_tree_add_22_22_n_390);
  or csa_tree_add_22_22_g3440__9945(csa_tree_add_22_22_n_421 ,csa_tree_add_22_22_n_336 ,csa_tree_add_22_22_n_387);
  nor csa_tree_add_22_22_g3441__2883(csa_tree_add_22_22_n_420 ,csa_tree_add_22_22_n_335 ,csa_tree_add_22_22_n_388);
  or csa_tree_add_22_22_g3442__2346(csa_tree_add_22_22_n_419 ,csa_tree_add_22_22_n_394 ,csa_tree_add_22_22_n_380);
  or csa_tree_add_22_22_g3443__1666(csa_tree_add_22_22_n_418 ,csa_tree_add_22_22_n_369 ,csa_tree_add_22_22_n_378);
  or csa_tree_add_22_22_g3444__7410(csa_tree_add_22_22_n_417 ,csa_tree_add_22_22_n_338 ,csa_tree_add_22_22_n_357);
  or csa_tree_add_22_22_g3445__6417(csa_tree_add_22_22_n_416 ,csa_tree_add_22_22_n_376 ,csa_tree_add_22_22_n_365);
  nor csa_tree_add_22_22_g3446__5477(csa_tree_add_22_22_n_415 ,csa_tree_add_22_22_n_386 ,csa_tree_add_22_22_n_351);
  nor csa_tree_add_22_22_g3447__2398(csa_tree_add_22_22_n_414 ,csa_tree_add_22_22_n_337 ,csa_tree_add_22_22_n_358);
  or csa_tree_add_22_22_g3448__5107(csa_tree_add_22_22_n_413 ,csa_tree_add_22_22_n_385 ,csa_tree_add_22_22_n_350);
  nor csa_tree_add_22_22_g3449__6260(csa_tree_add_22_22_n_412 ,csa_tree_add_22_22_n_319 ,csa_tree_add_22_22_n_348);
  and csa_tree_add_22_22_g3450__4319(csa_tree_add_22_22_n_427 ,csa_tree_add_22_22_n_298 ,csa_tree_add_22_22_n_375);
  or csa_tree_add_22_22_g3451__8428(csa_tree_add_22_22_n_410 ,csa_tree_add_22_22_n_367 ,csa_tree_add_22_22_n_382);
  or csa_tree_add_22_22_g3452__5526(csa_tree_add_22_22_n_409 ,csa_tree_add_22_22_n_325 ,csa_tree_add_22_22_n_362);
  nor csa_tree_add_22_22_g3453__6783(csa_tree_add_22_22_n_408 ,csa_tree_add_22_22_n_313 ,csa_tree_add_22_22_n_370);
  nor csa_tree_add_22_22_g3454__3680(csa_tree_add_22_22_n_407 ,csa_tree_add_22_22_n_324 ,csa_tree_add_22_22_n_363);
  or csa_tree_add_22_22_g3455__1617(n_597 ,csa_tree_add_22_22_n_243 ,csa_tree_add_22_22_n_371);
  nor csa_tree_add_22_22_g3456__2802(csa_tree_add_22_22_n_405 ,csa_tree_add_22_22_n_322 ,csa_tree_add_22_22_n_361);
  xnor csa_tree_add_22_22_g3457__1705(n_470 ,csa_tree_add_22_22_n_326 ,csa_tree_add_22_22_n_278);
  xnor csa_tree_add_22_22_g3458__5122(csa_tree_add_22_22_n_403 ,csa_tree_add_22_22_n_323 ,csa_tree_add_22_22_n_317);
  xnor csa_tree_add_22_22_g3459__8246(csa_tree_add_22_22_n_402 ,csa_tree_add_22_22_n_329 ,csa_tree_add_22_22_n_341);
  xnor csa_tree_add_22_22_g3460__7098(csa_tree_add_22_22_n_401 ,csa_tree_add_22_22_n_336 ,csa_tree_add_22_22_n_340);
  xnor csa_tree_add_22_22_g3461__6131(csa_tree_add_22_22_n_400 ,csa_tree_add_22_22_n_332 ,csa_tree_add_22_22_n_331);
  xnor csa_tree_add_22_22_g3462__1881(csa_tree_add_22_22_n_399 ,csa_tree_add_22_22_n_333 ,csa_tree_add_22_22_n_334);
  xnor csa_tree_add_22_22_g3463__5115(csa_tree_add_22_22_n_398 ,csa_tree_add_22_22_n_281 ,csa_tree_add_22_22_n_321);
  xnor csa_tree_add_22_22_g3464__7482(csa_tree_add_22_22_n_397 ,csa_tree_add_22_22_n_338 ,csa_tree_add_22_22_n_342);
  xnor csa_tree_add_22_22_g3465__4733(csa_tree_add_22_22_n_396 ,csa_tree_add_22_22_n_325 ,csa_tree_add_22_22_n_327);
  xnor csa_tree_add_22_22_g3466__6161(csa_tree_add_22_22_n_395 ,csa_tree_add_22_22_n_256 ,csa_tree_add_22_22_n_330);
  xnor csa_tree_add_22_22_g3467__9315(csa_tree_add_22_22_n_411 ,csa_tree_add_22_22_n_339 ,csa_tree_add_22_22_n_312);
  not csa_tree_add_22_22_g3468(csa_tree_add_22_22_n_394 ,csa_tree_add_22_22_n_393);
  not csa_tree_add_22_22_g3469(csa_tree_add_22_22_n_392 ,csa_tree_add_22_22_n_391);
  not csa_tree_add_22_22_g3470(csa_tree_add_22_22_n_389 ,csa_tree_add_22_22_n_390);
  not csa_tree_add_22_22_g3471(csa_tree_add_22_22_n_387 ,csa_tree_add_22_22_n_388);
  not csa_tree_add_22_22_g3472(csa_tree_add_22_22_n_386 ,csa_tree_add_22_22_n_385);
  or csa_tree_add_22_22_g3473__9945(csa_tree_add_22_22_n_384 ,csa_tree_add_22_22_n_280 ,csa_tree_add_22_22_n_321);
  nor csa_tree_add_22_22_g3474__2883(csa_tree_add_22_22_n_383 ,csa_tree_add_22_22_n_281 ,csa_tree_add_22_22_n_320);
  and csa_tree_add_22_22_g3475__2346(csa_tree_add_22_22_n_382 ,csa_tree_add_22_22_n_317 ,csa_tree_add_22_22_n_323);
  or csa_tree_add_22_22_g3476__1666(csa_tree_add_22_22_n_381 ,csa_tree_add_22_22_n_331 ,csa_tree_add_22_22_n_332);
  and csa_tree_add_22_22_g3477__7410(csa_tree_add_22_22_n_380 ,csa_tree_add_22_22_n_331 ,csa_tree_add_22_22_n_332);
  or csa_tree_add_22_22_g3478__6417(csa_tree_add_22_22_n_379 ,csa_tree_add_22_22_n_334 ,csa_tree_add_22_22_n_333);
  and csa_tree_add_22_22_g3479__5477(csa_tree_add_22_22_n_378 ,csa_tree_add_22_22_n_334 ,csa_tree_add_22_22_n_333);
  or csa_tree_add_22_22_g3480__2398(csa_tree_add_22_22_n_377 ,csa_tree_add_22_22_n_256 ,csa_tree_add_22_22_n_330);
  and csa_tree_add_22_22_g3481__5107(csa_tree_add_22_22_n_376 ,csa_tree_add_22_22_n_256 ,csa_tree_add_22_22_n_330);
  or csa_tree_add_22_22_g3482__6260(csa_tree_add_22_22_n_375 ,csa_tree_add_22_22_n_295 ,csa_tree_add_22_22_n_339);
  xnor csa_tree_add_22_22_g3483__4319(n_612 ,csa_tree_add_22_22_n_285 ,csa_tree_add_22_22_n_262);
  or csa_tree_add_22_22_g3484__8428(csa_tree_add_22_22_n_373 ,csa_tree_add_22_22_n_317 ,csa_tree_add_22_22_n_323);
  or csa_tree_add_22_22_g3485__5526(n_483 ,csa_tree_add_22_22_n_206 ,csa_tree_add_22_22_n_316);
  nor csa_tree_add_22_22_g3486__6783(csa_tree_add_22_22_n_371 ,csa_tree_add_22_22_n_229 ,csa_tree_add_22_22_n_326);
  xnor csa_tree_add_22_22_g3487__3680(csa_tree_add_22_22_n_393 ,csa_tree_add_22_22_n_171 ,csa_tree_add_22_22_n_272);
  xnor csa_tree_add_22_22_g3488__1617(csa_tree_add_22_22_n_391 ,csa_tree_add_22_22_n_148 ,csa_tree_add_22_22_n_271);
  xnor csa_tree_add_22_22_g3489__2802(csa_tree_add_22_22_n_390 ,csa_tree_add_22_22_n_151 ,csa_tree_add_22_22_n_268);
  xnor csa_tree_add_22_22_g3490__1705(csa_tree_add_22_22_n_388 ,csa_tree_add_22_22_n_134 ,csa_tree_add_22_22_n_273);
  or csa_tree_add_22_22_g3491__5122(csa_tree_add_22_22_n_385 ,csa_tree_add_22_22_n_297 ,csa_tree_add_22_22_n_314);
  not csa_tree_add_22_22_g3492(csa_tree_add_22_22_n_369 ,csa_tree_add_22_22_n_368);
  not csa_tree_add_22_22_g3493(csa_tree_add_22_22_n_367 ,csa_tree_add_22_22_n_366);
  not csa_tree_add_22_22_g3494(csa_tree_add_22_22_n_365 ,csa_tree_add_22_22_n_364);
  not csa_tree_add_22_22_g3495(csa_tree_add_22_22_n_362 ,csa_tree_add_22_22_n_363);
  not csa_tree_add_22_22_g3496(csa_tree_add_22_22_n_361 ,csa_tree_add_22_22_n_360);
  not csa_tree_add_22_22_g3497(csa_tree_add_22_22_n_357 ,csa_tree_add_22_22_n_358);
  not csa_tree_add_22_22_g3498(csa_tree_add_22_22_n_350 ,csa_tree_add_22_22_n_351);
  not csa_tree_add_22_22_g3499(csa_tree_add_22_22_n_347 ,csa_tree_add_22_22_n_348);
  xnor csa_tree_add_22_22_g3500__8246(csa_tree_add_22_22_n_345 ,csa_tree_add_22_22_n_252 ,csa_tree_add_22_22_n_282);
  xnor csa_tree_add_22_22_g3501__7098(csa_tree_add_22_22_n_344 ,csa_tree_add_22_22_n_139 ,csa_tree_add_22_22_n_284);
  xnor csa_tree_add_22_22_g3502__6131(csa_tree_add_22_22_n_370 ,csa_tree_add_22_22_n_191 ,csa_tree_add_22_22_n_265);
  xnor csa_tree_add_22_22_g3503__1881(csa_tree_add_22_22_n_368 ,csa_tree_add_22_22_n_179 ,csa_tree_add_22_22_n_269);
  xnor csa_tree_add_22_22_g3504__5115(csa_tree_add_22_22_n_366 ,csa_tree_add_22_22_n_129 ,csa_tree_add_22_22_n_279);
  xnor csa_tree_add_22_22_g3505__7482(csa_tree_add_22_22_n_364 ,csa_tree_add_22_22_n_146 ,csa_tree_add_22_22_n_276);
  xnor csa_tree_add_22_22_g3506__4733(csa_tree_add_22_22_n_363 ,csa_tree_add_22_22_n_142 ,csa_tree_add_22_22_n_275);
  xnor csa_tree_add_22_22_g3507__6161(csa_tree_add_22_22_n_360 ,csa_tree_add_22_22_n_186 ,csa_tree_add_22_22_n_270);
  xnor csa_tree_add_22_22_g3508__9315(csa_tree_add_22_22_n_359 ,csa_tree_add_22_22_n_140 ,csa_tree_add_22_22_n_258);
  xnor csa_tree_add_22_22_g3509__9945(csa_tree_add_22_22_n_358 ,csa_tree_add_22_22_n_183 ,csa_tree_add_22_22_n_274);
  xnor csa_tree_add_22_22_g3510__2883(csa_tree_add_22_22_n_356 ,csa_tree_add_22_22_n_176 ,csa_tree_add_22_22_n_261);
  xnor csa_tree_add_22_22_g3511__2346(csa_tree_add_22_22_n_355 ,csa_tree_add_22_22_n_132 ,csa_tree_add_22_22_n_260);
  xnor csa_tree_add_22_22_g3512__1666(csa_tree_add_22_22_n_354 ,csa_tree_add_22_22_n_143 ,csa_tree_add_22_22_n_259);
  xnor csa_tree_add_22_22_g3513__7410(csa_tree_add_22_22_n_353 ,csa_tree_add_22_22_n_189 ,csa_tree_add_22_22_n_267);
  xnor csa_tree_add_22_22_g3514__6417(csa_tree_add_22_22_n_352 ,csa_tree_add_22_22_n_155 ,csa_tree_add_22_22_n_266);
  xnor csa_tree_add_22_22_g3515__5477(csa_tree_add_22_22_n_351 ,csa_tree_add_22_22_n_128 ,csa_tree_add_22_22_n_277);
  xnor csa_tree_add_22_22_g3516__2398(csa_tree_add_22_22_n_349 ,csa_tree_add_22_22_n_174 ,csa_tree_add_22_22_n_257);
  xnor csa_tree_add_22_22_g3517__5107(csa_tree_add_22_22_n_348 ,csa_tree_add_22_22_n_159 ,csa_tree_add_22_22_n_263);
  xnor csa_tree_add_22_22_g3518__6260(csa_tree_add_22_22_n_346 ,csa_tree_add_22_22_n_131 ,csa_tree_add_22_22_n_264);
  not csa_tree_add_22_22_g3519(csa_tree_add_22_22_n_337 ,csa_tree_add_22_22_n_338);
  not csa_tree_add_22_22_g3520(csa_tree_add_22_22_n_335 ,csa_tree_add_22_22_n_336);
  not csa_tree_add_22_22_g3521(csa_tree_add_22_22_n_328 ,csa_tree_add_22_22_n_329);
  and csa_tree_add_22_22_g3522__4319(csa_tree_add_22_22_n_343 ,csa_tree_add_22_22_n_207 ,csa_tree_add_22_22_n_303);
  and csa_tree_add_22_22_g3523__8428(csa_tree_add_22_22_n_342 ,csa_tree_add_22_22_n_232 ,csa_tree_add_22_22_n_311);
  and csa_tree_add_22_22_g3524__5526(csa_tree_add_22_22_n_341 ,csa_tree_add_22_22_n_234 ,csa_tree_add_22_22_n_310);
  and csa_tree_add_22_22_g3525__6783(csa_tree_add_22_22_n_340 ,csa_tree_add_22_22_n_238 ,csa_tree_add_22_22_n_304);
  and csa_tree_add_22_22_g3526__3680(csa_tree_add_22_22_n_339 ,csa_tree_add_22_22_n_220 ,csa_tree_add_22_22_n_306);
  and csa_tree_add_22_22_g3527__1617(csa_tree_add_22_22_n_338 ,csa_tree_add_22_22_n_210 ,csa_tree_add_22_22_n_300);
  and csa_tree_add_22_22_g3528__2802(csa_tree_add_22_22_n_336 ,csa_tree_add_22_22_n_230 ,csa_tree_add_22_22_n_307);
  and csa_tree_add_22_22_g3529__1705(csa_tree_add_22_22_n_334 ,csa_tree_add_22_22_n_237 ,csa_tree_add_22_22_n_302);
  and csa_tree_add_22_22_g3530__5122(csa_tree_add_22_22_n_333 ,csa_tree_add_22_22_n_211 ,csa_tree_add_22_22_n_301);
  and csa_tree_add_22_22_g3531__8246(csa_tree_add_22_22_n_332 ,csa_tree_add_22_22_n_216 ,csa_tree_add_22_22_n_305);
  and csa_tree_add_22_22_g3532__7098(csa_tree_add_22_22_n_331 ,csa_tree_add_22_22_n_242 ,csa_tree_add_22_22_n_308);
  and csa_tree_add_22_22_g3533__6131(csa_tree_add_22_22_n_330 ,csa_tree_add_22_22_n_205 ,csa_tree_add_22_22_n_299);
  and csa_tree_add_22_22_g3534__1881(csa_tree_add_22_22_n_329 ,csa_tree_add_22_22_n_227 ,csa_tree_add_22_22_n_309);
  not csa_tree_add_22_22_g3535(csa_tree_add_22_22_n_324 ,csa_tree_add_22_22_n_325);
  not csa_tree_add_22_22_g3536(csa_tree_add_22_22_n_321 ,csa_tree_add_22_22_n_320);
  not csa_tree_add_22_22_g3537(csa_tree_add_22_22_n_318 ,csa_tree_add_22_22_n_319);
  and csa_tree_add_22_22_g3538__5115(csa_tree_add_22_22_n_316 ,csa_tree_add_22_22_n_224 ,csa_tree_add_22_22_n_285);
  nor csa_tree_add_22_22_g3539__7482(csa_tree_add_22_22_n_315 ,csa_tree_add_22_22_n_252 ,csa_tree_add_22_22_n_283);
  and csa_tree_add_22_22_g3540__4733(csa_tree_add_22_22_n_314 ,csa_tree_add_22_22_n_296 ,csa_tree_add_22_22_n_284);
  and csa_tree_add_22_22_g3541__6161(csa_tree_add_22_22_n_313 ,csa_tree_add_22_22_n_252 ,csa_tree_add_22_22_n_283);
  xnor csa_tree_add_22_22_g3542__9315(csa_tree_add_22_22_n_312 ,csa_tree_add_22_22_n_173 ,csa_tree_add_22_22_n_253);
  and csa_tree_add_22_22_g3543__9945(csa_tree_add_22_22_n_327 ,csa_tree_add_22_22_n_217 ,csa_tree_add_22_22_n_288);
  and csa_tree_add_22_22_g3544__2883(csa_tree_add_22_22_n_326 ,csa_tree_add_22_22_n_235 ,csa_tree_add_22_22_n_292);
  and csa_tree_add_22_22_g3545__2346(csa_tree_add_22_22_n_325 ,csa_tree_add_22_22_n_223 ,csa_tree_add_22_22_n_291);
  and csa_tree_add_22_22_g3546__1666(csa_tree_add_22_22_n_323 ,csa_tree_add_22_22_n_221 ,csa_tree_add_22_22_n_290);
  and csa_tree_add_22_22_g3547__7410(csa_tree_add_22_22_n_322 ,csa_tree_add_22_22_n_239 ,csa_tree_add_22_22_n_289);
  or csa_tree_add_22_22_g3548__6417(csa_tree_add_22_22_n_320 ,csa_tree_add_22_22_n_247 ,csa_tree_add_22_22_n_287);
  and csa_tree_add_22_22_g3549__5477(csa_tree_add_22_22_n_319 ,csa_tree_add_22_22_n_219 ,csa_tree_add_22_22_n_293);
  and csa_tree_add_22_22_g3550__2398(csa_tree_add_22_22_n_317 ,csa_tree_add_22_22_n_244 ,csa_tree_add_22_22_n_294);
  or csa_tree_add_22_22_g3551__5107(csa_tree_add_22_22_n_311 ,csa_tree_add_22_22_n_199 ,csa_tree_add_22_22_n_233);
  or csa_tree_add_22_22_g3552__6260(csa_tree_add_22_22_n_310 ,csa_tree_add_22_22_n_156 ,csa_tree_add_22_22_n_249);
  or csa_tree_add_22_22_g3553__4319(csa_tree_add_22_22_n_309 ,csa_tree_add_22_22_n_194 ,csa_tree_add_22_22_n_208);
  or csa_tree_add_22_22_g3554__8428(csa_tree_add_22_22_n_308 ,csa_tree_add_22_22_n_160 ,csa_tree_add_22_22_n_240);
  or csa_tree_add_22_22_g3555__5526(csa_tree_add_22_22_n_307 ,csa_tree_add_22_22_n_164 ,csa_tree_add_22_22_n_215);
  or csa_tree_add_22_22_g3556__6783(csa_tree_add_22_22_n_306 ,csa_tree_add_22_22_n_189 ,csa_tree_add_22_22_n_213);
  or csa_tree_add_22_22_g3557__3680(csa_tree_add_22_22_n_305 ,csa_tree_add_22_22_n_192 ,csa_tree_add_22_22_n_214);
  or csa_tree_add_22_22_g3558__1617(csa_tree_add_22_22_n_304 ,csa_tree_add_22_22_n_161 ,csa_tree_add_22_22_n_251);
  or csa_tree_add_22_22_g3559__2802(csa_tree_add_22_22_n_303 ,csa_tree_add_22_22_n_198 ,csa_tree_add_22_22_n_209);
  or csa_tree_add_22_22_g3560__1705(csa_tree_add_22_22_n_302 ,csa_tree_add_22_22_n_204 ,csa_tree_add_22_22_n_245);
  or csa_tree_add_22_22_g3561__5122(csa_tree_add_22_22_n_301 ,csa_tree_add_22_22_n_158 ,csa_tree_add_22_22_n_228);
  or csa_tree_add_22_22_g3562__8246(csa_tree_add_22_22_n_300 ,csa_tree_add_22_22_n_203 ,csa_tree_add_22_22_n_212);
  or csa_tree_add_22_22_g3563__7098(csa_tree_add_22_22_n_299 ,csa_tree_add_22_22_n_159 ,csa_tree_add_22_22_n_218);
  or csa_tree_add_22_22_g3564__6131(csa_tree_add_22_22_n_298 ,csa_tree_add_22_22_n_173 ,csa_tree_add_22_22_n_253);
  nor csa_tree_add_22_22_g3565__1881(csa_tree_add_22_22_n_297 ,csa_tree_add_22_22_n_139 ,csa_tree_add_22_22_n_255);
  or csa_tree_add_22_22_g3566__5115(csa_tree_add_22_22_n_296 ,csa_tree_add_22_22_n_138 ,csa_tree_add_22_22_n_254);
  and csa_tree_add_22_22_g3567__7482(csa_tree_add_22_22_n_295 ,csa_tree_add_22_22_n_173 ,csa_tree_add_22_22_n_253);
  or csa_tree_add_22_22_g3568__4733(csa_tree_add_22_22_n_294 ,csa_tree_add_22_22_n_197 ,csa_tree_add_22_22_n_250);
  or csa_tree_add_22_22_g3569__6161(csa_tree_add_22_22_n_293 ,csa_tree_add_22_22_n_191 ,csa_tree_add_22_22_n_225);
  or csa_tree_add_22_22_g3570__9315(csa_tree_add_22_22_n_292 ,csa_tree_add_22_22_n_196 ,csa_tree_add_22_22_n_246);
  or csa_tree_add_22_22_g3571__9945(csa_tree_add_22_22_n_291 ,csa_tree_add_22_22_n_195 ,csa_tree_add_22_22_n_222);
  or csa_tree_add_22_22_g3572__2883(csa_tree_add_22_22_n_290 ,csa_tree_add_22_22_n_190 ,csa_tree_add_22_22_n_226);
  or csa_tree_add_22_22_g3573__2346(csa_tree_add_22_22_n_289 ,csa_tree_add_22_22_n_157 ,csa_tree_add_22_22_n_236);
  or csa_tree_add_22_22_g3574__1666(csa_tree_add_22_22_n_288 ,csa_tree_add_22_22_n_201 ,csa_tree_add_22_22_n_241);
  nor csa_tree_add_22_22_g3575__7410(csa_tree_add_22_22_n_287 ,csa_tree_add_22_22_n_165 ,csa_tree_add_22_22_n_248);
  xnor csa_tree_add_22_22_g3576__6417(n_613 ,csa_tree_add_22_22_n_166 ,in9[1]);
  not csa_tree_add_22_22_g3577(csa_tree_add_22_22_n_283 ,csa_tree_add_22_22_n_282);
  not csa_tree_add_22_22_g3578(csa_tree_add_22_22_n_280 ,csa_tree_add_22_22_n_281);
  xnor csa_tree_add_22_22_g3579__5477(csa_tree_add_22_22_n_279 ,csa_tree_add_22_22_n_165 ,in9[12]);
  xnor csa_tree_add_22_22_g3580__2398(csa_tree_add_22_22_n_278 ,csa_tree_add_22_22_n_175 ,in9[16]);
  xnor csa_tree_add_22_22_g3581__5107(csa_tree_add_22_22_n_277 ,csa_tree_add_22_22_n_177 ,csa_tree_add_22_22_n_158);
  xnor csa_tree_add_22_22_g3582__6260(csa_tree_add_22_22_n_276 ,csa_tree_add_22_22_n_204 ,in9[5]);
  xnor csa_tree_add_22_22_g3583__4319(csa_tree_add_22_22_n_275 ,csa_tree_add_22_22_n_199 ,in9[9]);
  xnor csa_tree_add_22_22_g3584__8428(csa_tree_add_22_22_n_274 ,csa_tree_add_22_22_n_160 ,in9[10]);
  xnor csa_tree_add_22_22_g3585__5526(csa_tree_add_22_22_n_273 ,csa_tree_add_22_22_n_156 ,in9[7]);
  xnor csa_tree_add_22_22_g3586__6783(csa_tree_add_22_22_n_272 ,csa_tree_add_22_22_n_197 ,in9[11]);
  xnor csa_tree_add_22_22_g3587__3680(csa_tree_add_22_22_n_271 ,csa_tree_add_22_22_n_157 ,in9[14]);
  xnor csa_tree_add_22_22_g3588__1617(csa_tree_add_22_22_n_270 ,csa_tree_add_22_22_n_196 ,in9[15]);
  xnor csa_tree_add_22_22_g3589__2802(csa_tree_add_22_22_n_269 ,csa_tree_add_22_22_n_161 ,in9[6]);
  xnor csa_tree_add_22_22_g3590__1705(csa_tree_add_22_22_n_268 ,csa_tree_add_22_22_n_201 ,in9[8]);
  xnor csa_tree_add_22_22_g3591__5122(csa_tree_add_22_22_n_267 ,csa_tree_add_22_22_n_172 ,csa_tree_add_22_22_n_149);
  xnor csa_tree_add_22_22_g3592__8246(csa_tree_add_22_22_n_266 ,csa_tree_add_22_22_n_154 ,csa_tree_add_22_22_n_164);
  xnor csa_tree_add_22_22_g3593__7098(csa_tree_add_22_22_n_265 ,csa_tree_add_22_22_n_153 ,csa_tree_add_22_22_n_137);
  xnor csa_tree_add_22_22_g3594__6131(csa_tree_add_22_22_n_264 ,csa_tree_add_22_22_n_126 ,csa_tree_add_22_22_n_198);
  xnor csa_tree_add_22_22_g3595__1881(csa_tree_add_22_22_n_263 ,csa_tree_add_22_22_n_144 ,csa_tree_add_22_22_n_152);
  xnor csa_tree_add_22_22_g3596__5115(csa_tree_add_22_22_n_262 ,csa_tree_add_22_22_n_136 ,csa_tree_add_22_22_n_188);
  xnor csa_tree_add_22_22_g3597__7482(csa_tree_add_22_22_n_261 ,csa_tree_add_22_22_n_180 ,csa_tree_add_22_22_n_195);
  xnor csa_tree_add_22_22_g3598__4733(csa_tree_add_22_22_n_260 ,csa_tree_add_22_22_n_184 ,csa_tree_add_22_22_n_194);
  xnor csa_tree_add_22_22_g3599__6161(csa_tree_add_22_22_n_259 ,csa_tree_add_22_22_n_130 ,csa_tree_add_22_22_n_190);
  xnor csa_tree_add_22_22_g3600__9315(csa_tree_add_22_22_n_258 ,csa_tree_add_22_22_n_181 ,csa_tree_add_22_22_n_203);
  xnor csa_tree_add_22_22_g3601__9945(csa_tree_add_22_22_n_257 ,csa_tree_add_22_22_n_127 ,csa_tree_add_22_22_n_192);
  xnor csa_tree_add_22_22_g3602__2883(csa_tree_add_22_22_n_285 ,csa_tree_add_22_22_n_200 ,in9[2]);
  xnor csa_tree_add_22_22_g3603__2346(csa_tree_add_22_22_n_284 ,csa_tree_add_22_22_n_193 ,in9[4]);
  xnor csa_tree_add_22_22_g3604__1666(csa_tree_add_22_22_n_282 ,csa_tree_add_22_22_n_162 ,in9[3]);
  xnor csa_tree_add_22_22_g3605__7410(csa_tree_add_22_22_n_281 ,csa_tree_add_22_22_n_202 ,in9[13]);
  not csa_tree_add_22_22_g3606(csa_tree_add_22_22_n_255 ,csa_tree_add_22_22_n_254);
  nor csa_tree_add_22_22_g3607__6417(csa_tree_add_22_22_n_251 ,in9[6] ,csa_tree_add_22_22_n_178);
  nor csa_tree_add_22_22_g3608__5477(csa_tree_add_22_22_n_250 ,in9[11] ,csa_tree_add_22_22_n_170);
  nor csa_tree_add_22_22_g3609__2398(csa_tree_add_22_22_n_249 ,in9[7] ,csa_tree_add_22_22_n_133);
  and csa_tree_add_22_22_g3610__5107(csa_tree_add_22_22_n_248 ,csa_tree_add_22_22_n_121 ,csa_tree_add_22_22_n_129);
  nor csa_tree_add_22_22_g3611__6260(csa_tree_add_22_22_n_247 ,csa_tree_add_22_22_n_121 ,csa_tree_add_22_22_n_129);
  nor csa_tree_add_22_22_g3612__4319(csa_tree_add_22_22_n_246 ,in9[15] ,csa_tree_add_22_22_n_185);
  nor csa_tree_add_22_22_g3613__8428(csa_tree_add_22_22_n_245 ,in9[5] ,csa_tree_add_22_22_n_145);
  or csa_tree_add_22_22_g3614__5526(csa_tree_add_22_22_n_244 ,csa_tree_add_22_22_n_123 ,csa_tree_add_22_22_n_171);
  nor csa_tree_add_22_22_g3615__6783(csa_tree_add_22_22_n_243 ,csa_tree_add_22_22_n_120 ,csa_tree_add_22_22_n_175);
  or csa_tree_add_22_22_g3616__3680(csa_tree_add_22_22_n_242 ,csa_tree_add_22_22_n_122 ,csa_tree_add_22_22_n_183);
  nor csa_tree_add_22_22_g3617__1617(csa_tree_add_22_22_n_241 ,in9[8] ,csa_tree_add_22_22_n_150);
  nor csa_tree_add_22_22_g3618__2802(csa_tree_add_22_22_n_240 ,in9[10] ,csa_tree_add_22_22_n_182);
  or csa_tree_add_22_22_g3619__1705(csa_tree_add_22_22_n_239 ,csa_tree_add_22_22_n_124 ,csa_tree_add_22_22_n_148);
  or csa_tree_add_22_22_g3620__5122(csa_tree_add_22_22_n_238 ,csa_tree_add_22_22_n_104 ,csa_tree_add_22_22_n_179);
  or csa_tree_add_22_22_g3621__8246(csa_tree_add_22_22_n_237 ,csa_tree_add_22_22_n_108 ,csa_tree_add_22_22_n_146);
  nor csa_tree_add_22_22_g3622__7098(csa_tree_add_22_22_n_236 ,in9[14] ,csa_tree_add_22_22_n_147);
  or csa_tree_add_22_22_g3623__6131(csa_tree_add_22_22_n_235 ,csa_tree_add_22_22_n_107 ,csa_tree_add_22_22_n_186);
  or csa_tree_add_22_22_g3624__1881(csa_tree_add_22_22_n_234 ,csa_tree_add_22_22_n_119 ,csa_tree_add_22_22_n_134);
  nor csa_tree_add_22_22_g3625__5115(csa_tree_add_22_22_n_233 ,in9[9] ,csa_tree_add_22_22_n_141);
  or csa_tree_add_22_22_g3626__7482(csa_tree_add_22_22_n_232 ,csa_tree_add_22_22_n_106 ,csa_tree_add_22_22_n_142);
  and csa_tree_add_22_22_g3627__4733(n_484 ,in9[1] ,csa_tree_add_22_22_n_167);
  or csa_tree_add_22_22_g3628__6161(csa_tree_add_22_22_n_256 ,csa_tree_add_22_22_n_125 ,csa_tree_add_22_22_n_193);
  and csa_tree_add_22_22_g3629__9315(csa_tree_add_22_22_n_254 ,in9[3] ,csa_tree_add_22_22_n_163);
  or csa_tree_add_22_22_g3630__9945(csa_tree_add_22_22_n_253 ,csa_tree_add_22_22_n_110 ,csa_tree_add_22_22_n_202);
  or csa_tree_add_22_22_g3631__2883(csa_tree_add_22_22_n_252 ,csa_tree_add_22_22_n_109 ,csa_tree_add_22_22_n_200);
  or csa_tree_add_22_22_g3632__2346(csa_tree_add_22_22_n_230 ,csa_tree_add_22_22_n_155 ,csa_tree_add_22_22_n_154);
  and csa_tree_add_22_22_g3633__1666(csa_tree_add_22_22_n_229 ,csa_tree_add_22_22_n_120 ,csa_tree_add_22_22_n_175);
  and csa_tree_add_22_22_g3634__7410(csa_tree_add_22_22_n_228 ,csa_tree_add_22_22_n_128 ,csa_tree_add_22_22_n_177);
  or csa_tree_add_22_22_g3635__6417(csa_tree_add_22_22_n_227 ,csa_tree_add_22_22_n_132 ,csa_tree_add_22_22_n_184);
  and csa_tree_add_22_22_g3636__5477(csa_tree_add_22_22_n_226 ,csa_tree_add_22_22_n_143 ,csa_tree_add_22_22_n_130);
  and csa_tree_add_22_22_g3637__2398(csa_tree_add_22_22_n_225 ,csa_tree_add_22_22_n_153 ,csa_tree_add_22_22_n_137);
  or csa_tree_add_22_22_g3638__5107(csa_tree_add_22_22_n_224 ,csa_tree_add_22_22_n_135 ,csa_tree_add_22_22_n_187);
  or csa_tree_add_22_22_g3639__6260(csa_tree_add_22_22_n_223 ,csa_tree_add_22_22_n_176 ,csa_tree_add_22_22_n_180);
  and csa_tree_add_22_22_g3640__4319(csa_tree_add_22_22_n_222 ,csa_tree_add_22_22_n_176 ,csa_tree_add_22_22_n_180);
  or csa_tree_add_22_22_g3641__8428(csa_tree_add_22_22_n_221 ,csa_tree_add_22_22_n_143 ,csa_tree_add_22_22_n_130);
  or csa_tree_add_22_22_g3642__5526(csa_tree_add_22_22_n_220 ,csa_tree_add_22_22_n_172 ,csa_tree_add_22_22_n_149);
  or csa_tree_add_22_22_g3643__6783(csa_tree_add_22_22_n_219 ,csa_tree_add_22_22_n_153 ,csa_tree_add_22_22_n_137);
  and csa_tree_add_22_22_g3644__3680(csa_tree_add_22_22_n_218 ,csa_tree_add_22_22_n_144 ,csa_tree_add_22_22_n_152);
  or csa_tree_add_22_22_g3645__1617(csa_tree_add_22_22_n_217 ,csa_tree_add_22_22_n_105 ,csa_tree_add_22_22_n_151);
  or csa_tree_add_22_22_g3646__2802(csa_tree_add_22_22_n_216 ,csa_tree_add_22_22_n_174 ,csa_tree_add_22_22_n_127);
  and csa_tree_add_22_22_g3647__1705(csa_tree_add_22_22_n_215 ,csa_tree_add_22_22_n_155 ,csa_tree_add_22_22_n_154);
  and csa_tree_add_22_22_g3648__5122(csa_tree_add_22_22_n_214 ,csa_tree_add_22_22_n_174 ,csa_tree_add_22_22_n_127);
  and csa_tree_add_22_22_g3649__8246(csa_tree_add_22_22_n_213 ,csa_tree_add_22_22_n_172 ,csa_tree_add_22_22_n_149);
  and csa_tree_add_22_22_g3650__7098(csa_tree_add_22_22_n_212 ,csa_tree_add_22_22_n_140 ,csa_tree_add_22_22_n_181);
  or csa_tree_add_22_22_g3651__6131(csa_tree_add_22_22_n_211 ,csa_tree_add_22_22_n_128 ,csa_tree_add_22_22_n_177);
  or csa_tree_add_22_22_g3652__1881(csa_tree_add_22_22_n_210 ,csa_tree_add_22_22_n_140 ,csa_tree_add_22_22_n_181);
  and csa_tree_add_22_22_g3653__5115(csa_tree_add_22_22_n_209 ,csa_tree_add_22_22_n_131 ,csa_tree_add_22_22_n_126);
  and csa_tree_add_22_22_g3654__7482(csa_tree_add_22_22_n_208 ,csa_tree_add_22_22_n_132 ,csa_tree_add_22_22_n_184);
  or csa_tree_add_22_22_g3655__4733(csa_tree_add_22_22_n_207 ,csa_tree_add_22_22_n_131 ,csa_tree_add_22_22_n_126);
  nor csa_tree_add_22_22_g3656__6161(csa_tree_add_22_22_n_206 ,csa_tree_add_22_22_n_136 ,csa_tree_add_22_22_n_188);
  or csa_tree_add_22_22_g3657__9315(csa_tree_add_22_22_n_205 ,csa_tree_add_22_22_n_144 ,csa_tree_add_22_22_n_152);
  not csa_tree_add_22_22_g3658(csa_tree_add_22_22_n_187 ,csa_tree_add_22_22_n_188);
  not csa_tree_add_22_22_g3659(csa_tree_add_22_22_n_185 ,csa_tree_add_22_22_n_186);
  not csa_tree_add_22_22_g3660(csa_tree_add_22_22_n_182 ,csa_tree_add_22_22_n_183);
  not csa_tree_add_22_22_g3661(csa_tree_add_22_22_n_178 ,csa_tree_add_22_22_n_179);
  not csa_tree_add_22_22_g3662(csa_tree_add_22_22_n_170 ,csa_tree_add_22_22_n_171);
  and csa_tree_add_22_22_g3663__9945(n_614 ,in1[0] ,in10[0]);
  and csa_tree_add_22_22_g3664__2883(n_485 ,in1[1] ,in10[0]);
  or csa_tree_add_22_22_g3665__2346(csa_tree_add_22_22_n_204 ,csa_tree_add_22_22_n_90 ,csa_tree_add_22_22_n_33);
  or csa_tree_add_22_22_g3666__1666(csa_tree_add_22_22_n_203 ,csa_tree_add_22_22_n_51 ,csa_tree_add_22_22_n_9);
  or csa_tree_add_22_22_g3667__7410(csa_tree_add_22_22_n_202 ,csa_tree_add_22_22_n_60 ,csa_tree_add_22_22_n_80);
  or csa_tree_add_22_22_g3668__6417(csa_tree_add_22_22_n_201 ,csa_tree_add_22_22_n_98 ,csa_tree_add_22_22_n_71);
  or csa_tree_add_22_22_g3669__5477(csa_tree_add_22_22_n_200 ,csa_tree_add_22_22_n_63 ,csa_tree_add_22_22_n_28);
  or csa_tree_add_22_22_g3670__2398(csa_tree_add_22_22_n_199 ,csa_tree_add_22_22_n_54 ,csa_tree_add_22_22_n_71);
  or csa_tree_add_22_22_g3671__5107(csa_tree_add_22_22_n_198 ,csa_tree_add_22_22_n_57 ,csa_tree_add_22_22_n_2);
  or csa_tree_add_22_22_g3672__6260(csa_tree_add_22_22_n_197 ,csa_tree_add_22_22_n_118 ,csa_tree_add_22_22_n_71);
  or csa_tree_add_22_22_g3673__4319(csa_tree_add_22_22_n_196 ,csa_tree_add_22_22_n_117 ,csa_tree_add_22_22_n_13);
  or csa_tree_add_22_22_g3674__8428(csa_tree_add_22_22_n_195 ,csa_tree_add_22_22_n_88 ,csa_tree_add_22_22_n_9);
  or csa_tree_add_22_22_g3675__5526(csa_tree_add_22_22_n_194 ,csa_tree_add_22_22_n_84 ,csa_tree_add_22_22_n_80);
  or csa_tree_add_22_22_g3676__6783(csa_tree_add_22_22_n_193 ,csa_tree_add_22_22_n_48 ,csa_tree_add_22_22_n_28);
  or csa_tree_add_22_22_g3677__3680(csa_tree_add_22_22_n_192 ,csa_tree_add_22_22_n_103 ,csa_tree_add_22_22_n_80);
  or csa_tree_add_22_22_g3678__1617(csa_tree_add_22_22_n_191 ,csa_tree_add_22_22_n_116 ,csa_tree_add_22_22_n_1);
  or csa_tree_add_22_22_g3679__2802(csa_tree_add_22_22_n_190 ,csa_tree_add_22_22_n_92 ,csa_tree_add_22_22_n_80);
  or csa_tree_add_22_22_g3680__1705(csa_tree_add_22_22_n_189 ,csa_tree_add_22_22_n_57 ,csa_tree_add_22_22_n_36);
  or csa_tree_add_22_22_g3681__5122(csa_tree_add_22_22_n_188 ,csa_tree_add_22_22_n_82 ,csa_tree_add_22_22_n_80);
  or csa_tree_add_22_22_g3682__8246(csa_tree_add_22_22_n_186 ,csa_tree_add_22_22_n_118 ,csa_tree_add_22_22_n_74);
  or csa_tree_add_22_22_g3683__7098(csa_tree_add_22_22_n_184 ,csa_tree_add_22_22_n_97 ,csa_tree_add_22_22_n_77);
  or csa_tree_add_22_22_g3684__6131(csa_tree_add_22_22_n_183 ,csa_tree_add_22_22_n_51 ,csa_tree_add_22_22_n_4);
  or csa_tree_add_22_22_g3685__1881(csa_tree_add_22_22_n_181 ,csa_tree_add_22_22_n_84 ,csa_tree_add_22_22_n_7);
  or csa_tree_add_22_22_g3686__5115(csa_tree_add_22_22_n_180 ,csa_tree_add_22_22_n_90 ,csa_tree_add_22_22_n_13);
  or csa_tree_add_22_22_g3687__7482(csa_tree_add_22_22_n_179 ,csa_tree_add_22_22_n_48 ,csa_tree_add_22_22_n_68);
  or csa_tree_add_22_22_g3688__4733(csa_tree_add_22_22_n_177 ,csa_tree_add_22_22_n_63 ,csa_tree_add_22_22_n_77);
  or csa_tree_add_22_22_g3689__6161(csa_tree_add_22_22_n_176 ,csa_tree_add_22_22_n_97 ,csa_tree_add_22_22_n_23);
  or csa_tree_add_22_22_g3690__9315(csa_tree_add_22_22_n_175 ,csa_tree_add_22_22_n_60 ,csa_tree_add_22_22_n_23);
  or csa_tree_add_22_22_g3691__9945(csa_tree_add_22_22_n_174 ,csa_tree_add_22_22_n_96 ,csa_tree_add_22_22_n_18);
  or csa_tree_add_22_22_g3692__2883(csa_tree_add_22_22_n_173 ,csa_tree_add_22_22_n_57 ,csa_tree_add_22_22_n_77);
  or csa_tree_add_22_22_g3693__2346(csa_tree_add_22_22_n_172 ,csa_tree_add_22_22_n_54 ,csa_tree_add_22_22_n_74);
  or csa_tree_add_22_22_g3694__1666(csa_tree_add_22_22_n_171 ,csa_tree_add_22_22_n_103 ,csa_tree_add_22_22_n_68);
  not csa_tree_add_22_22_g3695(csa_tree_add_22_22_n_167 ,csa_tree_add_22_22_n_166);
  not csa_tree_add_22_22_g3696(csa_tree_add_22_22_n_163 ,csa_tree_add_22_22_n_162);
  not csa_tree_add_22_22_g3697(csa_tree_add_22_22_n_151 ,csa_tree_add_22_22_n_150);
  not csa_tree_add_22_22_g3698(csa_tree_add_22_22_n_148 ,csa_tree_add_22_22_n_147);
  not csa_tree_add_22_22_g3699(csa_tree_add_22_22_n_145 ,csa_tree_add_22_22_n_146);
  not csa_tree_add_22_22_g3700(csa_tree_add_22_22_n_142 ,csa_tree_add_22_22_n_141);
  not csa_tree_add_22_22_g3701(csa_tree_add_22_22_n_138 ,csa_tree_add_22_22_n_139);
  not csa_tree_add_22_22_g3702(csa_tree_add_22_22_n_135 ,csa_tree_add_22_22_n_136);
  not csa_tree_add_22_22_g3703(csa_tree_add_22_22_n_134 ,csa_tree_add_22_22_n_133);
  or csa_tree_add_22_22_g3704__7410(csa_tree_add_22_22_n_166 ,csa_tree_add_22_22_n_86 ,csa_tree_add_22_22_n_9);
  or csa_tree_add_22_22_g3705__6417(csa_tree_add_22_22_n_165 ,csa_tree_add_22_22_n_117 ,csa_tree_add_22_22_n_27);
  or csa_tree_add_22_22_g3706__5477(csa_tree_add_22_22_n_164 ,csa_tree_add_22_22_n_114 ,csa_tree_add_22_22_n_2);
  or csa_tree_add_22_22_g3707__2398(csa_tree_add_22_22_n_162 ,csa_tree_add_22_22_n_45 ,csa_tree_add_22_22_n_71);
  or csa_tree_add_22_22_g3708__5107(csa_tree_add_22_22_n_161 ,csa_tree_add_22_22_n_96 ,csa_tree_add_22_22_n_71);
  or csa_tree_add_22_22_g3709__6260(csa_tree_add_22_22_n_160 ,csa_tree_add_22_22_n_92 ,csa_tree_add_22_22_n_71);
  or csa_tree_add_22_22_g3710__4319(csa_tree_add_22_22_n_159 ,csa_tree_add_22_22_n_102 ,csa_tree_add_22_22_n_9);
  or csa_tree_add_22_22_g3711__8428(csa_tree_add_22_22_n_158 ,csa_tree_add_22_22_n_48 ,csa_tree_add_22_22_n_80);
  or csa_tree_add_22_22_g3712__5526(csa_tree_add_22_22_n_157 ,csa_tree_add_22_22_n_60 ,csa_tree_add_22_22_n_4);
  or csa_tree_add_22_22_g3713__6783(csa_tree_add_22_22_n_156 ,csa_tree_add_22_22_n_88 ,csa_tree_add_22_22_n_33);
  or csa_tree_add_22_22_g3714__3680(csa_tree_add_22_22_n_155 ,csa_tree_add_22_22_n_116 ,csa_tree_add_22_22_n_18);
  or csa_tree_add_22_22_g3715__1617(csa_tree_add_22_22_n_154 ,csa_tree_add_22_22_n_45 ,csa_tree_add_22_22_n_6);
  or csa_tree_add_22_22_g3716__2802(csa_tree_add_22_22_n_153 ,csa_tree_add_22_22_n_86 ,csa_tree_add_22_22_n_77);
  or csa_tree_add_22_22_g3717__1705(csa_tree_add_22_22_n_152 ,csa_tree_add_22_22_n_63 ,csa_tree_add_22_22_n_36);
  and csa_tree_add_22_22_g3718__5122(csa_tree_add_22_22_n_150 ,in1[6] ,in10[2]);
  or csa_tree_add_22_22_g3719__8246(csa_tree_add_22_22_n_149 ,csa_tree_add_22_22_n_115 ,csa_tree_add_22_22_n_77);
  and csa_tree_add_22_22_g3720__7098(csa_tree_add_22_22_n_147 ,in1[10] ,in10[4]);
  or csa_tree_add_22_22_g3721__6131(csa_tree_add_22_22_n_146 ,csa_tree_add_22_22_n_102 ,csa_tree_add_22_22_n_68);
  or csa_tree_add_22_22_g3722__1881(csa_tree_add_22_22_n_144 ,csa_tree_add_22_22_n_82 ,csa_tree_add_22_22_n_13);
  or csa_tree_add_22_22_g3723__5115(csa_tree_add_22_22_n_143 ,csa_tree_add_22_22_n_100 ,csa_tree_add_22_22_n_74);
  and csa_tree_add_22_22_g3724__7482(csa_tree_add_22_22_n_141 ,in1[7] ,in10[2]);
  or csa_tree_add_22_22_g3725__4733(csa_tree_add_22_22_n_140 ,csa_tree_add_22_22_n_114 ,csa_tree_add_22_22_n_17);
  or csa_tree_add_22_22_g3726__6161(csa_tree_add_22_22_n_139 ,csa_tree_add_22_22_n_99 ,csa_tree_add_22_22_n_23);
  or csa_tree_add_22_22_g3727__9315(csa_tree_add_22_22_n_137 ,csa_tree_add_22_22_n_101 ,csa_tree_add_22_22_n_68);
  or csa_tree_add_22_22_g3728__9945(csa_tree_add_22_22_n_136 ,csa_tree_add_22_22_n_99 ,csa_tree_add_22_22_n_68);
  and csa_tree_add_22_22_g3729__2883(csa_tree_add_22_22_n_133 ,in1[5] ,in10[2]);
  or csa_tree_add_22_22_g3730__2346(csa_tree_add_22_22_n_132 ,csa_tree_add_22_22_n_45 ,csa_tree_add_22_22_n_74);
  or csa_tree_add_22_22_g3731__1666(csa_tree_add_22_22_n_131 ,csa_tree_add_22_22_n_98 ,csa_tree_add_22_22_n_23);
  or csa_tree_add_22_22_g3732__7410(csa_tree_add_22_22_n_130 ,csa_tree_add_22_22_n_51 ,csa_tree_add_22_22_n_7);
  or csa_tree_add_22_22_g3733__6417(csa_tree_add_22_22_n_129 ,csa_tree_add_22_22_n_115 ,csa_tree_add_22_22_n_35);
  or csa_tree_add_22_22_g3734__5477(csa_tree_add_22_22_n_128 ,csa_tree_add_22_22_n_101 ,csa_tree_add_22_22_n_74);
  or csa_tree_add_22_22_g3735__2398(csa_tree_add_22_22_n_127 ,csa_tree_add_22_22_n_100 ,csa_tree_add_22_22_n_13);
  or csa_tree_add_22_22_g3736__5107(csa_tree_add_22_22_n_126 ,csa_tree_add_22_22_n_54 ,csa_tree_add_22_22_n_77);
  not csa_tree_add_22_22_g3737(csa_tree_add_22_22_n_125 ,in9[4]);
  not csa_tree_add_22_22_g3738(csa_tree_add_22_22_n_124 ,in9[14]);
  not csa_tree_add_22_22_g3739(csa_tree_add_22_22_n_123 ,in9[11]);
  not csa_tree_add_22_22_g3740(csa_tree_add_22_22_n_122 ,in9[10]);
  not csa_tree_add_22_22_g3741(csa_tree_add_22_22_n_121 ,in9[12]);
  not csa_tree_add_22_22_g3742(csa_tree_add_22_22_n_120 ,in9[16]);
  not csa_tree_add_22_22_g3743(csa_tree_add_22_22_n_119 ,in9[7]);
  not csa_tree_add_22_22_g3744(csa_tree_add_22_22_n_118 ,in1[11]);
  not csa_tree_add_22_22_g3745(csa_tree_add_22_22_n_117 ,in1[12]);
  not csa_tree_add_22_22_g3746(csa_tree_add_22_22_n_116 ,in1[2]);
  not csa_tree_add_22_22_g3747(csa_tree_add_22_22_n_115 ,in1[10]);
  not csa_tree_add_22_22_g3748(csa_tree_add_22_22_n_114 ,in1[5]);
  not csa_tree_add_22_22_g3749(csa_tree_add_22_22_n_113 ,in10[1]);
  not csa_tree_add_22_22_g3750(csa_tree_add_22_22_n_112 ,in10[3]);
  not csa_tree_add_22_22_g3751(csa_tree_add_22_22_n_111 ,in10[4]);
  not csa_tree_add_22_22_g3752(csa_tree_add_22_22_n_110 ,in9[13]);
  not csa_tree_add_22_22_g3753(csa_tree_add_22_22_n_109 ,in9[2]);
  not csa_tree_add_22_22_g3754(csa_tree_add_22_22_n_108 ,in9[5]);
  not csa_tree_add_22_22_g3755(csa_tree_add_22_22_n_107 ,in9[15]);
  not csa_tree_add_22_22_g3756(csa_tree_add_22_22_n_106 ,in9[9]);
  not csa_tree_add_22_22_g3757(csa_tree_add_22_22_n_105 ,in9[8]);
  not csa_tree_add_22_22_g3758(csa_tree_add_22_22_n_104 ,in9[6]);
  not csa_tree_add_22_22_g3759(csa_tree_add_22_22_n_103 ,in1[9]);
  not csa_tree_add_22_22_g3760(csa_tree_add_22_22_n_102 ,in1[3]);
  not csa_tree_add_22_22_g3761(csa_tree_add_22_22_n_101 ,in1[1]);
  not csa_tree_add_22_22_g3762(csa_tree_add_22_22_n_100 ,in1[7]);
  not csa_tree_add_22_22_g3763(csa_tree_add_22_22_n_99 ,in1[0]);
  not csa_tree_add_22_22_g3764(csa_tree_add_22_22_n_98 ,in1[8]);
  not csa_tree_add_22_22_g3765(csa_tree_add_22_22_n_97 ,in1[4]);
  not csa_tree_add_22_22_g3766(csa_tree_add_22_22_n_96 ,in1[6]);
  not csa_tree_add_22_22_g3767(csa_tree_add_22_22_n_95 ,in10[2]);
  not csa_tree_add_22_22_g3768(csa_tree_add_22_22_n_94 ,in10[0]);
  not csa_tree_add_22_22_drc_bufs3825(csa_tree_add_22_22_n_92 ,csa_tree_add_22_22_n_91);
  not csa_tree_add_22_22_drc_bufs3826(csa_tree_add_22_22_n_91 ,csa_tree_add_22_22_n_115);
  not csa_tree_add_22_22_drc_bufs3829(csa_tree_add_22_22_n_90 ,csa_tree_add_22_22_n_89);
  not csa_tree_add_22_22_drc_bufs3830(csa_tree_add_22_22_n_89 ,csa_tree_add_22_22_n_114);
  not csa_tree_add_22_22_drc_bufs3833(csa_tree_add_22_22_n_88 ,csa_tree_add_22_22_n_87);
  not csa_tree_add_22_22_drc_bufs3834(csa_tree_add_22_22_n_87 ,csa_tree_add_22_22_n_100);
  not csa_tree_add_22_22_drc_bufs3837(csa_tree_add_22_22_n_86 ,csa_tree_add_22_22_n_85);
  not csa_tree_add_22_22_drc_bufs3838(csa_tree_add_22_22_n_85 ,csa_tree_add_22_22_n_99);
  not csa_tree_add_22_22_drc_bufs3841(csa_tree_add_22_22_n_84 ,csa_tree_add_22_22_n_83);
  not csa_tree_add_22_22_drc_bufs3842(csa_tree_add_22_22_n_83 ,csa_tree_add_22_22_n_96);
  not csa_tree_add_22_22_drc_bufs3845(csa_tree_add_22_22_n_82 ,csa_tree_add_22_22_n_81);
  not csa_tree_add_22_22_drc_bufs3846(csa_tree_add_22_22_n_81 ,csa_tree_add_22_22_n_101);
  not csa_tree_add_22_22_drc_bufs3856(csa_tree_add_22_22_n_80 ,csa_tree_add_22_22_n_78);
  not csa_tree_add_22_22_drc_bufs3858(csa_tree_add_22_22_n_78 ,csa_tree_add_22_22_n_113);
  not csa_tree_add_22_22_drc_bufs3860(csa_tree_add_22_22_n_77 ,csa_tree_add_22_22_n_75);
  not csa_tree_add_22_22_drc_bufs3862(csa_tree_add_22_22_n_75 ,csa_tree_add_22_22_n_112);
  not csa_tree_add_22_22_drc_bufs3868(csa_tree_add_22_22_n_74 ,csa_tree_add_22_22_n_72);
  not csa_tree_add_22_22_drc_bufs3870(csa_tree_add_22_22_n_72 ,csa_tree_add_22_22_n_111);
  not csa_tree_add_22_22_drc_bufs3876(csa_tree_add_22_22_n_71 ,csa_tree_add_22_22_n_69);
  not csa_tree_add_22_22_drc_bufs3878(csa_tree_add_22_22_n_69 ,csa_tree_add_22_22_n_94);
  not csa_tree_add_22_22_drc_bufs3881(csa_tree_add_22_22_n_68 ,csa_tree_add_22_22_n_67);
  not csa_tree_add_22_22_drc_bufs3882(csa_tree_add_22_22_n_67 ,csa_tree_add_22_22_n_95);
  not csa_tree_add_22_22_drc_bufs3888(csa_tree_add_22_22_n_63 ,csa_tree_add_22_22_n_61);
  not csa_tree_add_22_22_drc_bufs3890(csa_tree_add_22_22_n_61 ,csa_tree_add_22_22_n_116);
  not csa_tree_add_22_22_drc_bufs3892(csa_tree_add_22_22_n_60 ,csa_tree_add_22_22_n_58);
  not csa_tree_add_22_22_drc_bufs3894(csa_tree_add_22_22_n_58 ,csa_tree_add_22_22_n_117);
  not csa_tree_add_22_22_drc_bufs3896(csa_tree_add_22_22_n_57 ,csa_tree_add_22_22_n_55);
  not csa_tree_add_22_22_drc_bufs3898(csa_tree_add_22_22_n_55 ,csa_tree_add_22_22_n_118);
  not csa_tree_add_22_22_drc_bufs3900(csa_tree_add_22_22_n_54 ,csa_tree_add_22_22_n_52);
  not csa_tree_add_22_22_drc_bufs3902(csa_tree_add_22_22_n_52 ,csa_tree_add_22_22_n_103);
  not csa_tree_add_22_22_drc_bufs3904(csa_tree_add_22_22_n_51 ,csa_tree_add_22_22_n_49);
  not csa_tree_add_22_22_drc_bufs3906(csa_tree_add_22_22_n_49 ,csa_tree_add_22_22_n_98);
  not csa_tree_add_22_22_drc_bufs3908(csa_tree_add_22_22_n_48 ,csa_tree_add_22_22_n_46);
  not csa_tree_add_22_22_drc_bufs3910(csa_tree_add_22_22_n_46 ,csa_tree_add_22_22_n_97);
  not csa_tree_add_22_22_drc_bufs3912(csa_tree_add_22_22_n_45 ,csa_tree_add_22_22_n_43);
  not csa_tree_add_22_22_drc_bufs3914(csa_tree_add_22_22_n_43 ,csa_tree_add_22_22_n_102);
  not csa_tree_add_22_22_drc_bufs3924(csa_tree_add_22_22_n_36 ,csa_tree_add_22_22_n_34);
  not csa_tree_add_22_22_drc_bufs3925(csa_tree_add_22_22_n_35 ,csa_tree_add_22_22_n_34);
  not csa_tree_add_22_22_drc_bufs3926(csa_tree_add_22_22_n_34 ,csa_tree_add_22_22_n_95);
  not csa_tree_add_22_22_drc_bufs3928(csa_tree_add_22_22_n_33 ,csa_tree_add_22_22_n_32);
  not csa_tree_add_22_22_drc_bufs3930(csa_tree_add_22_22_n_32 ,csa_tree_add_22_22_n_71);
  not csa_tree_add_22_22_drc_bufs3936(csa_tree_add_22_22_n_28 ,csa_tree_add_22_22_n_26);
  not csa_tree_add_22_22_drc_bufs3937(csa_tree_add_22_22_n_27 ,csa_tree_add_22_22_n_26);
  not csa_tree_add_22_22_drc_bufs3938(csa_tree_add_22_22_n_26 ,csa_tree_add_22_22_n_94);
  not csa_tree_add_22_22_drc_bufs3944(csa_tree_add_22_22_n_23 ,csa_tree_add_22_22_n_22);
  not csa_tree_add_22_22_drc_bufs3946(csa_tree_add_22_22_n_22 ,csa_tree_add_22_22_n_74);
  not csa_tree_add_22_22_drc_bufs3952(csa_tree_add_22_22_n_18 ,csa_tree_add_22_22_n_16);
  not csa_tree_add_22_22_drc_bufs3953(csa_tree_add_22_22_n_17 ,csa_tree_add_22_22_n_16);
  not csa_tree_add_22_22_drc_bufs3954(csa_tree_add_22_22_n_16 ,csa_tree_add_22_22_n_111);
  not csa_tree_add_22_22_drc_bufs3960(csa_tree_add_22_22_n_13 ,csa_tree_add_22_22_n_12);
  not csa_tree_add_22_22_drc_bufs3962(csa_tree_add_22_22_n_12 ,csa_tree_add_22_22_n_77);
  not csa_tree_add_22_22_drc_bufs3968(csa_tree_add_22_22_n_9 ,csa_tree_add_22_22_n_8);
  not csa_tree_add_22_22_drc_bufs3970(csa_tree_add_22_22_n_8 ,csa_tree_add_22_22_n_80);
  not csa_tree_add_22_22_drc_bufs3972(csa_tree_add_22_22_n_7 ,csa_tree_add_22_22_n_5);
  not csa_tree_add_22_22_drc_bufs3973(csa_tree_add_22_22_n_6 ,csa_tree_add_22_22_n_5);
  not csa_tree_add_22_22_drc_bufs3974(csa_tree_add_22_22_n_5 ,csa_tree_add_22_22_n_112);
  not csa_tree_add_22_22_drc_bufs3976(csa_tree_add_22_22_n_4 ,csa_tree_add_22_22_n_3);
  not csa_tree_add_22_22_drc_bufs3978(csa_tree_add_22_22_n_3 ,csa_tree_add_22_22_n_68);
  not csa_tree_add_22_22_drc_bufs3980(csa_tree_add_22_22_n_2 ,csa_tree_add_22_22_n_0);
  not csa_tree_add_22_22_drc_bufs3981(csa_tree_add_22_22_n_1 ,csa_tree_add_22_22_n_0);
  not csa_tree_add_22_22_drc_bufs3982(csa_tree_add_22_22_n_0 ,csa_tree_add_22_22_n_113);
  xnor csa_tree_add_24_21_groupi_g5525__6260(out1[32] ,csa_tree_add_24_21_groupi_n_2027 ,csa_tree_add_24_21_groupi_n_376);
  nor csa_tree_add_24_21_groupi_g5526__4319(csa_tree_add_24_21_groupi_n_2027 ,csa_tree_add_24_21_groupi_n_1457 ,csa_tree_add_24_21_groupi_n_2025);
  xnor csa_tree_add_24_21_groupi_g5527__8428(csa_tree_add_24_21_groupi_n_2026 ,csa_tree_add_24_21_groupi_n_2024 ,csa_tree_add_24_21_groupi_n_1527);
  nor csa_tree_add_24_21_groupi_g5528__5526(csa_tree_add_24_21_groupi_n_2025 ,csa_tree_add_24_21_groupi_n_1487 ,csa_tree_add_24_21_groupi_n_2024);
  and csa_tree_add_24_21_groupi_g5529__6783(csa_tree_add_24_21_groupi_n_2024 ,csa_tree_add_24_21_groupi_n_1536 ,csa_tree_add_24_21_groupi_n_2022);
  xnor csa_tree_add_24_21_groupi_g5530__3680(csa_tree_add_24_21_groupi_n_2023 ,csa_tree_add_24_21_groupi_n_2021 ,csa_tree_add_24_21_groupi_n_1588);
  or csa_tree_add_24_21_groupi_g5531__1617(csa_tree_add_24_21_groupi_n_2022 ,csa_tree_add_24_21_groupi_n_1534 ,csa_tree_add_24_21_groupi_n_2021);
  and csa_tree_add_24_21_groupi_g5532__2802(csa_tree_add_24_21_groupi_n_2021 ,csa_tree_add_24_21_groupi_n_1680 ,csa_tree_add_24_21_groupi_n_2019);
  xnor csa_tree_add_24_21_groupi_g5533__1705(csa_tree_add_24_21_groupi_n_2020 ,csa_tree_add_24_21_groupi_n_2018 ,csa_tree_add_24_21_groupi_n_1704);
  or csa_tree_add_24_21_groupi_g5534__5122(csa_tree_add_24_21_groupi_n_2019 ,csa_tree_add_24_21_groupi_n_1681 ,csa_tree_add_24_21_groupi_n_2018);
  and csa_tree_add_24_21_groupi_g5535__8246(csa_tree_add_24_21_groupi_n_2018 ,csa_tree_add_24_21_groupi_n_1717 ,csa_tree_add_24_21_groupi_n_2016);
  xnor csa_tree_add_24_21_groupi_g5536__7098(csa_tree_add_24_21_groupi_n_2017 ,csa_tree_add_24_21_groupi_n_2015 ,csa_tree_add_24_21_groupi_n_1755);
  or csa_tree_add_24_21_groupi_g5537__6131(csa_tree_add_24_21_groupi_n_2016 ,csa_tree_add_24_21_groupi_n_1712 ,csa_tree_add_24_21_groupi_n_2015);
  and csa_tree_add_24_21_groupi_g5538__1881(csa_tree_add_24_21_groupi_n_2015 ,csa_tree_add_24_21_groupi_n_1806 ,csa_tree_add_24_21_groupi_n_2013);
  xnor csa_tree_add_24_21_groupi_g5539__5115(csa_tree_add_24_21_groupi_n_2014 ,csa_tree_add_24_21_groupi_n_2012 ,csa_tree_add_24_21_groupi_n_1839);
  or csa_tree_add_24_21_groupi_g5540__7482(csa_tree_add_24_21_groupi_n_2013 ,csa_tree_add_24_21_groupi_n_1807 ,csa_tree_add_24_21_groupi_n_2012);
  and csa_tree_add_24_21_groupi_g5541__4733(csa_tree_add_24_21_groupi_n_2012 ,csa_tree_add_24_21_groupi_n_1861 ,csa_tree_add_24_21_groupi_n_2010);
  xnor csa_tree_add_24_21_groupi_g5542__6161(csa_tree_add_24_21_groupi_n_2011 ,csa_tree_add_24_21_groupi_n_2009 ,csa_tree_add_24_21_groupi_n_1878);
  or csa_tree_add_24_21_groupi_g5543__9315(csa_tree_add_24_21_groupi_n_2010 ,csa_tree_add_24_21_groupi_n_1863 ,csa_tree_add_24_21_groupi_n_2009);
  and csa_tree_add_24_21_groupi_g5544__9945(csa_tree_add_24_21_groupi_n_2009 ,csa_tree_add_24_21_groupi_n_1867 ,csa_tree_add_24_21_groupi_n_2007);
  xnor csa_tree_add_24_21_groupi_g5545__2883(csa_tree_add_24_21_groupi_n_2008 ,csa_tree_add_24_21_groupi_n_2006 ,csa_tree_add_24_21_groupi_n_1877);
  or csa_tree_add_24_21_groupi_g5546__2346(csa_tree_add_24_21_groupi_n_2007 ,csa_tree_add_24_21_groupi_n_1842 ,csa_tree_add_24_21_groupi_n_2006);
  and csa_tree_add_24_21_groupi_g5547__1666(csa_tree_add_24_21_groupi_n_2006 ,csa_tree_add_24_21_groupi_n_2004 ,csa_tree_add_24_21_groupi_n_1896);
  xnor csa_tree_add_24_21_groupi_g5548__7410(csa_tree_add_24_21_groupi_n_2005 ,csa_tree_add_24_21_groupi_n_2003 ,csa_tree_add_24_21_groupi_n_1909);
  or csa_tree_add_24_21_groupi_g5549__6417(csa_tree_add_24_21_groupi_n_2004 ,csa_tree_add_24_21_groupi_n_1881 ,csa_tree_add_24_21_groupi_n_2003);
  and csa_tree_add_24_21_groupi_g5550__5477(csa_tree_add_24_21_groupi_n_2003 ,csa_tree_add_24_21_groupi_n_1925 ,csa_tree_add_24_21_groupi_n_2001);
  xnor csa_tree_add_24_21_groupi_g5551__2398(csa_tree_add_24_21_groupi_n_2002 ,csa_tree_add_24_21_groupi_n_2000 ,csa_tree_add_24_21_groupi_n_1936);
  or csa_tree_add_24_21_groupi_g5552__5107(csa_tree_add_24_21_groupi_n_2001 ,csa_tree_add_24_21_groupi_n_1924 ,csa_tree_add_24_21_groupi_n_2000);
  and csa_tree_add_24_21_groupi_g5553__6260(csa_tree_add_24_21_groupi_n_2000 ,csa_tree_add_24_21_groupi_n_1998 ,csa_tree_add_24_21_groupi_n_1911);
  xnor csa_tree_add_24_21_groupi_g5554__4319(csa_tree_add_24_21_groupi_n_1999 ,csa_tree_add_24_21_groupi_n_1997 ,csa_tree_add_24_21_groupi_n_1935);
  or csa_tree_add_24_21_groupi_g5555__8428(csa_tree_add_24_21_groupi_n_1998 ,csa_tree_add_24_21_groupi_n_1913 ,csa_tree_add_24_21_groupi_n_1997);
  and csa_tree_add_24_21_groupi_g5556__5526(csa_tree_add_24_21_groupi_n_1997 ,csa_tree_add_24_21_groupi_n_1995 ,csa_tree_add_24_21_groupi_n_1926);
  xnor csa_tree_add_24_21_groupi_g5557__6783(csa_tree_add_24_21_groupi_n_1996 ,csa_tree_add_24_21_groupi_n_1994 ,csa_tree_add_24_21_groupi_n_1934);
  or csa_tree_add_24_21_groupi_g5558__3680(csa_tree_add_24_21_groupi_n_1995 ,csa_tree_add_24_21_groupi_n_1922 ,csa_tree_add_24_21_groupi_n_1994);
  and csa_tree_add_24_21_groupi_g5559__1617(csa_tree_add_24_21_groupi_n_1994 ,csa_tree_add_24_21_groupi_n_1992 ,csa_tree_add_24_21_groupi_n_1944);
  xnor csa_tree_add_24_21_groupi_g5560__2802(csa_tree_add_24_21_groupi_n_1993 ,csa_tree_add_24_21_groupi_n_1991 ,csa_tree_add_24_21_groupi_n_1954);
  or csa_tree_add_24_21_groupi_g5561__1705(csa_tree_add_24_21_groupi_n_1992 ,csa_tree_add_24_21_groupi_n_1947 ,csa_tree_add_24_21_groupi_n_1991);
  and csa_tree_add_24_21_groupi_g5562__5122(csa_tree_add_24_21_groupi_n_1991 ,csa_tree_add_24_21_groupi_n_1989 ,csa_tree_add_24_21_groupi_n_1927);
  xnor csa_tree_add_24_21_groupi_g5563__8246(csa_tree_add_24_21_groupi_n_1990 ,csa_tree_add_24_21_groupi_n_1988 ,csa_tree_add_24_21_groupi_n_1937);
  or csa_tree_add_24_21_groupi_g5564__7098(csa_tree_add_24_21_groupi_n_1989 ,csa_tree_add_24_21_groupi_n_1929 ,csa_tree_add_24_21_groupi_n_1988);
  and csa_tree_add_24_21_groupi_g5565__6131(csa_tree_add_24_21_groupi_n_1988 ,csa_tree_add_24_21_groupi_n_1986 ,csa_tree_add_24_21_groupi_n_1942);
  xnor csa_tree_add_24_21_groupi_g5566__1881(csa_tree_add_24_21_groupi_n_1987 ,csa_tree_add_24_21_groupi_n_1985 ,csa_tree_add_24_21_groupi_n_1953);
  or csa_tree_add_24_21_groupi_g5567__5115(csa_tree_add_24_21_groupi_n_1986 ,csa_tree_add_24_21_groupi_n_1985 ,csa_tree_add_24_21_groupi_n_1943);
  and csa_tree_add_24_21_groupi_g5568__7482(csa_tree_add_24_21_groupi_n_1985 ,csa_tree_add_24_21_groupi_n_1983 ,csa_tree_add_24_21_groupi_n_1948);
  xnor csa_tree_add_24_21_groupi_g5569__4733(csa_tree_add_24_21_groupi_n_1984 ,csa_tree_add_24_21_groupi_n_1982 ,csa_tree_add_24_21_groupi_n_1952);
  or csa_tree_add_24_21_groupi_g5570__6161(csa_tree_add_24_21_groupi_n_1983 ,csa_tree_add_24_21_groupi_n_1982 ,csa_tree_add_24_21_groupi_n_1945);
  and csa_tree_add_24_21_groupi_g5571__9315(csa_tree_add_24_21_groupi_n_1982 ,csa_tree_add_24_21_groupi_n_1980 ,csa_tree_add_24_21_groupi_n_1938);
  xnor csa_tree_add_24_21_groupi_g5572__9945(csa_tree_add_24_21_groupi_n_1981 ,csa_tree_add_24_21_groupi_n_1979 ,csa_tree_add_24_21_groupi_n_1951);
  or csa_tree_add_24_21_groupi_g5573__2883(csa_tree_add_24_21_groupi_n_1980 ,csa_tree_add_24_21_groupi_n_1940 ,csa_tree_add_24_21_groupi_n_1979);
  and csa_tree_add_24_21_groupi_g5574__2346(csa_tree_add_24_21_groupi_n_1979 ,csa_tree_add_24_21_groupi_n_1977 ,csa_tree_add_24_21_groupi_n_1941);
  xnor csa_tree_add_24_21_groupi_g5575__1666(csa_tree_add_24_21_groupi_n_1978 ,csa_tree_add_24_21_groupi_n_1976 ,csa_tree_add_24_21_groupi_n_1950);
  or csa_tree_add_24_21_groupi_g5576__7410(csa_tree_add_24_21_groupi_n_1977 ,csa_tree_add_24_21_groupi_n_1939 ,csa_tree_add_24_21_groupi_n_1976);
  and csa_tree_add_24_21_groupi_g5577__6417(csa_tree_add_24_21_groupi_n_1976 ,csa_tree_add_24_21_groupi_n_1974 ,csa_tree_add_24_21_groupi_n_1928);
  xnor csa_tree_add_24_21_groupi_g5578__5477(csa_tree_add_24_21_groupi_n_1975 ,csa_tree_add_24_21_groupi_n_1973 ,csa_tree_add_24_21_groupi_n_1933);
  or csa_tree_add_24_21_groupi_g5579__2398(csa_tree_add_24_21_groupi_n_1974 ,csa_tree_add_24_21_groupi_n_1923 ,csa_tree_add_24_21_groupi_n_1973);
  and csa_tree_add_24_21_groupi_g5580__5107(csa_tree_add_24_21_groupi_n_1973 ,csa_tree_add_24_21_groupi_n_1880 ,csa_tree_add_24_21_groupi_n_1971);
  xnor csa_tree_add_24_21_groupi_g5581__6260(csa_tree_add_24_21_groupi_n_1972 ,csa_tree_add_24_21_groupi_n_1970 ,csa_tree_add_24_21_groupi_n_1908);
  or csa_tree_add_24_21_groupi_g5582__4319(csa_tree_add_24_21_groupi_n_1971 ,csa_tree_add_24_21_groupi_n_1882 ,csa_tree_add_24_21_groupi_n_1970);
  and csa_tree_add_24_21_groupi_g5583__8428(csa_tree_add_24_21_groupi_n_1970 ,csa_tree_add_24_21_groupi_n_1968 ,csa_tree_add_24_21_groupi_n_1897);
  xnor csa_tree_add_24_21_groupi_g5584__5526(csa_tree_add_24_21_groupi_n_1969 ,csa_tree_add_24_21_groupi_n_1967 ,csa_tree_add_24_21_groupi_n_1907);
  or csa_tree_add_24_21_groupi_g5585__6783(csa_tree_add_24_21_groupi_n_1968 ,csa_tree_add_24_21_groupi_n_1898 ,csa_tree_add_24_21_groupi_n_1967);
  and csa_tree_add_24_21_groupi_g5586__3680(csa_tree_add_24_21_groupi_n_1967 ,csa_tree_add_24_21_groupi_n_1857 ,csa_tree_add_24_21_groupi_n_1965);
  xnor csa_tree_add_24_21_groupi_g5587__1617(csa_tree_add_24_21_groupi_n_1966 ,csa_tree_add_24_21_groupi_n_1964 ,csa_tree_add_24_21_groupi_n_1879);
  or csa_tree_add_24_21_groupi_g5588__2802(csa_tree_add_24_21_groupi_n_1965 ,csa_tree_add_24_21_groupi_n_1860 ,csa_tree_add_24_21_groupi_n_1964);
  and csa_tree_add_24_21_groupi_g5589__1705(csa_tree_add_24_21_groupi_n_1964 ,csa_tree_add_24_21_groupi_n_1894 ,csa_tree_add_24_21_groupi_n_1962);
  xnor csa_tree_add_24_21_groupi_g5590__5122(csa_tree_add_24_21_groupi_n_1963 ,csa_tree_add_24_21_groupi_n_1961 ,csa_tree_add_24_21_groupi_n_1910);
  or csa_tree_add_24_21_groupi_g5591__8246(csa_tree_add_24_21_groupi_n_1962 ,csa_tree_add_24_21_groupi_n_1895 ,csa_tree_add_24_21_groupi_n_1961);
  and csa_tree_add_24_21_groupi_g5592__7098(csa_tree_add_24_21_groupi_n_1961 ,csa_tree_add_24_21_groupi_n_1801 ,csa_tree_add_24_21_groupi_n_1959);
  xnor csa_tree_add_24_21_groupi_g5593__6131(csa_tree_add_24_21_groupi_n_1960 ,csa_tree_add_24_21_groupi_n_1958 ,csa_tree_add_24_21_groupi_n_1838);
  or csa_tree_add_24_21_groupi_g5594__1881(csa_tree_add_24_21_groupi_n_1959 ,csa_tree_add_24_21_groupi_n_1804 ,csa_tree_add_24_21_groupi_n_1958);
  and csa_tree_add_24_21_groupi_g5595__5115(csa_tree_add_24_21_groupi_n_1958 ,csa_tree_add_24_21_groupi_n_1818 ,csa_tree_add_24_21_groupi_n_1956);
  xnor csa_tree_add_24_21_groupi_g5596__7482(csa_tree_add_24_21_groupi_n_1957 ,csa_tree_add_24_21_groupi_n_1955 ,csa_tree_add_24_21_groupi_n_1837);
  or csa_tree_add_24_21_groupi_g5597__4733(csa_tree_add_24_21_groupi_n_1956 ,csa_tree_add_24_21_groupi_n_1817 ,csa_tree_add_24_21_groupi_n_1955);
  and csa_tree_add_24_21_groupi_g5598__6161(csa_tree_add_24_21_groupi_n_1955 ,csa_tree_add_24_21_groupi_n_1741 ,csa_tree_add_24_21_groupi_n_1946);
  xnor csa_tree_add_24_21_groupi_g5599__9315(csa_tree_add_24_21_groupi_n_1954 ,csa_tree_add_24_21_groupi_n_1931 ,csa_tree_add_24_21_groupi_n_1888);
  xnor csa_tree_add_24_21_groupi_g5600__9945(csa_tree_add_24_21_groupi_n_1953 ,csa_tree_add_24_21_groupi_n_1900 ,csa_tree_add_24_21_groupi_n_1915);
  xnor csa_tree_add_24_21_groupi_g5601__2883(csa_tree_add_24_21_groupi_n_1952 ,csa_tree_add_24_21_groupi_n_1856 ,csa_tree_add_24_21_groupi_n_1921);
  xnor csa_tree_add_24_21_groupi_g5602__2346(csa_tree_add_24_21_groupi_n_1951 ,csa_tree_add_24_21_groupi_n_1906 ,csa_tree_add_24_21_groupi_n_1917);
  xnor csa_tree_add_24_21_groupi_g5603__1666(csa_tree_add_24_21_groupi_n_1950 ,csa_tree_add_24_21_groupi_n_1844 ,csa_tree_add_24_21_groupi_n_1918);
  xnor csa_tree_add_24_21_groupi_g5604__7410(csa_tree_add_24_21_groupi_n_1949 ,csa_tree_add_24_21_groupi_n_1932 ,csa_tree_add_24_21_groupi_n_1754);
  or csa_tree_add_24_21_groupi_g5605__6417(csa_tree_add_24_21_groupi_n_1948 ,csa_tree_add_24_21_groupi_n_1855 ,csa_tree_add_24_21_groupi_n_1921);
  nor csa_tree_add_24_21_groupi_g5606__5477(csa_tree_add_24_21_groupi_n_1947 ,csa_tree_add_24_21_groupi_n_1930 ,csa_tree_add_24_21_groupi_n_1888);
  or csa_tree_add_24_21_groupi_g5607__2398(csa_tree_add_24_21_groupi_n_1946 ,csa_tree_add_24_21_groupi_n_1711 ,csa_tree_add_24_21_groupi_n_1932);
  nor csa_tree_add_24_21_groupi_g5608__5107(csa_tree_add_24_21_groupi_n_1945 ,csa_tree_add_24_21_groupi_n_1856 ,csa_tree_add_24_21_groupi_n_1920);
  or csa_tree_add_24_21_groupi_g5609__6260(csa_tree_add_24_21_groupi_n_1944 ,csa_tree_add_24_21_groupi_n_1931 ,csa_tree_add_24_21_groupi_n_1887);
  nor csa_tree_add_24_21_groupi_g5610__4319(csa_tree_add_24_21_groupi_n_1943 ,csa_tree_add_24_21_groupi_n_1899 ,csa_tree_add_24_21_groupi_n_1915);
  or csa_tree_add_24_21_groupi_g5611__8428(csa_tree_add_24_21_groupi_n_1942 ,csa_tree_add_24_21_groupi_n_1900 ,csa_tree_add_24_21_groupi_n_1914);
  or csa_tree_add_24_21_groupi_g5612__5526(csa_tree_add_24_21_groupi_n_1941 ,csa_tree_add_24_21_groupi_n_1844 ,csa_tree_add_24_21_groupi_n_1919);
  nor csa_tree_add_24_21_groupi_g5613__6783(csa_tree_add_24_21_groupi_n_1940 ,csa_tree_add_24_21_groupi_n_1905 ,csa_tree_add_24_21_groupi_n_1917);
  and csa_tree_add_24_21_groupi_g5614__3680(csa_tree_add_24_21_groupi_n_1939 ,csa_tree_add_24_21_groupi_n_1844 ,csa_tree_add_24_21_groupi_n_1919);
  or csa_tree_add_24_21_groupi_g5615__1617(csa_tree_add_24_21_groupi_n_1938 ,csa_tree_add_24_21_groupi_n_1906 ,csa_tree_add_24_21_groupi_n_1916);
  xnor csa_tree_add_24_21_groupi_g5616__2802(csa_tree_add_24_21_groupi_n_1937 ,csa_tree_add_24_21_groupi_n_1902 ,csa_tree_add_24_21_groupi_n_1884);
  xnor csa_tree_add_24_21_groupi_g5617__1705(csa_tree_add_24_21_groupi_n_1936 ,csa_tree_add_24_21_groupi_n_1869 ,csa_tree_add_24_21_groupi_n_1889);
  xnor csa_tree_add_24_21_groupi_g5618__5122(csa_tree_add_24_21_groupi_n_1935 ,csa_tree_add_24_21_groupi_n_1871 ,csa_tree_add_24_21_groupi_n_1891);
  xnor csa_tree_add_24_21_groupi_g5619__8246(csa_tree_add_24_21_groupi_n_1934 ,csa_tree_add_24_21_groupi_n_1873 ,csa_tree_add_24_21_groupi_n_1886);
  xnor csa_tree_add_24_21_groupi_g5620__7098(csa_tree_add_24_21_groupi_n_1933 ,csa_tree_add_24_21_groupi_n_1904 ,csa_tree_add_24_21_groupi_n_1850);
  not csa_tree_add_24_21_groupi_g5621(csa_tree_add_24_21_groupi_n_1930 ,csa_tree_add_24_21_groupi_n_1931);
  nor csa_tree_add_24_21_groupi_g5622__6131(csa_tree_add_24_21_groupi_n_1929 ,csa_tree_add_24_21_groupi_n_1901 ,csa_tree_add_24_21_groupi_n_1884);
  or csa_tree_add_24_21_groupi_g5623__1881(csa_tree_add_24_21_groupi_n_1928 ,csa_tree_add_24_21_groupi_n_1904 ,csa_tree_add_24_21_groupi_n_1849);
  or csa_tree_add_24_21_groupi_g5624__5115(csa_tree_add_24_21_groupi_n_1927 ,csa_tree_add_24_21_groupi_n_1902 ,csa_tree_add_24_21_groupi_n_1883);
  or csa_tree_add_24_21_groupi_g5625__7482(csa_tree_add_24_21_groupi_n_1926 ,csa_tree_add_24_21_groupi_n_1873 ,csa_tree_add_24_21_groupi_n_1885);
  or csa_tree_add_24_21_groupi_g5626__4733(csa_tree_add_24_21_groupi_n_1925 ,csa_tree_add_24_21_groupi_n_1869 ,csa_tree_add_24_21_groupi_n_0);
  nor csa_tree_add_24_21_groupi_g5627__6161(csa_tree_add_24_21_groupi_n_1924 ,csa_tree_add_24_21_groupi_n_1868 ,csa_tree_add_24_21_groupi_n_1889);
  nor csa_tree_add_24_21_groupi_g5628__9315(csa_tree_add_24_21_groupi_n_1923 ,csa_tree_add_24_21_groupi_n_1903 ,csa_tree_add_24_21_groupi_n_1850);
  nor csa_tree_add_24_21_groupi_g5629__9945(csa_tree_add_24_21_groupi_n_1922 ,csa_tree_add_24_21_groupi_n_1872 ,csa_tree_add_24_21_groupi_n_1886);
  and csa_tree_add_24_21_groupi_g5630__2883(csa_tree_add_24_21_groupi_n_1932 ,csa_tree_add_24_21_groupi_n_1716 ,csa_tree_add_24_21_groupi_n_1893);
  and csa_tree_add_24_21_groupi_g5631__2346(csa_tree_add_24_21_groupi_n_1931 ,csa_tree_add_24_21_groupi_n_1859 ,csa_tree_add_24_21_groupi_n_1892);
  not csa_tree_add_24_21_groupi_g5632(csa_tree_add_24_21_groupi_n_1920 ,csa_tree_add_24_21_groupi_n_1921);
  not csa_tree_add_24_21_groupi_g5633(csa_tree_add_24_21_groupi_n_1919 ,csa_tree_add_24_21_groupi_n_1918);
  not csa_tree_add_24_21_groupi_g5634(csa_tree_add_24_21_groupi_n_1917 ,csa_tree_add_24_21_groupi_n_1916);
  not csa_tree_add_24_21_groupi_g5635(csa_tree_add_24_21_groupi_n_1914 ,csa_tree_add_24_21_groupi_n_1915);
  nor csa_tree_add_24_21_groupi_g5636__1666(csa_tree_add_24_21_groupi_n_1913 ,csa_tree_add_24_21_groupi_n_1870 ,csa_tree_add_24_21_groupi_n_1891);
  xnor csa_tree_add_24_21_groupi_g5637__7410(csa_tree_add_24_21_groupi_n_1912 ,csa_tree_add_24_21_groupi_n_1876 ,csa_tree_add_24_21_groupi_n_1756);
  or csa_tree_add_24_21_groupi_g5638__6417(csa_tree_add_24_21_groupi_n_1911 ,csa_tree_add_24_21_groupi_n_1871 ,csa_tree_add_24_21_groupi_n_1890);
  xnor csa_tree_add_24_21_groupi_g5639__5477(csa_tree_add_24_21_groupi_n_1910 ,csa_tree_add_24_21_groupi_n_1743 ,csa_tree_add_24_21_groupi_n_1852);
  xnor csa_tree_add_24_21_groupi_g5640__2398(csa_tree_add_24_21_groupi_n_1909 ,csa_tree_add_24_21_groupi_n_1843 ,csa_tree_add_24_21_groupi_n_1853);
  xnor csa_tree_add_24_21_groupi_g5641__5107(csa_tree_add_24_21_groupi_n_1908 ,csa_tree_add_24_21_groupi_n_1811 ,csa_tree_add_24_21_groupi_n_1848);
  xnor csa_tree_add_24_21_groupi_g5642__6260(csa_tree_add_24_21_groupi_n_1907 ,csa_tree_add_24_21_groupi_n_1875 ,csa_tree_add_24_21_groupi_n_1846);
  xnor csa_tree_add_24_21_groupi_g5643__4319(csa_tree_add_24_21_groupi_n_1921 ,csa_tree_add_24_21_groupi_n_1746 ,csa_tree_add_24_21_groupi_n_1840);
  xnor csa_tree_add_24_21_groupi_g5644__8428(csa_tree_add_24_21_groupi_n_1918 ,csa_tree_add_24_21_groupi_n_1748 ,csa_tree_add_24_21_groupi_n_1836);
  xnor csa_tree_add_24_21_groupi_g5645__5526(csa_tree_add_24_21_groupi_n_1916 ,csa_tree_add_24_21_groupi_n_1745 ,csa_tree_add_24_21_groupi_n_1);
  xnor csa_tree_add_24_21_groupi_g5646__6783(csa_tree_add_24_21_groupi_n_1915 ,csa_tree_add_24_21_groupi_n_1751 ,csa_tree_add_24_21_groupi_n_1835);
  not csa_tree_add_24_21_groupi_g5647(csa_tree_add_24_21_groupi_n_1906 ,csa_tree_add_24_21_groupi_n_1905);
  not csa_tree_add_24_21_groupi_g5648(csa_tree_add_24_21_groupi_n_1903 ,csa_tree_add_24_21_groupi_n_1904);
  not csa_tree_add_24_21_groupi_g5649(csa_tree_add_24_21_groupi_n_1901 ,csa_tree_add_24_21_groupi_n_1902);
  not csa_tree_add_24_21_groupi_g5650(csa_tree_add_24_21_groupi_n_1900 ,csa_tree_add_24_21_groupi_n_1899);
  nor csa_tree_add_24_21_groupi_g5651__3680(csa_tree_add_24_21_groupi_n_1898 ,csa_tree_add_24_21_groupi_n_1874 ,csa_tree_add_24_21_groupi_n_1846);
  or csa_tree_add_24_21_groupi_g5652__1617(csa_tree_add_24_21_groupi_n_1897 ,csa_tree_add_24_21_groupi_n_1875 ,csa_tree_add_24_21_groupi_n_1845);
  or csa_tree_add_24_21_groupi_g5653__2802(csa_tree_add_24_21_groupi_n_1896 ,csa_tree_add_24_21_groupi_n_1843 ,csa_tree_add_24_21_groupi_n_1854);
  nor csa_tree_add_24_21_groupi_g5654__1705(csa_tree_add_24_21_groupi_n_1895 ,csa_tree_add_24_21_groupi_n_1742 ,csa_tree_add_24_21_groupi_n_1852);
  or csa_tree_add_24_21_groupi_g5655__5122(csa_tree_add_24_21_groupi_n_1894 ,csa_tree_add_24_21_groupi_n_1743 ,csa_tree_add_24_21_groupi_n_1851);
  or csa_tree_add_24_21_groupi_g5656__8246(csa_tree_add_24_21_groupi_n_1893 ,csa_tree_add_24_21_groupi_n_1713 ,csa_tree_add_24_21_groupi_n_1876);
  or csa_tree_add_24_21_groupi_g5657__7098(csa_tree_add_24_21_groupi_n_1892 ,csa_tree_add_24_21_groupi_n_1750 ,csa_tree_add_24_21_groupi_n_1858);
  or csa_tree_add_24_21_groupi_g5658__6131(csa_tree_add_24_21_groupi_n_1905 ,csa_tree_add_24_21_groupi_n_1827 ,csa_tree_add_24_21_groupi_n_1864);
  and csa_tree_add_24_21_groupi_g5659__1881(csa_tree_add_24_21_groupi_n_1904 ,csa_tree_add_24_21_groupi_n_1820 ,csa_tree_add_24_21_groupi_n_1862);
  and csa_tree_add_24_21_groupi_g5660__5115(csa_tree_add_24_21_groupi_n_1902 ,csa_tree_add_24_21_groupi_n_1831 ,csa_tree_add_24_21_groupi_n_1865);
  or csa_tree_add_24_21_groupi_g5661__7482(csa_tree_add_24_21_groupi_n_1899 ,csa_tree_add_24_21_groupi_n_1830 ,csa_tree_add_24_21_groupi_n_1866);
  not csa_tree_add_24_21_groupi_g5662(csa_tree_add_24_21_groupi_n_1891 ,csa_tree_add_24_21_groupi_n_1890);
  not csa_tree_add_24_21_groupi_g5663(csa_tree_add_24_21_groupi_n_1889 ,csa_tree_add_24_21_groupi_n_0);
  not csa_tree_add_24_21_groupi_g5664(csa_tree_add_24_21_groupi_n_1887 ,csa_tree_add_24_21_groupi_n_1888);
  not csa_tree_add_24_21_groupi_g5665(csa_tree_add_24_21_groupi_n_1886 ,csa_tree_add_24_21_groupi_n_1885);
  not csa_tree_add_24_21_groupi_g5666(csa_tree_add_24_21_groupi_n_1883 ,csa_tree_add_24_21_groupi_n_1884);
  nor csa_tree_add_24_21_groupi_g5667__4733(csa_tree_add_24_21_groupi_n_1882 ,csa_tree_add_24_21_groupi_n_1810 ,csa_tree_add_24_21_groupi_n_1848);
  and csa_tree_add_24_21_groupi_g5668__6161(csa_tree_add_24_21_groupi_n_1881 ,csa_tree_add_24_21_groupi_n_1843 ,csa_tree_add_24_21_groupi_n_1854);
  or csa_tree_add_24_21_groupi_g5669__9315(csa_tree_add_24_21_groupi_n_1880 ,csa_tree_add_24_21_groupi_n_1811 ,csa_tree_add_24_21_groupi_n_1847);
  xnor csa_tree_add_24_21_groupi_g5670__9945(csa_tree_add_24_21_groupi_n_1879 ,csa_tree_add_24_21_groupi_n_1834 ,csa_tree_add_24_21_groupi_n_1813);
  xnor csa_tree_add_24_21_groupi_g5671__2883(csa_tree_add_24_21_groupi_n_1878 ,csa_tree_add_24_21_groupi_n_1794 ,csa_tree_add_24_21_groupi_n_1815);
  xnor csa_tree_add_24_21_groupi_g5672__2346(csa_tree_add_24_21_groupi_n_1877 ,csa_tree_add_24_21_groupi_n_1832 ,csa_tree_add_24_21_groupi_n_1808);
  xnor csa_tree_add_24_21_groupi_g5673__1666(csa_tree_add_24_21_groupi_n_1890 ,csa_tree_add_24_21_groupi_n_1747 ,csa_tree_add_24_21_groupi_n_1796);
  xnor csa_tree_add_24_21_groupi_g5675__7410(csa_tree_add_24_21_groupi_n_1888 ,csa_tree_add_24_21_groupi_n_1725 ,csa_tree_add_24_21_groupi_n_1799);
  xnor csa_tree_add_24_21_groupi_g5676__6417(csa_tree_add_24_21_groupi_n_1885 ,csa_tree_add_24_21_groupi_n_1752 ,csa_tree_add_24_21_groupi_n_1798);
  xnor csa_tree_add_24_21_groupi_g5677__5477(csa_tree_add_24_21_groupi_n_1884 ,csa_tree_add_24_21_groupi_n_1816 ,csa_tree_add_24_21_groupi_n_1800);
  not csa_tree_add_24_21_groupi_g5678(csa_tree_add_24_21_groupi_n_1874 ,csa_tree_add_24_21_groupi_n_1875);
  not csa_tree_add_24_21_groupi_g5679(csa_tree_add_24_21_groupi_n_1872 ,csa_tree_add_24_21_groupi_n_1873);
  not csa_tree_add_24_21_groupi_g5680(csa_tree_add_24_21_groupi_n_1870 ,csa_tree_add_24_21_groupi_n_1871);
  not csa_tree_add_24_21_groupi_g5681(csa_tree_add_24_21_groupi_n_1868 ,csa_tree_add_24_21_groupi_n_1869);
  or csa_tree_add_24_21_groupi_g5682__2398(csa_tree_add_24_21_groupi_n_1867 ,csa_tree_add_24_21_groupi_n_1832 ,csa_tree_add_24_21_groupi_n_1809);
  nor csa_tree_add_24_21_groupi_g5683__5107(csa_tree_add_24_21_groupi_n_1866 ,csa_tree_add_24_21_groupi_n_1746 ,csa_tree_add_24_21_groupi_n_1829);
  or csa_tree_add_24_21_groupi_g5684__6260(csa_tree_add_24_21_groupi_n_1865 ,csa_tree_add_24_21_groupi_n_1751 ,csa_tree_add_24_21_groupi_n_1828);
  nor csa_tree_add_24_21_groupi_g5685__4319(csa_tree_add_24_21_groupi_n_1864 ,csa_tree_add_24_21_groupi_n_1748 ,csa_tree_add_24_21_groupi_n_1825);
  nor csa_tree_add_24_21_groupi_g5686__8428(csa_tree_add_24_21_groupi_n_1863 ,csa_tree_add_24_21_groupi_n_1793 ,csa_tree_add_24_21_groupi_n_1815);
  or csa_tree_add_24_21_groupi_g5687__5526(csa_tree_add_24_21_groupi_n_1862 ,csa_tree_add_24_21_groupi_n_1637 ,csa_tree_add_24_21_groupi_n_1819);
  or csa_tree_add_24_21_groupi_g5688__6783(csa_tree_add_24_21_groupi_n_1861 ,csa_tree_add_24_21_groupi_n_1794 ,csa_tree_add_24_21_groupi_n_1814);
  nor csa_tree_add_24_21_groupi_g5689__3680(csa_tree_add_24_21_groupi_n_1860 ,csa_tree_add_24_21_groupi_n_1833 ,csa_tree_add_24_21_groupi_n_1813);
  or csa_tree_add_24_21_groupi_g5690__1617(csa_tree_add_24_21_groupi_n_1859 ,csa_tree_add_24_21_groupi_n_1662 ,csa_tree_add_24_21_groupi_n_1816);
  and csa_tree_add_24_21_groupi_g5691__2802(csa_tree_add_24_21_groupi_n_1858 ,csa_tree_add_24_21_groupi_n_1662 ,csa_tree_add_24_21_groupi_n_1816);
  or csa_tree_add_24_21_groupi_g5692__1705(csa_tree_add_24_21_groupi_n_1857 ,csa_tree_add_24_21_groupi_n_1834 ,csa_tree_add_24_21_groupi_n_1812);
  and csa_tree_add_24_21_groupi_g5693__5122(csa_tree_add_24_21_groupi_n_1876 ,csa_tree_add_24_21_groupi_n_1652 ,csa_tree_add_24_21_groupi_n_1823);
  and csa_tree_add_24_21_groupi_g5694__8246(csa_tree_add_24_21_groupi_n_1875 ,csa_tree_add_24_21_groupi_n_1761 ,csa_tree_add_24_21_groupi_n_1821);
  and csa_tree_add_24_21_groupi_g5695__7098(csa_tree_add_24_21_groupi_n_1873 ,csa_tree_add_24_21_groupi_n_1786 ,csa_tree_add_24_21_groupi_n_1822);
  and csa_tree_add_24_21_groupi_g5696__6131(csa_tree_add_24_21_groupi_n_1871 ,csa_tree_add_24_21_groupi_n_1782 ,csa_tree_add_24_21_groupi_n_1824);
  and csa_tree_add_24_21_groupi_g5697__1881(csa_tree_add_24_21_groupi_n_1869 ,csa_tree_add_24_21_groupi_n_1780 ,csa_tree_add_24_21_groupi_n_1826);
  not csa_tree_add_24_21_groupi_g5698(csa_tree_add_24_21_groupi_n_1856 ,csa_tree_add_24_21_groupi_n_1855);
  not csa_tree_add_24_21_groupi_g5699(csa_tree_add_24_21_groupi_n_1854 ,csa_tree_add_24_21_groupi_n_1853);
  not csa_tree_add_24_21_groupi_g5700(csa_tree_add_24_21_groupi_n_1851 ,csa_tree_add_24_21_groupi_n_1852);
  not csa_tree_add_24_21_groupi_g5701(csa_tree_add_24_21_groupi_n_1850 ,csa_tree_add_24_21_groupi_n_1849);
  not csa_tree_add_24_21_groupi_g5702(csa_tree_add_24_21_groupi_n_1848 ,csa_tree_add_24_21_groupi_n_1847);
  not csa_tree_add_24_21_groupi_g5703(csa_tree_add_24_21_groupi_n_1846 ,csa_tree_add_24_21_groupi_n_1845);
  and csa_tree_add_24_21_groupi_g5704__5115(csa_tree_add_24_21_groupi_n_1842 ,csa_tree_add_24_21_groupi_n_1832 ,csa_tree_add_24_21_groupi_n_1809);
  xnor csa_tree_add_24_21_groupi_g5705__7482(csa_tree_add_24_21_groupi_n_1841 ,csa_tree_add_24_21_groupi_n_1795 ,csa_tree_add_24_21_groupi_n_1705);
  xnor csa_tree_add_24_21_groupi_g5706__4733(csa_tree_add_24_21_groupi_n_1840 ,csa_tree_add_24_21_groupi_n_1673 ,csa_tree_add_24_21_groupi_n_1764);
  xnor csa_tree_add_24_21_groupi_g5707__6161(csa_tree_add_24_21_groupi_n_1839 ,csa_tree_add_24_21_groupi_n_1729 ,csa_tree_add_24_21_groupi_n_1792);
  xnor csa_tree_add_24_21_groupi_g5708__9315(csa_tree_add_24_21_groupi_n_1838 ,csa_tree_add_24_21_groupi_n_1790 ,csa_tree_add_24_21_groupi_n_1770);
  xnor csa_tree_add_24_21_groupi_g5709__9945(csa_tree_add_24_21_groupi_n_1837 ,csa_tree_add_24_21_groupi_n_1603 ,csa_tree_add_24_21_groupi_n_1772);
  xnor csa_tree_add_24_21_groupi_g5711__2883(csa_tree_add_24_21_groupi_n_1836 ,csa_tree_add_24_21_groupi_n_1671 ,csa_tree_add_24_21_groupi_n_1768);
  xnor csa_tree_add_24_21_groupi_g5712__2346(csa_tree_add_24_21_groupi_n_1835 ,csa_tree_add_24_21_groupi_n_1655 ,csa_tree_add_24_21_groupi_n_1767);
  and csa_tree_add_24_21_groupi_g5713__1666(csa_tree_add_24_21_groupi_n_1855 ,csa_tree_add_24_21_groupi_n_1788 ,csa_tree_add_24_21_groupi_n_1802);
  xnor csa_tree_add_24_21_groupi_g5714__7410(csa_tree_add_24_21_groupi_n_1853 ,csa_tree_add_24_21_groupi_n_1730 ,csa_tree_add_24_21_groupi_n_1757);
  xnor csa_tree_add_24_21_groupi_g5715__6417(csa_tree_add_24_21_groupi_n_1852 ,csa_tree_add_24_21_groupi_n_1584 ,csa_tree_add_24_21_groupi_n_1759);
  xnor csa_tree_add_24_21_groupi_g5716__5477(csa_tree_add_24_21_groupi_n_1849 ,csa_tree_add_24_21_groupi_n_1773 ,csa_tree_add_24_21_groupi_n_1760);
  xnor csa_tree_add_24_21_groupi_g5717__2398(csa_tree_add_24_21_groupi_n_1847 ,csa_tree_add_24_21_groupi_n_1765 ,csa_tree_add_24_21_groupi_n_1707);
  xnor csa_tree_add_24_21_groupi_g5718__5107(csa_tree_add_24_21_groupi_n_1845 ,csa_tree_add_24_21_groupi_n_1701 ,csa_tree_add_24_21_groupi_n_1758);
  and csa_tree_add_24_21_groupi_g5719__6260(csa_tree_add_24_21_groupi_n_1844 ,csa_tree_add_24_21_groupi_n_1735 ,csa_tree_add_24_21_groupi_n_1803);
  and csa_tree_add_24_21_groupi_g5720__4319(csa_tree_add_24_21_groupi_n_1843 ,csa_tree_add_24_21_groupi_n_1777 ,csa_tree_add_24_21_groupi_n_1805);
  not csa_tree_add_24_21_groupi_g5721(csa_tree_add_24_21_groupi_n_1833 ,csa_tree_add_24_21_groupi_n_1834);
  or csa_tree_add_24_21_groupi_g5722__8428(csa_tree_add_24_21_groupi_n_1831 ,csa_tree_add_24_21_groupi_n_1654 ,csa_tree_add_24_21_groupi_n_1767);
  and csa_tree_add_24_21_groupi_g5723__5526(csa_tree_add_24_21_groupi_n_1830 ,csa_tree_add_24_21_groupi_n_1673 ,csa_tree_add_24_21_groupi_n_1764);
  nor csa_tree_add_24_21_groupi_g5724__6783(csa_tree_add_24_21_groupi_n_1829 ,csa_tree_add_24_21_groupi_n_1673 ,csa_tree_add_24_21_groupi_n_1764);
  nor csa_tree_add_24_21_groupi_g5725__3680(csa_tree_add_24_21_groupi_n_1828 ,csa_tree_add_24_21_groupi_n_1655 ,csa_tree_add_24_21_groupi_n_1766);
  nor csa_tree_add_24_21_groupi_g5726__1617(csa_tree_add_24_21_groupi_n_1827 ,csa_tree_add_24_21_groupi_n_1672 ,csa_tree_add_24_21_groupi_n_1768);
  or csa_tree_add_24_21_groupi_g5727__2802(csa_tree_add_24_21_groupi_n_1826 ,csa_tree_add_24_21_groupi_n_1747 ,csa_tree_add_24_21_groupi_n_1783);
  and csa_tree_add_24_21_groupi_g5728__1705(csa_tree_add_24_21_groupi_n_1825 ,csa_tree_add_24_21_groupi_n_1672 ,csa_tree_add_24_21_groupi_n_1768);
  or csa_tree_add_24_21_groupi_g5729__5122(csa_tree_add_24_21_groupi_n_1824 ,csa_tree_add_24_21_groupi_n_1752 ,csa_tree_add_24_21_groupi_n_1781);
  or csa_tree_add_24_21_groupi_g5730__8246(csa_tree_add_24_21_groupi_n_1823 ,csa_tree_add_24_21_groupi_n_1653 ,csa_tree_add_24_21_groupi_n_1795);
  or csa_tree_add_24_21_groupi_g5731__7098(csa_tree_add_24_21_groupi_n_1822 ,csa_tree_add_24_21_groupi_n_1753 ,csa_tree_add_24_21_groupi_n_1784);
  or csa_tree_add_24_21_groupi_g5732__6131(csa_tree_add_24_21_groupi_n_1821 ,csa_tree_add_24_21_groupi_n_1640 ,csa_tree_add_24_21_groupi_n_1763);
  or csa_tree_add_24_21_groupi_g5733__1881(csa_tree_add_24_21_groupi_n_1820 ,csa_tree_add_24_21_groupi_n_1608 ,csa_tree_add_24_21_groupi_n_1765);
  and csa_tree_add_24_21_groupi_g5734__5115(csa_tree_add_24_21_groupi_n_1819 ,csa_tree_add_24_21_groupi_n_1608 ,csa_tree_add_24_21_groupi_n_1765);
  or csa_tree_add_24_21_groupi_g5735__7482(csa_tree_add_24_21_groupi_n_1818 ,csa_tree_add_24_21_groupi_n_1603 ,csa_tree_add_24_21_groupi_n_1771);
  nor csa_tree_add_24_21_groupi_g5736__4733(csa_tree_add_24_21_groupi_n_1817 ,csa_tree_add_24_21_groupi_n_1602 ,csa_tree_add_24_21_groupi_n_1772);
  and csa_tree_add_24_21_groupi_g5737__6161(csa_tree_add_24_21_groupi_n_1834 ,csa_tree_add_24_21_groupi_n_1739 ,csa_tree_add_24_21_groupi_n_1779);
  and csa_tree_add_24_21_groupi_g5738__9315(csa_tree_add_24_21_groupi_n_1832 ,csa_tree_add_24_21_groupi_n_1731 ,csa_tree_add_24_21_groupi_n_1785);
  not csa_tree_add_24_21_groupi_g5739(csa_tree_add_24_21_groupi_n_1815 ,csa_tree_add_24_21_groupi_n_1814);
  not csa_tree_add_24_21_groupi_g5740(csa_tree_add_24_21_groupi_n_1813 ,csa_tree_add_24_21_groupi_n_1812);
  not csa_tree_add_24_21_groupi_g5741(csa_tree_add_24_21_groupi_n_1811 ,csa_tree_add_24_21_groupi_n_1810);
  not csa_tree_add_24_21_groupi_g5742(csa_tree_add_24_21_groupi_n_1809 ,csa_tree_add_24_21_groupi_n_1808);
  nor csa_tree_add_24_21_groupi_g5743__9945(csa_tree_add_24_21_groupi_n_1807 ,csa_tree_add_24_21_groupi_n_1729 ,csa_tree_add_24_21_groupi_n_1791);
  or csa_tree_add_24_21_groupi_g5744__2883(csa_tree_add_24_21_groupi_n_1806 ,csa_tree_add_24_21_groupi_n_1728 ,csa_tree_add_24_21_groupi_n_1792);
  or csa_tree_add_24_21_groupi_g5745__2346(csa_tree_add_24_21_groupi_n_1805 ,csa_tree_add_24_21_groupi_n_1749 ,csa_tree_add_24_21_groupi_n_1776);
  nor csa_tree_add_24_21_groupi_g5746__1666(csa_tree_add_24_21_groupi_n_1804 ,csa_tree_add_24_21_groupi_n_1789 ,csa_tree_add_24_21_groupi_n_1770);
  or csa_tree_add_24_21_groupi_g5747__7410(csa_tree_add_24_21_groupi_n_1803 ,csa_tree_add_24_21_groupi_n_1774 ,csa_tree_add_24_21_groupi_n_1733);
  or csa_tree_add_24_21_groupi_g5748__6417(csa_tree_add_24_21_groupi_n_1802 ,csa_tree_add_24_21_groupi_n_1787 ,csa_tree_add_24_21_groupi_n_1775);
  or csa_tree_add_24_21_groupi_g5749__5477(csa_tree_add_24_21_groupi_n_1801 ,csa_tree_add_24_21_groupi_n_1790 ,csa_tree_add_24_21_groupi_n_1769);
  xor csa_tree_add_24_21_groupi_g5750__2398(csa_tree_add_24_21_groupi_n_1800 ,csa_tree_add_24_21_groupi_n_1750 ,csa_tree_add_24_21_groupi_n_1662);
  xnor csa_tree_add_24_21_groupi_g5751__5107(csa_tree_add_24_21_groupi_n_1799 ,csa_tree_add_24_21_groupi_n_1675 ,csa_tree_add_24_21_groupi_n_1753);
  xnor csa_tree_add_24_21_groupi_g5752__6260(csa_tree_add_24_21_groupi_n_1798 ,csa_tree_add_24_21_groupi_n_1610 ,csa_tree_add_24_21_groupi_n_1723);
  xnor csa_tree_add_24_21_groupi_g5753__4319(csa_tree_add_24_21_groupi_n_1797 ,csa_tree_add_24_21_groupi_n_1580 ,csa_tree_add_24_21_groupi_n_1727);
  xnor csa_tree_add_24_21_groupi_g5754__8428(csa_tree_add_24_21_groupi_n_1796 ,csa_tree_add_24_21_groupi_n_1612 ,csa_tree_add_24_21_groupi_n_1721);
  xnor csa_tree_add_24_21_groupi_g5755__5526(csa_tree_add_24_21_groupi_n_1816 ,csa_tree_add_24_21_groupi_n_1543 ,csa_tree_add_24_21_groupi_n_1706);
  xnor csa_tree_add_24_21_groupi_g5756__6783(csa_tree_add_24_21_groupi_n_1814 ,csa_tree_add_24_21_groupi_n_1615 ,csa_tree_add_24_21_groupi_n_1703);
  xnor csa_tree_add_24_21_groupi_g5757__3680(csa_tree_add_24_21_groupi_n_1812 ,csa_tree_add_24_21_groupi_n_1719 ,csa_tree_add_24_21_groupi_n_1709);
  or csa_tree_add_24_21_groupi_g5758__1617(csa_tree_add_24_21_groupi_n_1810 ,csa_tree_add_24_21_groupi_n_1732 ,csa_tree_add_24_21_groupi_n_1778);
  xnor csa_tree_add_24_21_groupi_g5759__2802(csa_tree_add_24_21_groupi_n_1808 ,csa_tree_add_24_21_groupi_n_1702 ,csa_tree_add_24_21_groupi_n_1708);
  not csa_tree_add_24_21_groupi_g5760(csa_tree_add_24_21_groupi_n_1793 ,csa_tree_add_24_21_groupi_n_1794);
  not csa_tree_add_24_21_groupi_g5761(csa_tree_add_24_21_groupi_n_1791 ,csa_tree_add_24_21_groupi_n_1792);
  not csa_tree_add_24_21_groupi_g5762(csa_tree_add_24_21_groupi_n_1790 ,csa_tree_add_24_21_groupi_n_1789);
  or csa_tree_add_24_21_groupi_g5763__1705(csa_tree_add_24_21_groupi_n_1788 ,csa_tree_add_24_21_groupi_n_1745 ,csa_tree_add_24_21_groupi_n_1669);
  nor csa_tree_add_24_21_groupi_g5764__5122(csa_tree_add_24_21_groupi_n_1787 ,csa_tree_add_24_21_groupi_n_1744 ,csa_tree_add_24_21_groupi_n_1670);
  or csa_tree_add_24_21_groupi_g5765__8246(csa_tree_add_24_21_groupi_n_1786 ,csa_tree_add_24_21_groupi_n_1674 ,csa_tree_add_24_21_groupi_n_1725);
  or csa_tree_add_24_21_groupi_g5766__7098(csa_tree_add_24_21_groupi_n_1785 ,csa_tree_add_24_21_groupi_n_1730 ,csa_tree_add_24_21_groupi_n_1736);
  nor csa_tree_add_24_21_groupi_g5767__6131(csa_tree_add_24_21_groupi_n_1784 ,csa_tree_add_24_21_groupi_n_1675 ,csa_tree_add_24_21_groupi_n_1724);
  nor csa_tree_add_24_21_groupi_g5768__1881(csa_tree_add_24_21_groupi_n_1783 ,csa_tree_add_24_21_groupi_n_1612 ,csa_tree_add_24_21_groupi_n_1721);
  or csa_tree_add_24_21_groupi_g5769__5115(csa_tree_add_24_21_groupi_n_1782 ,csa_tree_add_24_21_groupi_n_1609 ,csa_tree_add_24_21_groupi_n_1722);
  nor csa_tree_add_24_21_groupi_g5770__7482(csa_tree_add_24_21_groupi_n_1781 ,csa_tree_add_24_21_groupi_n_1610 ,csa_tree_add_24_21_groupi_n_1723);
  or csa_tree_add_24_21_groupi_g5771__4733(csa_tree_add_24_21_groupi_n_1780 ,csa_tree_add_24_21_groupi_n_1611 ,csa_tree_add_24_21_groupi_n_1720);
  or csa_tree_add_24_21_groupi_g5772__6161(csa_tree_add_24_21_groupi_n_1779 ,csa_tree_add_24_21_groupi_n_1584 ,csa_tree_add_24_21_groupi_n_1740);
  and csa_tree_add_24_21_groupi_g5773__9315(csa_tree_add_24_21_groupi_n_1778 ,csa_tree_add_24_21_groupi_n_1701 ,csa_tree_add_24_21_groupi_n_1734);
  or csa_tree_add_24_21_groupi_g5774__9945(csa_tree_add_24_21_groupi_n_1777 ,csa_tree_add_24_21_groupi_n_1580 ,csa_tree_add_24_21_groupi_n_1726);
  nor csa_tree_add_24_21_groupi_g5775__2883(csa_tree_add_24_21_groupi_n_1776 ,csa_tree_add_24_21_groupi_n_1579 ,csa_tree_add_24_21_groupi_n_1727);
  and csa_tree_add_24_21_groupi_g5776__2346(csa_tree_add_24_21_groupi_n_1795 ,csa_tree_add_24_21_groupi_n_1448 ,csa_tree_add_24_21_groupi_n_1714);
  and csa_tree_add_24_21_groupi_g5777__1666(csa_tree_add_24_21_groupi_n_1794 ,csa_tree_add_24_21_groupi_n_1692 ,csa_tree_add_24_21_groupi_n_1715);
  and csa_tree_add_24_21_groupi_g5778__7410(csa_tree_add_24_21_groupi_n_1792 ,csa_tree_add_24_21_groupi_n_1688 ,csa_tree_add_24_21_groupi_n_1738);
  or csa_tree_add_24_21_groupi_g5779__6417(csa_tree_add_24_21_groupi_n_1789 ,csa_tree_add_24_21_groupi_n_1454 ,csa_tree_add_24_21_groupi_n_1737);
  not csa_tree_add_24_21_groupi_g5781(csa_tree_add_24_21_groupi_n_1774 ,csa_tree_add_24_21_groupi_n_1773);
  not csa_tree_add_24_21_groupi_g5782(csa_tree_add_24_21_groupi_n_1772 ,csa_tree_add_24_21_groupi_n_1771);
  not csa_tree_add_24_21_groupi_g5783(csa_tree_add_24_21_groupi_n_1770 ,csa_tree_add_24_21_groupi_n_1769);
  not csa_tree_add_24_21_groupi_g5784(csa_tree_add_24_21_groupi_n_1766 ,csa_tree_add_24_21_groupi_n_1767);
  nor csa_tree_add_24_21_groupi_g5785__5477(csa_tree_add_24_21_groupi_n_1763 ,csa_tree_add_24_21_groupi_n_1550 ,csa_tree_add_24_21_groupi_n_1719);
  xnor csa_tree_add_24_21_groupi_g5786__2398(csa_tree_add_24_21_groupi_n_1762 ,csa_tree_add_24_21_groupi_n_1700 ,csa_tree_add_24_21_groupi_n_1531);
  or csa_tree_add_24_21_groupi_g5787__5107(csa_tree_add_24_21_groupi_n_1761 ,csa_tree_add_24_21_groupi_n_1549 ,csa_tree_add_24_21_groupi_n_1718);
  xnor csa_tree_add_24_21_groupi_g5788__6260(csa_tree_add_24_21_groupi_n_1760 ,csa_tree_add_24_21_groupi_n_1664 ,csa_tree_add_24_21_groupi_n_1699);
  xnor csa_tree_add_24_21_groupi_g5789__4319(csa_tree_add_24_21_groupi_n_1759 ,csa_tree_add_24_21_groupi_n_1368 ,csa_tree_add_24_21_groupi_n_1657);
  xnor csa_tree_add_24_21_groupi_g5790__8428(csa_tree_add_24_21_groupi_n_1758 ,csa_tree_add_24_21_groupi_n_1614 ,csa_tree_add_24_21_groupi_n_1659);
  xnor csa_tree_add_24_21_groupi_g5791__5526(csa_tree_add_24_21_groupi_n_1757 ,csa_tree_add_24_21_groupi_n_1463 ,csa_tree_add_24_21_groupi_n_1668);
  xnor csa_tree_add_24_21_groupi_g5792__6783(csa_tree_add_24_21_groupi_n_1756 ,csa_tree_add_24_21_groupi_n_1633 ,csa_tree_add_24_21_groupi_n_1677);
  xnor csa_tree_add_24_21_groupi_g5793__3680(csa_tree_add_24_21_groupi_n_1755 ,csa_tree_add_24_21_groupi_n_1661 ,csa_tree_add_24_21_groupi_n_1697);
  xnor csa_tree_add_24_21_groupi_g5794__1617(csa_tree_add_24_21_groupi_n_1754 ,csa_tree_add_24_21_groupi_n_1599 ,csa_tree_add_24_21_groupi_n_1665);
  xnor csa_tree_add_24_21_groupi_g5795__2802(csa_tree_add_24_21_groupi_n_1775 ,csa_tree_add_24_21_groupi_n_1636 ,csa_tree_add_24_21_groupi_n_1650);
  xnor csa_tree_add_24_21_groupi_g5796__1705(csa_tree_add_24_21_groupi_n_1773 ,csa_tree_add_24_21_groupi_n_1639 ,csa_tree_add_24_21_groupi_n_1649);
  xnor csa_tree_add_24_21_groupi_g5797__5122(csa_tree_add_24_21_groupi_n_1771 ,csa_tree_add_24_21_groupi_n_1678 ,csa_tree_add_24_21_groupi_n_1529);
  xnor csa_tree_add_24_21_groupi_g5798__8246(csa_tree_add_24_21_groupi_n_1769 ,csa_tree_add_24_21_groupi_n_1616 ,csa_tree_add_24_21_groupi_n_1651);
  xnor csa_tree_add_24_21_groupi_g5799__7098(csa_tree_add_24_21_groupi_n_1768 ,csa_tree_add_24_21_groupi_n_1644 ,csa_tree_add_24_21_groupi_n_1647);
  xnor csa_tree_add_24_21_groupi_g5800__6131(csa_tree_add_24_21_groupi_n_1767 ,csa_tree_add_24_21_groupi_n_1635 ,csa_tree_add_24_21_groupi_n_1648);
  xnor csa_tree_add_24_21_groupi_g5801__1881(csa_tree_add_24_21_groupi_n_1765 ,csa_tree_add_24_21_groupi_n_1465 ,csa_tree_add_24_21_groupi_n_1646);
  xnor csa_tree_add_24_21_groupi_g5802__5115(csa_tree_add_24_21_groupi_n_1764 ,csa_tree_add_24_21_groupi_n_1634 ,csa_tree_add_24_21_groupi_n_1645);
  not csa_tree_add_24_21_groupi_g5804(csa_tree_add_24_21_groupi_n_1744 ,csa_tree_add_24_21_groupi_n_1745);
  not csa_tree_add_24_21_groupi_g5805(csa_tree_add_24_21_groupi_n_1743 ,csa_tree_add_24_21_groupi_n_1742);
  or csa_tree_add_24_21_groupi_g5806__7482(csa_tree_add_24_21_groupi_n_1741 ,csa_tree_add_24_21_groupi_n_1599 ,csa_tree_add_24_21_groupi_n_1666);
  nor csa_tree_add_24_21_groupi_g5807__4733(csa_tree_add_24_21_groupi_n_1740 ,csa_tree_add_24_21_groupi_n_1368 ,csa_tree_add_24_21_groupi_n_1656);
  or csa_tree_add_24_21_groupi_g5808__6161(csa_tree_add_24_21_groupi_n_1739 ,csa_tree_add_24_21_groupi_n_1367 ,csa_tree_add_24_21_groupi_n_1657);
  or csa_tree_add_24_21_groupi_g5809__9315(csa_tree_add_24_21_groupi_n_1738 ,csa_tree_add_24_21_groupi_n_1615 ,csa_tree_add_24_21_groupi_n_1685);
  and csa_tree_add_24_21_groupi_g5810__9945(csa_tree_add_24_21_groupi_n_1737 ,csa_tree_add_24_21_groupi_n_1452 ,csa_tree_add_24_21_groupi_n_1678);
  nor csa_tree_add_24_21_groupi_g5811__2883(csa_tree_add_24_21_groupi_n_1736 ,csa_tree_add_24_21_groupi_n_1462 ,csa_tree_add_24_21_groupi_n_1668);
  or csa_tree_add_24_21_groupi_g5812__2346(csa_tree_add_24_21_groupi_n_1735 ,csa_tree_add_24_21_groupi_n_1663 ,csa_tree_add_24_21_groupi_n_1699);
  or csa_tree_add_24_21_groupi_g5813__1666(csa_tree_add_24_21_groupi_n_1734 ,csa_tree_add_24_21_groupi_n_1614 ,csa_tree_add_24_21_groupi_n_1658);
  nor csa_tree_add_24_21_groupi_g5814__7410(csa_tree_add_24_21_groupi_n_1733 ,csa_tree_add_24_21_groupi_n_1664 ,csa_tree_add_24_21_groupi_n_1698);
  nor csa_tree_add_24_21_groupi_g5815__6417(csa_tree_add_24_21_groupi_n_1732 ,csa_tree_add_24_21_groupi_n_1613 ,csa_tree_add_24_21_groupi_n_1659);
  or csa_tree_add_24_21_groupi_g5816__5477(csa_tree_add_24_21_groupi_n_1731 ,csa_tree_add_24_21_groupi_n_1463 ,csa_tree_add_24_21_groupi_n_1667);
  and csa_tree_add_24_21_groupi_g5817__2398(csa_tree_add_24_21_groupi_n_1753 ,csa_tree_add_24_21_groupi_n_1629 ,csa_tree_add_24_21_groupi_n_1695);
  and csa_tree_add_24_21_groupi_g5818__5107(csa_tree_add_24_21_groupi_n_1752 ,csa_tree_add_24_21_groupi_n_1567 ,csa_tree_add_24_21_groupi_n_1687);
  and csa_tree_add_24_21_groupi_g5819__6260(csa_tree_add_24_21_groupi_n_1751 ,csa_tree_add_24_21_groupi_n_1625 ,csa_tree_add_24_21_groupi_n_1693);
  and csa_tree_add_24_21_groupi_g5820__4319(csa_tree_add_24_21_groupi_n_1750 ,csa_tree_add_24_21_groupi_n_1619 ,csa_tree_add_24_21_groupi_n_1682);
  and csa_tree_add_24_21_groupi_g5821__8428(csa_tree_add_24_21_groupi_n_1749 ,csa_tree_add_24_21_groupi_n_1501 ,csa_tree_add_24_21_groupi_n_1684);
  and csa_tree_add_24_21_groupi_g5822__5526(csa_tree_add_24_21_groupi_n_1748 ,csa_tree_add_24_21_groupi_n_1628 ,csa_tree_add_24_21_groupi_n_1690);
  and csa_tree_add_24_21_groupi_g5823__6783(csa_tree_add_24_21_groupi_n_1747 ,csa_tree_add_24_21_groupi_n_1576 ,csa_tree_add_24_21_groupi_n_1691);
  and csa_tree_add_24_21_groupi_g5824__3680(csa_tree_add_24_21_groupi_n_1746 ,csa_tree_add_24_21_groupi_n_1592 ,csa_tree_add_24_21_groupi_n_1694);
  and csa_tree_add_24_21_groupi_g5825__1617(csa_tree_add_24_21_groupi_n_1745 ,csa_tree_add_24_21_groupi_n_1594 ,csa_tree_add_24_21_groupi_n_1689);
  or csa_tree_add_24_21_groupi_g5826__2802(csa_tree_add_24_21_groupi_n_1742 ,csa_tree_add_24_21_groupi_n_1621 ,csa_tree_add_24_21_groupi_n_1683);
  not csa_tree_add_24_21_groupi_g5827(csa_tree_add_24_21_groupi_n_1729 ,csa_tree_add_24_21_groupi_n_1728);
  not csa_tree_add_24_21_groupi_g5828(csa_tree_add_24_21_groupi_n_1726 ,csa_tree_add_24_21_groupi_n_1727);
  not csa_tree_add_24_21_groupi_g5829(csa_tree_add_24_21_groupi_n_1724 ,csa_tree_add_24_21_groupi_n_1725);
  not csa_tree_add_24_21_groupi_g5830(csa_tree_add_24_21_groupi_n_1722 ,csa_tree_add_24_21_groupi_n_1723);
  not csa_tree_add_24_21_groupi_g5831(csa_tree_add_24_21_groupi_n_1721 ,csa_tree_add_24_21_groupi_n_1720);
  not csa_tree_add_24_21_groupi_g5832(csa_tree_add_24_21_groupi_n_1719 ,csa_tree_add_24_21_groupi_n_1718);
  or csa_tree_add_24_21_groupi_g5833__1705(csa_tree_add_24_21_groupi_n_1717 ,csa_tree_add_24_21_groupi_n_1661 ,csa_tree_add_24_21_groupi_n_1696);
  or csa_tree_add_24_21_groupi_g5834__5122(csa_tree_add_24_21_groupi_n_1716 ,csa_tree_add_24_21_groupi_n_1633 ,csa_tree_add_24_21_groupi_n_1676);
  or csa_tree_add_24_21_groupi_g5835__8246(csa_tree_add_24_21_groupi_n_1715 ,csa_tree_add_24_21_groupi_n_1702 ,csa_tree_add_24_21_groupi_n_1686);
  or csa_tree_add_24_21_groupi_g5836__7098(csa_tree_add_24_21_groupi_n_1714 ,csa_tree_add_24_21_groupi_n_1447 ,csa_tree_add_24_21_groupi_n_1700);
  nor csa_tree_add_24_21_groupi_g5837__6131(csa_tree_add_24_21_groupi_n_1713 ,csa_tree_add_24_21_groupi_n_1632 ,csa_tree_add_24_21_groupi_n_1677);
  nor csa_tree_add_24_21_groupi_g5838__1881(csa_tree_add_24_21_groupi_n_1712 ,csa_tree_add_24_21_groupi_n_1660 ,csa_tree_add_24_21_groupi_n_1697);
  and csa_tree_add_24_21_groupi_g5839__5115(csa_tree_add_24_21_groupi_n_1711 ,csa_tree_add_24_21_groupi_n_1599 ,csa_tree_add_24_21_groupi_n_1666);
  xnor csa_tree_add_24_21_groupi_g5840__7482(csa_tree_add_24_21_groupi_n_1710 ,csa_tree_add_24_21_groupi_n_1472 ,csa_tree_add_24_21_groupi_n_1587);
  xnor csa_tree_add_24_21_groupi_g5841__4733(csa_tree_add_24_21_groupi_n_1709 ,csa_tree_add_24_21_groupi_n_1550 ,csa_tree_add_24_21_groupi_n_1640);
  xnor csa_tree_add_24_21_groupi_g5842__6161(csa_tree_add_24_21_groupi_n_1708 ,csa_tree_add_24_21_groupi_n_1506 ,csa_tree_add_24_21_groupi_n_1607);
  xnor csa_tree_add_24_21_groupi_g5843__9315(csa_tree_add_24_21_groupi_n_1707 ,csa_tree_add_24_21_groupi_n_1637 ,csa_tree_add_24_21_groupi_n_1608);
  xnor csa_tree_add_24_21_groupi_g5844__9945(csa_tree_add_24_21_groupi_n_1706 ,csa_tree_add_24_21_groupi_n_1638 ,csa_tree_add_24_21_groupi_n_1509);
  xnor csa_tree_add_24_21_groupi_g5845__2883(csa_tree_add_24_21_groupi_n_1705 ,csa_tree_add_24_21_groupi_n_1424 ,csa_tree_add_24_21_groupi_n_1601);
  xnor csa_tree_add_24_21_groupi_g5846__2346(csa_tree_add_24_21_groupi_n_1704 ,csa_tree_add_24_21_groupi_n_1552 ,csa_tree_add_24_21_groupi_n_1631);
  xnor csa_tree_add_24_21_groupi_g5847__1666(csa_tree_add_24_21_groupi_n_1703 ,csa_tree_add_24_21_groupi_n_1334 ,csa_tree_add_24_21_groupi_n_1605);
  and csa_tree_add_24_21_groupi_g5848__7410(csa_tree_add_24_21_groupi_n_1730 ,csa_tree_add_24_21_groupi_n_1478 ,csa_tree_add_24_21_groupi_n_1679);
  xnor csa_tree_add_24_21_groupi_g5849__6417(csa_tree_add_24_21_groupi_n_1728 ,csa_tree_add_24_21_groupi_n_1585 ,csa_tree_add_24_21_groupi_n_1589);
  xnor csa_tree_add_24_21_groupi_g5850__5477(csa_tree_add_24_21_groupi_n_1727 ,csa_tree_add_24_21_groupi_n_1617 ,csa_tree_add_24_21_groupi_n_1522);
  xnor csa_tree_add_24_21_groupi_g5851__2398(csa_tree_add_24_21_groupi_n_1725 ,csa_tree_add_24_21_groupi_n_1643 ,csa_tree_add_24_21_groupi_n_1590);
  xnor csa_tree_add_24_21_groupi_g5852__5107(csa_tree_add_24_21_groupi_n_1723 ,csa_tree_add_24_21_groupi_n_1641 ,csa_tree_add_24_21_groupi_n_1591);
  xnor csa_tree_add_24_21_groupi_g5853__6260(csa_tree_add_24_21_groupi_n_1720 ,csa_tree_add_24_21_groupi_n_1642 ,csa_tree_add_24_21_groupi_n_1516);
  xnor csa_tree_add_24_21_groupi_g5854__4319(csa_tree_add_24_21_groupi_n_1718 ,csa_tree_add_24_21_groupi_n_1429 ,csa_tree_add_24_21_groupi_n_1586);
  not csa_tree_add_24_21_groupi_g5855(csa_tree_add_24_21_groupi_n_1698 ,csa_tree_add_24_21_groupi_n_1699);
  not csa_tree_add_24_21_groupi_g5856(csa_tree_add_24_21_groupi_n_1696 ,csa_tree_add_24_21_groupi_n_1697);
  or csa_tree_add_24_21_groupi_g5857__8428(csa_tree_add_24_21_groupi_n_1695 ,csa_tree_add_24_21_groupi_n_1622 ,csa_tree_add_24_21_groupi_n_1638);
  or csa_tree_add_24_21_groupi_g5858__5526(csa_tree_add_24_21_groupi_n_1694 ,csa_tree_add_24_21_groupi_n_1596 ,csa_tree_add_24_21_groupi_n_1636);
  or csa_tree_add_24_21_groupi_g5859__6783(csa_tree_add_24_21_groupi_n_1693 ,csa_tree_add_24_21_groupi_n_1623 ,csa_tree_add_24_21_groupi_n_1634);
  or csa_tree_add_24_21_groupi_g5860__3680(csa_tree_add_24_21_groupi_n_1692 ,csa_tree_add_24_21_groupi_n_1506 ,csa_tree_add_24_21_groupi_n_1606);
  or csa_tree_add_24_21_groupi_g5861__1617(csa_tree_add_24_21_groupi_n_1691 ,csa_tree_add_24_21_groupi_n_1574 ,csa_tree_add_24_21_groupi_n_1641);
  or csa_tree_add_24_21_groupi_g5862__2802(csa_tree_add_24_21_groupi_n_1690 ,csa_tree_add_24_21_groupi_n_1639 ,csa_tree_add_24_21_groupi_n_1627);
  or csa_tree_add_24_21_groupi_g5863__1705(csa_tree_add_24_21_groupi_n_1689 ,csa_tree_add_24_21_groupi_n_1593 ,csa_tree_add_24_21_groupi_n_1644);
  or csa_tree_add_24_21_groupi_g5864__5122(csa_tree_add_24_21_groupi_n_1688 ,csa_tree_add_24_21_groupi_n_1333 ,csa_tree_add_24_21_groupi_n_1604);
  or csa_tree_add_24_21_groupi_g5865__8246(csa_tree_add_24_21_groupi_n_1687 ,csa_tree_add_24_21_groupi_n_1565 ,csa_tree_add_24_21_groupi_n_1643);
  nor csa_tree_add_24_21_groupi_g5866__7098(csa_tree_add_24_21_groupi_n_1686 ,csa_tree_add_24_21_groupi_n_1505 ,csa_tree_add_24_21_groupi_n_1607);
  nor csa_tree_add_24_21_groupi_g5867__6131(csa_tree_add_24_21_groupi_n_1685 ,csa_tree_add_24_21_groupi_n_1334 ,csa_tree_add_24_21_groupi_n_1605);
  or csa_tree_add_24_21_groupi_g5868__1881(csa_tree_add_24_21_groupi_n_1684 ,csa_tree_add_24_21_groupi_n_1496 ,csa_tree_add_24_21_groupi_n_1642);
  nor csa_tree_add_24_21_groupi_g5869__5115(csa_tree_add_24_21_groupi_n_1683 ,csa_tree_add_24_21_groupi_n_1620 ,csa_tree_add_24_21_groupi_n_1616);
  or csa_tree_add_24_21_groupi_g5870__7482(csa_tree_add_24_21_groupi_n_1682 ,csa_tree_add_24_21_groupi_n_1618 ,csa_tree_add_24_21_groupi_n_1635);
  nor csa_tree_add_24_21_groupi_g5871__4733(csa_tree_add_24_21_groupi_n_1681 ,csa_tree_add_24_21_groupi_n_1552 ,csa_tree_add_24_21_groupi_n_1630);
  or csa_tree_add_24_21_groupi_g5872__6161(csa_tree_add_24_21_groupi_n_1680 ,csa_tree_add_24_21_groupi_n_1551 ,csa_tree_add_24_21_groupi_n_1631);
  or csa_tree_add_24_21_groupi_g5873(csa_tree_add_24_21_groupi_n_1679 ,csa_tree_add_24_21_groupi_n_1489 ,csa_tree_add_24_21_groupi_n_1617);
  and csa_tree_add_24_21_groupi_g5874(csa_tree_add_24_21_groupi_n_1702 ,csa_tree_add_24_21_groupi_n_1439 ,csa_tree_add_24_21_groupi_n_1598);
  or csa_tree_add_24_21_groupi_g5875(csa_tree_add_24_21_groupi_n_1701 ,csa_tree_add_24_21_groupi_n_1578 ,csa_tree_add_24_21_groupi_n_1624);
  and csa_tree_add_24_21_groupi_g5876(csa_tree_add_24_21_groupi_n_1700 ,csa_tree_add_24_21_groupi_n_1537 ,csa_tree_add_24_21_groupi_n_1595);
  and csa_tree_add_24_21_groupi_g5877(csa_tree_add_24_21_groupi_n_1699 ,csa_tree_add_24_21_groupi_n_1568 ,csa_tree_add_24_21_groupi_n_1626);
  or csa_tree_add_24_21_groupi_g5878(csa_tree_add_24_21_groupi_n_1697 ,csa_tree_add_24_21_groupi_n_1575 ,csa_tree_add_24_21_groupi_n_1597);
  not csa_tree_add_24_21_groupi_g5879(csa_tree_add_24_21_groupi_n_1676 ,csa_tree_add_24_21_groupi_n_1677);
  not csa_tree_add_24_21_groupi_g5880(csa_tree_add_24_21_groupi_n_1674 ,csa_tree_add_24_21_groupi_n_1675);
  not csa_tree_add_24_21_groupi_g5881(csa_tree_add_24_21_groupi_n_1672 ,csa_tree_add_24_21_groupi_n_1671);
  not csa_tree_add_24_21_groupi_g5882(csa_tree_add_24_21_groupi_n_1669 ,csa_tree_add_24_21_groupi_n_1670);
  not csa_tree_add_24_21_groupi_g5883(csa_tree_add_24_21_groupi_n_1668 ,csa_tree_add_24_21_groupi_n_1667);
  not csa_tree_add_24_21_groupi_g5884(csa_tree_add_24_21_groupi_n_1666 ,csa_tree_add_24_21_groupi_n_1665);
  not csa_tree_add_24_21_groupi_g5885(csa_tree_add_24_21_groupi_n_1663 ,csa_tree_add_24_21_groupi_n_1664);
  not csa_tree_add_24_21_groupi_g5886(csa_tree_add_24_21_groupi_n_1660 ,csa_tree_add_24_21_groupi_n_1661);
  not csa_tree_add_24_21_groupi_g5887(csa_tree_add_24_21_groupi_n_1658 ,csa_tree_add_24_21_groupi_n_1659);
  not csa_tree_add_24_21_groupi_g5888(csa_tree_add_24_21_groupi_n_1656 ,csa_tree_add_24_21_groupi_n_1657);
  not csa_tree_add_24_21_groupi_g5889(csa_tree_add_24_21_groupi_n_1654 ,csa_tree_add_24_21_groupi_n_1655);
  nor csa_tree_add_24_21_groupi_g5890(csa_tree_add_24_21_groupi_n_1653 ,csa_tree_add_24_21_groupi_n_1423 ,csa_tree_add_24_21_groupi_n_1601);
  or csa_tree_add_24_21_groupi_g5891(csa_tree_add_24_21_groupi_n_1652 ,csa_tree_add_24_21_groupi_n_1424 ,csa_tree_add_24_21_groupi_n_1600);
  xnor csa_tree_add_24_21_groupi_g5892(csa_tree_add_24_21_groupi_n_1651 ,csa_tree_add_24_21_groupi_n_1581 ,csa_tree_add_24_21_groupi_n_1366);
  xnor csa_tree_add_24_21_groupi_g5893(csa_tree_add_24_21_groupi_n_1650 ,csa_tree_add_24_21_groupi_n_1419 ,csa_tree_add_24_21_groupi_n_1542);
  xnor csa_tree_add_24_21_groupi_g5894(csa_tree_add_24_21_groupi_n_1649 ,csa_tree_add_24_21_groupi_n_1512 ,csa_tree_add_24_21_groupi_n_1548);
  xnor csa_tree_add_24_21_groupi_g5895(csa_tree_add_24_21_groupi_n_1648 ,csa_tree_add_24_21_groupi_n_1544 ,csa_tree_add_24_21_groupi_n_1458);
  xnor csa_tree_add_24_21_groupi_g5896(csa_tree_add_24_21_groupi_n_1647 ,csa_tree_add_24_21_groupi_n_1471 ,csa_tree_add_24_21_groupi_n_1546);
  xnor csa_tree_add_24_21_groupi_g5897(csa_tree_add_24_21_groupi_n_1646 ,csa_tree_add_24_21_groupi_n_1583 ,csa_tree_add_24_21_groupi_n_1350);
  xnor csa_tree_add_24_21_groupi_g5898(csa_tree_add_24_21_groupi_n_1645 ,csa_tree_add_24_21_groupi_n_1504 ,csa_tree_add_24_21_groupi_n_1540);
  xnor csa_tree_add_24_21_groupi_g5899(csa_tree_add_24_21_groupi_n_1678 ,csa_tree_add_24_21_groupi_n_1179 ,csa_tree_add_24_21_groupi_n_1517);
  xnor csa_tree_add_24_21_groupi_g5900(csa_tree_add_24_21_groupi_n_1677 ,csa_tree_add_24_21_groupi_n_1377 ,csa_tree_add_24_21_groupi_n_1530);
  xnor csa_tree_add_24_21_groupi_g5901(csa_tree_add_24_21_groupi_n_1675 ,csa_tree_add_24_21_groupi_n_1375 ,csa_tree_add_24_21_groupi_n_1528);
  xnor csa_tree_add_24_21_groupi_g5902(csa_tree_add_24_21_groupi_n_1673 ,csa_tree_add_24_21_groupi_n_1406 ,csa_tree_add_24_21_groupi_n_1532);
  xnor csa_tree_add_24_21_groupi_g5903(csa_tree_add_24_21_groupi_n_1671 ,csa_tree_add_24_21_groupi_n_1414 ,csa_tree_add_24_21_groupi_n_1521);
  xnor csa_tree_add_24_21_groupi_g5904(csa_tree_add_24_21_groupi_n_1670 ,csa_tree_add_24_21_groupi_n_1416 ,csa_tree_add_24_21_groupi_n_1523);
  xnor csa_tree_add_24_21_groupi_g5905(csa_tree_add_24_21_groupi_n_1667 ,csa_tree_add_24_21_groupi_n_1582 ,csa_tree_add_24_21_groupi_n_1524);
  xnor csa_tree_add_24_21_groupi_g5906(csa_tree_add_24_21_groupi_n_1665 ,csa_tree_add_24_21_groupi_n_1370 ,csa_tree_add_24_21_groupi_n_1520);
  xnor csa_tree_add_24_21_groupi_g5907(csa_tree_add_24_21_groupi_n_1664 ,csa_tree_add_24_21_groupi_n_1188 ,csa_tree_add_24_21_groupi_n_1525);
  xor csa_tree_add_24_21_groupi_g5908(csa_tree_add_24_21_groupi_n_1662 ,csa_tree_add_24_21_groupi_n_1412 ,csa_tree_add_24_21_groupi_n_1533);
  xnor csa_tree_add_24_21_groupi_g5909(csa_tree_add_24_21_groupi_n_1661 ,csa_tree_add_24_21_groupi_n_1513 ,csa_tree_add_24_21_groupi_n_1519);
  xnor csa_tree_add_24_21_groupi_g5910(csa_tree_add_24_21_groupi_n_1659 ,csa_tree_add_24_21_groupi_n_1514 ,csa_tree_add_24_21_groupi_n_1526);
  xnor csa_tree_add_24_21_groupi_g5911(csa_tree_add_24_21_groupi_n_1657 ,csa_tree_add_24_21_groupi_n_1344 ,csa_tree_add_24_21_groupi_n_1518);
  xnor csa_tree_add_24_21_groupi_g5912(csa_tree_add_24_21_groupi_n_1655 ,csa_tree_add_24_21_groupi_n_1407 ,csa_tree_add_24_21_groupi_n_1515);
  not csa_tree_add_24_21_groupi_g5913(csa_tree_add_24_21_groupi_n_1632 ,csa_tree_add_24_21_groupi_n_1633);
  not csa_tree_add_24_21_groupi_g5914(csa_tree_add_24_21_groupi_n_1631 ,csa_tree_add_24_21_groupi_n_1630);
  or csa_tree_add_24_21_groupi_g5915(csa_tree_add_24_21_groupi_n_1629 ,csa_tree_add_24_21_groupi_n_1509 ,csa_tree_add_24_21_groupi_n_1543);
  or csa_tree_add_24_21_groupi_g5916(csa_tree_add_24_21_groupi_n_1628 ,csa_tree_add_24_21_groupi_n_1512 ,csa_tree_add_24_21_groupi_n_1547);
  nor csa_tree_add_24_21_groupi_g5917(csa_tree_add_24_21_groupi_n_1627 ,csa_tree_add_24_21_groupi_n_1511 ,csa_tree_add_24_21_groupi_n_1548);
  or csa_tree_add_24_21_groupi_g5918(csa_tree_add_24_21_groupi_n_1626 ,csa_tree_add_24_21_groupi_n_1583 ,csa_tree_add_24_21_groupi_n_1566);
  or csa_tree_add_24_21_groupi_g5919(csa_tree_add_24_21_groupi_n_1625 ,csa_tree_add_24_21_groupi_n_1504 ,csa_tree_add_24_21_groupi_n_1539);
  nor csa_tree_add_24_21_groupi_g5920(csa_tree_add_24_21_groupi_n_1624 ,csa_tree_add_24_21_groupi_n_1429 ,csa_tree_add_24_21_groupi_n_1561);
  nor csa_tree_add_24_21_groupi_g5921(csa_tree_add_24_21_groupi_n_1623 ,csa_tree_add_24_21_groupi_n_1503 ,csa_tree_add_24_21_groupi_n_1540);
  and csa_tree_add_24_21_groupi_g5922(csa_tree_add_24_21_groupi_n_1622 ,csa_tree_add_24_21_groupi_n_1509 ,csa_tree_add_24_21_groupi_n_1543);
  nor csa_tree_add_24_21_groupi_g5923(csa_tree_add_24_21_groupi_n_1621 ,csa_tree_add_24_21_groupi_n_1366 ,csa_tree_add_24_21_groupi_n_1581);
  and csa_tree_add_24_21_groupi_g5924(csa_tree_add_24_21_groupi_n_1620 ,csa_tree_add_24_21_groupi_n_1366 ,csa_tree_add_24_21_groupi_n_1581);
  or csa_tree_add_24_21_groupi_g5925(csa_tree_add_24_21_groupi_n_1619 ,csa_tree_add_24_21_groupi_n_1458 ,csa_tree_add_24_21_groupi_n_1544);
  and csa_tree_add_24_21_groupi_g5926(csa_tree_add_24_21_groupi_n_1618 ,csa_tree_add_24_21_groupi_n_1458 ,csa_tree_add_24_21_groupi_n_1544);
  and csa_tree_add_24_21_groupi_g5927(csa_tree_add_24_21_groupi_n_1644 ,csa_tree_add_24_21_groupi_n_1494 ,csa_tree_add_24_21_groupi_n_1577);
  and csa_tree_add_24_21_groupi_g5928(csa_tree_add_24_21_groupi_n_1643 ,csa_tree_add_24_21_groupi_n_1479 ,csa_tree_add_24_21_groupi_n_1563);
  and csa_tree_add_24_21_groupi_g5929(csa_tree_add_24_21_groupi_n_1642 ,csa_tree_add_24_21_groupi_n_1500 ,csa_tree_add_24_21_groupi_n_1553);
  and csa_tree_add_24_21_groupi_g5930(csa_tree_add_24_21_groupi_n_1641 ,csa_tree_add_24_21_groupi_n_1488 ,csa_tree_add_24_21_groupi_n_1573);
  and csa_tree_add_24_21_groupi_g5931(csa_tree_add_24_21_groupi_n_1640 ,csa_tree_add_24_21_groupi_n_1474 ,csa_tree_add_24_21_groupi_n_1560);
  and csa_tree_add_24_21_groupi_g5932(csa_tree_add_24_21_groupi_n_1639 ,csa_tree_add_24_21_groupi_n_1446 ,csa_tree_add_24_21_groupi_n_1572);
  and csa_tree_add_24_21_groupi_g5933(csa_tree_add_24_21_groupi_n_1638 ,csa_tree_add_24_21_groupi_n_1497 ,csa_tree_add_24_21_groupi_n_1556);
  and csa_tree_add_24_21_groupi_g5934(csa_tree_add_24_21_groupi_n_1637 ,csa_tree_add_24_21_groupi_n_1480 ,csa_tree_add_24_21_groupi_n_1564);
  and csa_tree_add_24_21_groupi_g5935(csa_tree_add_24_21_groupi_n_1636 ,csa_tree_add_24_21_groupi_n_1485 ,csa_tree_add_24_21_groupi_n_1570);
  and csa_tree_add_24_21_groupi_g5936(csa_tree_add_24_21_groupi_n_1635 ,csa_tree_add_24_21_groupi_n_1450 ,csa_tree_add_24_21_groupi_n_1554);
  and csa_tree_add_24_21_groupi_g5937(csa_tree_add_24_21_groupi_n_1634 ,csa_tree_add_24_21_groupi_n_1495 ,csa_tree_add_24_21_groupi_n_1562);
  and csa_tree_add_24_21_groupi_g5938(csa_tree_add_24_21_groupi_n_1633 ,csa_tree_add_24_21_groupi_n_1263 ,csa_tree_add_24_21_groupi_n_1555);
  or csa_tree_add_24_21_groupi_g5939(csa_tree_add_24_21_groupi_n_1630 ,csa_tree_add_24_21_groupi_n_1483 ,csa_tree_add_24_21_groupi_n_1559);
  not csa_tree_add_24_21_groupi_g5940(csa_tree_add_24_21_groupi_n_1613 ,csa_tree_add_24_21_groupi_n_1614);
  not csa_tree_add_24_21_groupi_g5941(csa_tree_add_24_21_groupi_n_1612 ,csa_tree_add_24_21_groupi_n_1611);
  not csa_tree_add_24_21_groupi_g5942(csa_tree_add_24_21_groupi_n_1610 ,csa_tree_add_24_21_groupi_n_1609);
  not csa_tree_add_24_21_groupi_g5943(csa_tree_add_24_21_groupi_n_1606 ,csa_tree_add_24_21_groupi_n_1607);
  not csa_tree_add_24_21_groupi_g5944(csa_tree_add_24_21_groupi_n_1605 ,csa_tree_add_24_21_groupi_n_1604);
  not csa_tree_add_24_21_groupi_g5945(csa_tree_add_24_21_groupi_n_1602 ,csa_tree_add_24_21_groupi_n_1603);
  not csa_tree_add_24_21_groupi_g5946(csa_tree_add_24_21_groupi_n_1601 ,csa_tree_add_24_21_groupi_n_1600);
  or csa_tree_add_24_21_groupi_g5947(csa_tree_add_24_21_groupi_n_1598 ,csa_tree_add_24_21_groupi_n_1440 ,csa_tree_add_24_21_groupi_n_1582);
  and csa_tree_add_24_21_groupi_g5948(csa_tree_add_24_21_groupi_n_1597 ,csa_tree_add_24_21_groupi_n_1585 ,csa_tree_add_24_21_groupi_n_1558);
  nor csa_tree_add_24_21_groupi_g5949(csa_tree_add_24_21_groupi_n_1596 ,csa_tree_add_24_21_groupi_n_1419 ,csa_tree_add_24_21_groupi_n_1542);
  or csa_tree_add_24_21_groupi_g5950(csa_tree_add_24_21_groupi_n_1595 ,csa_tree_add_24_21_groupi_n_1472 ,csa_tree_add_24_21_groupi_n_1538);
  or csa_tree_add_24_21_groupi_g5951(csa_tree_add_24_21_groupi_n_1594 ,csa_tree_add_24_21_groupi_n_1470 ,csa_tree_add_24_21_groupi_n_1545);
  nor csa_tree_add_24_21_groupi_g5952(csa_tree_add_24_21_groupi_n_1593 ,csa_tree_add_24_21_groupi_n_1471 ,csa_tree_add_24_21_groupi_n_1546);
  or csa_tree_add_24_21_groupi_g5953(csa_tree_add_24_21_groupi_n_1592 ,csa_tree_add_24_21_groupi_n_1418 ,csa_tree_add_24_21_groupi_n_1541);
  xnor csa_tree_add_24_21_groupi_g5954(csa_tree_add_24_21_groupi_n_1591 ,csa_tree_add_24_21_groupi_n_1508 ,csa_tree_add_24_21_groupi_n_1362);
  xnor csa_tree_add_24_21_groupi_g5955(csa_tree_add_24_21_groupi_n_1590 ,csa_tree_add_24_21_groupi_n_1464 ,csa_tree_add_24_21_groupi_n_1510);
  xnor csa_tree_add_24_21_groupi_g5956(csa_tree_add_24_21_groupi_n_1589 ,csa_tree_add_24_21_groupi_n_1165 ,csa_tree_add_24_21_groupi_n_1467);
  xnor csa_tree_add_24_21_groupi_g5957(csa_tree_add_24_21_groupi_n_1588 ,csa_tree_add_24_21_groupi_n_1373 ,csa_tree_add_24_21_groupi_n_1460);
  xnor csa_tree_add_24_21_groupi_g5958(csa_tree_add_24_21_groupi_n_1587 ,csa_tree_add_24_21_groupi_n_1246 ,csa_tree_add_24_21_groupi_n_1469);
  xnor csa_tree_add_24_21_groupi_g5959(csa_tree_add_24_21_groupi_n_1586 ,csa_tree_add_24_21_groupi_n_1345 ,csa_tree_add_24_21_groupi_n_1461);
  xnor csa_tree_add_24_21_groupi_g5960(csa_tree_add_24_21_groupi_n_1617 ,csa_tree_add_24_21_groupi_n_1285 ,csa_tree_add_24_21_groupi_n_1432);
  xnor csa_tree_add_24_21_groupi_g5961(csa_tree_add_24_21_groupi_n_1616 ,csa_tree_add_24_21_groupi_n_1378 ,csa_tree_add_24_21_groupi_n_1438);
  and csa_tree_add_24_21_groupi_g5962(csa_tree_add_24_21_groupi_n_1615 ,csa_tree_add_24_21_groupi_n_1451 ,csa_tree_add_24_21_groupi_n_1571);
  xnor csa_tree_add_24_21_groupi_g5963(csa_tree_add_24_21_groupi_n_1614 ,csa_tree_add_24_21_groupi_n_1430 ,csa_tree_add_24_21_groupi_n_1434);
  xnor csa_tree_add_24_21_groupi_g5964(csa_tree_add_24_21_groupi_n_1611 ,csa_tree_add_24_21_groupi_n_1376 ,csa_tree_add_24_21_groupi_n_1437);
  xnor csa_tree_add_24_21_groupi_g5965(csa_tree_add_24_21_groupi_n_1609 ,csa_tree_add_24_21_groupi_n_1357 ,csa_tree_add_24_21_groupi_n_1436);
  xnor csa_tree_add_24_21_groupi_g5966(csa_tree_add_24_21_groupi_n_1608 ,csa_tree_add_24_21_groupi_n_1363 ,csa_tree_add_24_21_groupi_n_1435);
  xnor csa_tree_add_24_21_groupi_g5967(csa_tree_add_24_21_groupi_n_1607 ,csa_tree_add_24_21_groupi_n_1404 ,csa_tree_add_24_21_groupi_n_1433);
  xnor csa_tree_add_24_21_groupi_g5968(csa_tree_add_24_21_groupi_n_1604 ,csa_tree_add_24_21_groupi_n_1253 ,csa_tree_add_24_21_groupi_n_1431);
  and csa_tree_add_24_21_groupi_g5969(csa_tree_add_24_21_groupi_n_1603 ,csa_tree_add_24_21_groupi_n_1441 ,csa_tree_add_24_21_groupi_n_1557);
  xnor csa_tree_add_24_21_groupi_g5970(csa_tree_add_24_21_groupi_n_1600 ,csa_tree_add_24_21_groupi_n_1473 ,csa_tree_add_24_21_groupi_n_1322);
  and csa_tree_add_24_21_groupi_g5971(csa_tree_add_24_21_groupi_n_1599 ,csa_tree_add_24_21_groupi_n_1443 ,csa_tree_add_24_21_groupi_n_1569);
  not csa_tree_add_24_21_groupi_g5972(csa_tree_add_24_21_groupi_n_1580 ,csa_tree_add_24_21_groupi_n_1579);
  nor csa_tree_add_24_21_groupi_g5973(csa_tree_add_24_21_groupi_n_1578 ,csa_tree_add_24_21_groupi_n_1461 ,csa_tree_add_24_21_groupi_n_1345);
  or csa_tree_add_24_21_groupi_g5974(csa_tree_add_24_21_groupi_n_1577 ,csa_tree_add_24_21_groupi_n_1312 ,csa_tree_add_24_21_groupi_n_1490);
  or csa_tree_add_24_21_groupi_g5975(csa_tree_add_24_21_groupi_n_1576 ,csa_tree_add_24_21_groupi_n_1508 ,csa_tree_add_24_21_groupi_n_1361);
  nor csa_tree_add_24_21_groupi_g5976(csa_tree_add_24_21_groupi_n_1575 ,csa_tree_add_24_21_groupi_n_1164 ,csa_tree_add_24_21_groupi_n_1467);
  nor csa_tree_add_24_21_groupi_g5977(csa_tree_add_24_21_groupi_n_1574 ,csa_tree_add_24_21_groupi_n_1507 ,csa_tree_add_24_21_groupi_n_1362);
  or csa_tree_add_24_21_groupi_g5978(csa_tree_add_24_21_groupi_n_1573 ,csa_tree_add_24_21_groupi_n_1321 ,csa_tree_add_24_21_groupi_n_1486);
  or csa_tree_add_24_21_groupi_g5979(csa_tree_add_24_21_groupi_n_1572 ,csa_tree_add_24_21_groupi_n_1311 ,csa_tree_add_24_21_groupi_n_1445);
  or csa_tree_add_24_21_groupi_g5980(csa_tree_add_24_21_groupi_n_1571 ,csa_tree_add_24_21_groupi_n_1319 ,csa_tree_add_24_21_groupi_n_1499);
  or csa_tree_add_24_21_groupi_g5981(csa_tree_add_24_21_groupi_n_1570 ,csa_tree_add_24_21_groupi_n_1317 ,csa_tree_add_24_21_groupi_n_1484);
  or csa_tree_add_24_21_groupi_g5982(csa_tree_add_24_21_groupi_n_1569 ,csa_tree_add_24_21_groupi_n_1377 ,csa_tree_add_24_21_groupi_n_1442);
  or csa_tree_add_24_21_groupi_g5983(csa_tree_add_24_21_groupi_n_1568 ,csa_tree_add_24_21_groupi_n_1350 ,csa_tree_add_24_21_groupi_n_1465);
  or csa_tree_add_24_21_groupi_g5984(csa_tree_add_24_21_groupi_n_1567 ,csa_tree_add_24_21_groupi_n_1510 ,csa_tree_add_24_21_groupi_n_1464);
  and csa_tree_add_24_21_groupi_g5985(csa_tree_add_24_21_groupi_n_1566 ,csa_tree_add_24_21_groupi_n_1350 ,csa_tree_add_24_21_groupi_n_1465);
  and csa_tree_add_24_21_groupi_g5986(csa_tree_add_24_21_groupi_n_1565 ,csa_tree_add_24_21_groupi_n_1510 ,csa_tree_add_24_21_groupi_n_1464);
  or csa_tree_add_24_21_groupi_g5987(csa_tree_add_24_21_groupi_n_1564 ,csa_tree_add_24_21_groupi_n_1514 ,csa_tree_add_24_21_groupi_n_1476);
  or csa_tree_add_24_21_groupi_g5988(csa_tree_add_24_21_groupi_n_1563 ,csa_tree_add_24_21_groupi_n_1287 ,csa_tree_add_24_21_groupi_n_1475);
  or csa_tree_add_24_21_groupi_g5989(csa_tree_add_24_21_groupi_n_1562 ,csa_tree_add_24_21_groupi_n_1307 ,csa_tree_add_24_21_groupi_n_1498);
  and csa_tree_add_24_21_groupi_g5990(csa_tree_add_24_21_groupi_n_1561 ,csa_tree_add_24_21_groupi_n_1461 ,csa_tree_add_24_21_groupi_n_1345);
  or csa_tree_add_24_21_groupi_g5991(csa_tree_add_24_21_groupi_n_1560 ,csa_tree_add_24_21_groupi_n_1427 ,csa_tree_add_24_21_groupi_n_1482);
  nor csa_tree_add_24_21_groupi_g5992(csa_tree_add_24_21_groupi_n_1559 ,csa_tree_add_24_21_groupi_n_1491 ,csa_tree_add_24_21_groupi_n_1513);
  or csa_tree_add_24_21_groupi_g5993(csa_tree_add_24_21_groupi_n_1558 ,csa_tree_add_24_21_groupi_n_1165 ,csa_tree_add_24_21_groupi_n_1466);
  or csa_tree_add_24_21_groupi_g5994(csa_tree_add_24_21_groupi_n_1557 ,csa_tree_add_24_21_groupi_n_1288 ,csa_tree_add_24_21_groupi_n_1453);
  or csa_tree_add_24_21_groupi_g5995(csa_tree_add_24_21_groupi_n_1556 ,csa_tree_add_24_21_groupi_n_1283 ,csa_tree_add_24_21_groupi_n_1456);
  or csa_tree_add_24_21_groupi_g5996(csa_tree_add_24_21_groupi_n_1555 ,csa_tree_add_24_21_groupi_n_1264 ,csa_tree_add_24_21_groupi_n_1473);
  or csa_tree_add_24_21_groupi_g5997(csa_tree_add_24_21_groupi_n_1554 ,csa_tree_add_24_21_groupi_n_1284 ,csa_tree_add_24_21_groupi_n_1492);
  or csa_tree_add_24_21_groupi_g5998(csa_tree_add_24_21_groupi_n_1553 ,csa_tree_add_24_21_groupi_n_1315 ,csa_tree_add_24_21_groupi_n_1493);
  or csa_tree_add_24_21_groupi_g5999(csa_tree_add_24_21_groupi_n_1585 ,csa_tree_add_24_21_groupi_n_1393 ,csa_tree_add_24_21_groupi_n_1477);
  and csa_tree_add_24_21_groupi_g6000(csa_tree_add_24_21_groupi_n_1584 ,csa_tree_add_24_21_groupi_n_1379 ,csa_tree_add_24_21_groupi_n_1502);
  and csa_tree_add_24_21_groupi_g6001(csa_tree_add_24_21_groupi_n_1583 ,csa_tree_add_24_21_groupi_n_1389 ,csa_tree_add_24_21_groupi_n_1444);
  and csa_tree_add_24_21_groupi_g6002(csa_tree_add_24_21_groupi_n_1582 ,csa_tree_add_24_21_groupi_n_1390 ,csa_tree_add_24_21_groupi_n_1481);
  and csa_tree_add_24_21_groupi_g6003(csa_tree_add_24_21_groupi_n_1581 ,csa_tree_add_24_21_groupi_n_1273 ,csa_tree_add_24_21_groupi_n_1455);
  or csa_tree_add_24_21_groupi_g6004(csa_tree_add_24_21_groupi_n_1579 ,csa_tree_add_24_21_groupi_n_1382 ,csa_tree_add_24_21_groupi_n_1449);
  not csa_tree_add_24_21_groupi_g6005(csa_tree_add_24_21_groupi_n_1551 ,csa_tree_add_24_21_groupi_n_1552);
  not csa_tree_add_24_21_groupi_g6006(csa_tree_add_24_21_groupi_n_1550 ,csa_tree_add_24_21_groupi_n_1549);
  not csa_tree_add_24_21_groupi_g6007(csa_tree_add_24_21_groupi_n_1548 ,csa_tree_add_24_21_groupi_n_1547);
  not csa_tree_add_24_21_groupi_g6008(csa_tree_add_24_21_groupi_n_1546 ,csa_tree_add_24_21_groupi_n_1545);
  not csa_tree_add_24_21_groupi_g6009(csa_tree_add_24_21_groupi_n_1541 ,csa_tree_add_24_21_groupi_n_1542);
  not csa_tree_add_24_21_groupi_g6010(csa_tree_add_24_21_groupi_n_1539 ,csa_tree_add_24_21_groupi_n_1540);
  nor csa_tree_add_24_21_groupi_g6011(csa_tree_add_24_21_groupi_n_1538 ,csa_tree_add_24_21_groupi_n_1246 ,csa_tree_add_24_21_groupi_n_1468);
  or csa_tree_add_24_21_groupi_g6012(csa_tree_add_24_21_groupi_n_1537 ,csa_tree_add_24_21_groupi_n_1245 ,csa_tree_add_24_21_groupi_n_1469);
  or csa_tree_add_24_21_groupi_g6013(csa_tree_add_24_21_groupi_n_1536 ,csa_tree_add_24_21_groupi_n_1372 ,csa_tree_add_24_21_groupi_n_1460);
  xnor csa_tree_add_24_21_groupi_g6014(csa_tree_add_24_21_groupi_n_1535 ,csa_tree_add_24_21_groupi_n_1251 ,csa_tree_add_24_21_groupi_n_1323);
  nor csa_tree_add_24_21_groupi_g6015(csa_tree_add_24_21_groupi_n_1534 ,csa_tree_add_24_21_groupi_n_1373 ,csa_tree_add_24_21_groupi_n_1459);
  xnor csa_tree_add_24_21_groupi_g6016(csa_tree_add_24_21_groupi_n_1533 ,csa_tree_add_24_21_groupi_n_1347 ,csa_tree_add_24_21_groupi_n_1287);
  xnor csa_tree_add_24_21_groupi_g6017(csa_tree_add_24_21_groupi_n_1532 ,csa_tree_add_24_21_groupi_n_1336 ,csa_tree_add_24_21_groupi_n_1284);
  xnor csa_tree_add_24_21_groupi_g6018(csa_tree_add_24_21_groupi_n_1531 ,csa_tree_add_24_21_groupi_n_1402 ,csa_tree_add_24_21_groupi_n_1343);
  xnor csa_tree_add_24_21_groupi_g6019(csa_tree_add_24_21_groupi_n_1530 ,csa_tree_add_24_21_groupi_n_1181 ,csa_tree_add_24_21_groupi_n_1426);
  xnor csa_tree_add_24_21_groupi_g6020(csa_tree_add_24_21_groupi_n_1529 ,csa_tree_add_24_21_groupi_n_1421 ,csa_tree_add_24_21_groupi_n_1338);
  xnor csa_tree_add_24_21_groupi_g6021(csa_tree_add_24_21_groupi_n_1528 ,csa_tree_add_24_21_groupi_n_1352 ,csa_tree_add_24_21_groupi_n_1321);
  xnor csa_tree_add_24_21_groupi_g6022(csa_tree_add_24_21_groupi_n_1527 ,csa_tree_add_24_21_groupi_n_405 ,csa_tree_add_24_21_groupi_n_1417);
  xnor csa_tree_add_24_21_groupi_g6023(csa_tree_add_24_21_groupi_n_1526 ,csa_tree_add_24_21_groupi_n_1348 ,csa_tree_add_24_21_groupi_n_1349);
  xnor csa_tree_add_24_21_groupi_g6024(csa_tree_add_24_21_groupi_n_1525 ,csa_tree_add_24_21_groupi_n_1354 ,csa_tree_add_24_21_groupi_n_1312);
  xnor csa_tree_add_24_21_groupi_g6025(csa_tree_add_24_21_groupi_n_1524 ,csa_tree_add_24_21_groupi_n_1242 ,csa_tree_add_24_21_groupi_n_1360);
  xnor csa_tree_add_24_21_groupi_g6026(csa_tree_add_24_21_groupi_n_1523 ,csa_tree_add_24_21_groupi_n_1340 ,csa_tree_add_24_21_groupi_n_1307);
  xnor csa_tree_add_24_21_groupi_g6027(csa_tree_add_24_21_groupi_n_1522 ,csa_tree_add_24_21_groupi_n_1177 ,csa_tree_add_24_21_groupi_n_1410);
  xnor csa_tree_add_24_21_groupi_g6028(csa_tree_add_24_21_groupi_n_1521 ,csa_tree_add_24_21_groupi_n_1356 ,csa_tree_add_24_21_groupi_n_1317);
  xnor csa_tree_add_24_21_groupi_g6029(csa_tree_add_24_21_groupi_n_1520 ,csa_tree_add_24_21_groupi_n_1365 ,csa_tree_add_24_21_groupi_n_1288);
  xnor csa_tree_add_24_21_groupi_g6030(csa_tree_add_24_21_groupi_n_1519 ,csa_tree_add_24_21_groupi_n_1247 ,csa_tree_add_24_21_groupi_n_1371);
  xnor csa_tree_add_24_21_groupi_g6031(csa_tree_add_24_21_groupi_n_1518 ,csa_tree_add_24_21_groupi_n_1278 ,csa_tree_add_24_21_groupi_n_1427);
  xnor csa_tree_add_24_21_groupi_g6032(csa_tree_add_24_21_groupi_n_1517 ,csa_tree_add_24_21_groupi_n_1428 ,csa_tree_add_24_21_groupi_n_865);
  xnor csa_tree_add_24_21_groupi_g6033(csa_tree_add_24_21_groupi_n_1516 ,csa_tree_add_24_21_groupi_n_1358 ,csa_tree_add_24_21_groupi_n_1422);
  xnor csa_tree_add_24_21_groupi_g6034(csa_tree_add_24_21_groupi_n_1515 ,csa_tree_add_24_21_groupi_n_1341 ,csa_tree_add_24_21_groupi_n_1283);
  xnor csa_tree_add_24_21_groupi_g6035(csa_tree_add_24_21_groupi_n_1552 ,csa_tree_add_24_21_groupi_n_1320 ,csa_tree_add_24_21_groupi_n_1329);
  xnor csa_tree_add_24_21_groupi_g6036(csa_tree_add_24_21_groupi_n_1549 ,csa_tree_add_24_21_groupi_n_1281 ,csa_tree_add_24_21_groupi_n_1324);
  xnor csa_tree_add_24_21_groupi_g6037(csa_tree_add_24_21_groupi_n_1547 ,csa_tree_add_24_21_groupi_n_1318 ,csa_tree_add_24_21_groupi_n_1327);
  xnor csa_tree_add_24_21_groupi_g6038(csa_tree_add_24_21_groupi_n_1545 ,csa_tree_add_24_21_groupi_n_1123 ,csa_tree_add_24_21_groupi_n_1328);
  xnor csa_tree_add_24_21_groupi_g6039(csa_tree_add_24_21_groupi_n_1544 ,csa_tree_add_24_21_groupi_n_1282 ,csa_tree_add_24_21_groupi_n_1325);
  xnor csa_tree_add_24_21_groupi_g6040(csa_tree_add_24_21_groupi_n_1543 ,csa_tree_add_24_21_groupi_n_1309 ,csa_tree_add_24_21_groupi_n_1331);
  xnor csa_tree_add_24_21_groupi_g6041(csa_tree_add_24_21_groupi_n_1542 ,csa_tree_add_24_21_groupi_n_1308 ,csa_tree_add_24_21_groupi_n_1326);
  xnor csa_tree_add_24_21_groupi_g6042(csa_tree_add_24_21_groupi_n_1540 ,csa_tree_add_24_21_groupi_n_1286 ,csa_tree_add_24_21_groupi_n_1330);
  not csa_tree_add_24_21_groupi_g6043(csa_tree_add_24_21_groupi_n_1511 ,csa_tree_add_24_21_groupi_n_1512);
  not csa_tree_add_24_21_groupi_g6044(csa_tree_add_24_21_groupi_n_1507 ,csa_tree_add_24_21_groupi_n_1508);
  not csa_tree_add_24_21_groupi_g6045(csa_tree_add_24_21_groupi_n_1505 ,csa_tree_add_24_21_groupi_n_1506);
  not csa_tree_add_24_21_groupi_g6046(csa_tree_add_24_21_groupi_n_1503 ,csa_tree_add_24_21_groupi_n_1504);
  or csa_tree_add_24_21_groupi_g6047(csa_tree_add_24_21_groupi_n_1502 ,csa_tree_add_24_21_groupi_n_1380 ,csa_tree_add_24_21_groupi_n_1378);
  or csa_tree_add_24_21_groupi_g6048(csa_tree_add_24_21_groupi_n_1501 ,csa_tree_add_24_21_groupi_n_1422 ,csa_tree_add_24_21_groupi_n_1358);
  or csa_tree_add_24_21_groupi_g6049(csa_tree_add_24_21_groupi_n_1500 ,csa_tree_add_24_21_groupi_n_1302 ,csa_tree_add_24_21_groupi_n_1357);
  nor csa_tree_add_24_21_groupi_g6050(csa_tree_add_24_21_groupi_n_1499 ,csa_tree_add_24_21_groupi_n_1175 ,csa_tree_add_24_21_groupi_n_1404);
  nor csa_tree_add_24_21_groupi_g6051(csa_tree_add_24_21_groupi_n_1498 ,csa_tree_add_24_21_groupi_n_1416 ,csa_tree_add_24_21_groupi_n_1339);
  or csa_tree_add_24_21_groupi_g6052(csa_tree_add_24_21_groupi_n_1497 ,csa_tree_add_24_21_groupi_n_1408 ,csa_tree_add_24_21_groupi_n_1341);
  and csa_tree_add_24_21_groupi_g6053(csa_tree_add_24_21_groupi_n_1496 ,csa_tree_add_24_21_groupi_n_1422 ,csa_tree_add_24_21_groupi_n_1358);
  or csa_tree_add_24_21_groupi_g6054(csa_tree_add_24_21_groupi_n_1495 ,csa_tree_add_24_21_groupi_n_1415 ,csa_tree_add_24_21_groupi_n_1340);
  or csa_tree_add_24_21_groupi_g6055(csa_tree_add_24_21_groupi_n_1494 ,csa_tree_add_24_21_groupi_n_1187 ,csa_tree_add_24_21_groupi_n_1354);
  and csa_tree_add_24_21_groupi_g6056(csa_tree_add_24_21_groupi_n_1493 ,csa_tree_add_24_21_groupi_n_1302 ,csa_tree_add_24_21_groupi_n_1357);
  nor csa_tree_add_24_21_groupi_g6057(csa_tree_add_24_21_groupi_n_1492 ,csa_tree_add_24_21_groupi_n_1406 ,csa_tree_add_24_21_groupi_n_1335);
  nor csa_tree_add_24_21_groupi_g6058(csa_tree_add_24_21_groupi_n_1491 ,csa_tree_add_24_21_groupi_n_1247 ,csa_tree_add_24_21_groupi_n_1371);
  nor csa_tree_add_24_21_groupi_g6059(csa_tree_add_24_21_groupi_n_1490 ,csa_tree_add_24_21_groupi_n_1188 ,csa_tree_add_24_21_groupi_n_1353);
  nor csa_tree_add_24_21_groupi_g6060(csa_tree_add_24_21_groupi_n_1489 ,csa_tree_add_24_21_groupi_n_1176 ,csa_tree_add_24_21_groupi_n_1410);
  or csa_tree_add_24_21_groupi_g6061(csa_tree_add_24_21_groupi_n_1488 ,csa_tree_add_24_21_groupi_n_1374 ,csa_tree_add_24_21_groupi_n_1352);
  and csa_tree_add_24_21_groupi_g6062(csa_tree_add_24_21_groupi_n_1487 ,csa_tree_add_24_21_groupi_n_406 ,csa_tree_add_24_21_groupi_n_1417);
  nor csa_tree_add_24_21_groupi_g6063(csa_tree_add_24_21_groupi_n_1486 ,csa_tree_add_24_21_groupi_n_1375 ,csa_tree_add_24_21_groupi_n_1351);
  or csa_tree_add_24_21_groupi_g6064(csa_tree_add_24_21_groupi_n_1485 ,csa_tree_add_24_21_groupi_n_1413 ,csa_tree_add_24_21_groupi_n_1356);
  nor csa_tree_add_24_21_groupi_g6065(csa_tree_add_24_21_groupi_n_1484 ,csa_tree_add_24_21_groupi_n_1414 ,csa_tree_add_24_21_groupi_n_1355);
  and csa_tree_add_24_21_groupi_g6066(csa_tree_add_24_21_groupi_n_1483 ,csa_tree_add_24_21_groupi_n_1247 ,csa_tree_add_24_21_groupi_n_1371);
  and csa_tree_add_24_21_groupi_g6067(csa_tree_add_24_21_groupi_n_1482 ,csa_tree_add_24_21_groupi_n_1278 ,csa_tree_add_24_21_groupi_n_1344);
  or csa_tree_add_24_21_groupi_g6068(csa_tree_add_24_21_groupi_n_1481 ,csa_tree_add_24_21_groupi_n_1285 ,csa_tree_add_24_21_groupi_n_1384);
  or csa_tree_add_24_21_groupi_g6069(csa_tree_add_24_21_groupi_n_1480 ,csa_tree_add_24_21_groupi_n_1349 ,csa_tree_add_24_21_groupi_n_1348);
  or csa_tree_add_24_21_groupi_g6070(csa_tree_add_24_21_groupi_n_1479 ,csa_tree_add_24_21_groupi_n_1411 ,csa_tree_add_24_21_groupi_n_1347);
  or csa_tree_add_24_21_groupi_g6071(csa_tree_add_24_21_groupi_n_1478 ,csa_tree_add_24_21_groupi_n_1177 ,csa_tree_add_24_21_groupi_n_1409);
  nor csa_tree_add_24_21_groupi_g6072(csa_tree_add_24_21_groupi_n_1477 ,csa_tree_add_24_21_groupi_n_1253 ,csa_tree_add_24_21_groupi_n_1400);
  and csa_tree_add_24_21_groupi_g6073(csa_tree_add_24_21_groupi_n_1476 ,csa_tree_add_24_21_groupi_n_1349 ,csa_tree_add_24_21_groupi_n_1348);
  nor csa_tree_add_24_21_groupi_g6074(csa_tree_add_24_21_groupi_n_1475 ,csa_tree_add_24_21_groupi_n_1412 ,csa_tree_add_24_21_groupi_n_1346);
  or csa_tree_add_24_21_groupi_g6075(csa_tree_add_24_21_groupi_n_1474 ,csa_tree_add_24_21_groupi_n_1278 ,csa_tree_add_24_21_groupi_n_1344);
  and csa_tree_add_24_21_groupi_g6076(csa_tree_add_24_21_groupi_n_1514 ,csa_tree_add_24_21_groupi_n_1275 ,csa_tree_add_24_21_groupi_n_1385);
  and csa_tree_add_24_21_groupi_g6077(csa_tree_add_24_21_groupi_n_1513 ,csa_tree_add_24_21_groupi_n_1035 ,csa_tree_add_24_21_groupi_n_1397);
  and csa_tree_add_24_21_groupi_g6078(csa_tree_add_24_21_groupi_n_1512 ,csa_tree_add_24_21_groupi_n_1078 ,csa_tree_add_24_21_groupi_n_1394);
  and csa_tree_add_24_21_groupi_g6079(csa_tree_add_24_21_groupi_n_1510 ,csa_tree_add_24_21_groupi_n_1296 ,csa_tree_add_24_21_groupi_n_1387);
  and csa_tree_add_24_21_groupi_g6080(csa_tree_add_24_21_groupi_n_1509 ,csa_tree_add_24_21_groupi_n_1270 ,csa_tree_add_24_21_groupi_n_1381);
  and csa_tree_add_24_21_groupi_g6081(csa_tree_add_24_21_groupi_n_1508 ,csa_tree_add_24_21_groupi_n_1226 ,csa_tree_add_24_21_groupi_n_1395);
  and csa_tree_add_24_21_groupi_g6082(csa_tree_add_24_21_groupi_n_1506 ,csa_tree_add_24_21_groupi_n_1092 ,csa_tree_add_24_21_groupi_n_1396);
  and csa_tree_add_24_21_groupi_g6083(csa_tree_add_24_21_groupi_n_1504 ,csa_tree_add_24_21_groupi_n_1297 ,csa_tree_add_24_21_groupi_n_1398);
  not csa_tree_add_24_21_groupi_g6084(csa_tree_add_24_21_groupi_n_1470 ,csa_tree_add_24_21_groupi_n_1471);
  not csa_tree_add_24_21_groupi_g6085(csa_tree_add_24_21_groupi_n_1468 ,csa_tree_add_24_21_groupi_n_1469);
  not csa_tree_add_24_21_groupi_g6086(csa_tree_add_24_21_groupi_n_1466 ,csa_tree_add_24_21_groupi_n_1467);
  not csa_tree_add_24_21_groupi_g6087(csa_tree_add_24_21_groupi_n_1462 ,csa_tree_add_24_21_groupi_n_1463);
  not csa_tree_add_24_21_groupi_g6088(csa_tree_add_24_21_groupi_n_1459 ,csa_tree_add_24_21_groupi_n_1460);
  nor csa_tree_add_24_21_groupi_g6089(csa_tree_add_24_21_groupi_n_1457 ,csa_tree_add_24_21_groupi_n_406 ,csa_tree_add_24_21_groupi_n_1417);
  and csa_tree_add_24_21_groupi_g6090(csa_tree_add_24_21_groupi_n_1456 ,csa_tree_add_24_21_groupi_n_1408 ,csa_tree_add_24_21_groupi_n_1341);
  or csa_tree_add_24_21_groupi_g6091(csa_tree_add_24_21_groupi_n_1455 ,csa_tree_add_24_21_groupi_n_1272 ,csa_tree_add_24_21_groupi_n_1428);
  nor csa_tree_add_24_21_groupi_g6092(csa_tree_add_24_21_groupi_n_1454 ,csa_tree_add_24_21_groupi_n_1420 ,csa_tree_add_24_21_groupi_n_1338);
  nor csa_tree_add_24_21_groupi_g6093(csa_tree_add_24_21_groupi_n_1453 ,csa_tree_add_24_21_groupi_n_1364 ,csa_tree_add_24_21_groupi_n_1370);
  or csa_tree_add_24_21_groupi_g6094(csa_tree_add_24_21_groupi_n_1452 ,csa_tree_add_24_21_groupi_n_1421 ,csa_tree_add_24_21_groupi_n_1337);
  or csa_tree_add_24_21_groupi_g6095(csa_tree_add_24_21_groupi_n_1451 ,csa_tree_add_24_21_groupi_n_1174 ,csa_tree_add_24_21_groupi_n_1403);
  or csa_tree_add_24_21_groupi_g6096(csa_tree_add_24_21_groupi_n_1450 ,csa_tree_add_24_21_groupi_n_1405 ,csa_tree_add_24_21_groupi_n_1336);
  and csa_tree_add_24_21_groupi_g6097(csa_tree_add_24_21_groupi_n_1449 ,csa_tree_add_24_21_groupi_n_1388 ,csa_tree_add_24_21_groupi_n_1376);
  or csa_tree_add_24_21_groupi_g6098(csa_tree_add_24_21_groupi_n_1448 ,csa_tree_add_24_21_groupi_n_1402 ,csa_tree_add_24_21_groupi_n_1342);
  nor csa_tree_add_24_21_groupi_g6099(csa_tree_add_24_21_groupi_n_1447 ,csa_tree_add_24_21_groupi_n_1401 ,csa_tree_add_24_21_groupi_n_1343);
  or csa_tree_add_24_21_groupi_g6100(csa_tree_add_24_21_groupi_n_1446 ,csa_tree_add_24_21_groupi_n_1243 ,csa_tree_add_24_21_groupi_n_1363);
  and csa_tree_add_24_21_groupi_g6101(csa_tree_add_24_21_groupi_n_1445 ,csa_tree_add_24_21_groupi_n_1243 ,csa_tree_add_24_21_groupi_n_1363);
  or csa_tree_add_24_21_groupi_g6102(csa_tree_add_24_21_groupi_n_1444 ,csa_tree_add_24_21_groupi_n_1430 ,csa_tree_add_24_21_groupi_n_1386);
  or csa_tree_add_24_21_groupi_g6103(csa_tree_add_24_21_groupi_n_1443 ,csa_tree_add_24_21_groupi_n_1180 ,csa_tree_add_24_21_groupi_n_1426);
  nor csa_tree_add_24_21_groupi_g6104(csa_tree_add_24_21_groupi_n_1442 ,csa_tree_add_24_21_groupi_n_1181 ,csa_tree_add_24_21_groupi_n_1425);
  or csa_tree_add_24_21_groupi_g6105(csa_tree_add_24_21_groupi_n_1441 ,csa_tree_add_24_21_groupi_n_1365 ,csa_tree_add_24_21_groupi_n_1369);
  nor csa_tree_add_24_21_groupi_g6106(csa_tree_add_24_21_groupi_n_1440 ,csa_tree_add_24_21_groupi_n_1242 ,csa_tree_add_24_21_groupi_n_1360);
  or csa_tree_add_24_21_groupi_g6107(csa_tree_add_24_21_groupi_n_1439 ,csa_tree_add_24_21_groupi_n_1241 ,csa_tree_add_24_21_groupi_n_1359);
  xnor csa_tree_add_24_21_groupi_g6108(csa_tree_add_24_21_groupi_n_1438 ,csa_tree_add_24_21_groupi_n_1277 ,csa_tree_add_24_21_groupi_n_1239);
  xnor csa_tree_add_24_21_groupi_g6109(csa_tree_add_24_21_groupi_n_1437 ,csa_tree_add_24_21_groupi_n_1249 ,csa_tree_add_24_21_groupi_n_1280);
  xnor csa_tree_add_24_21_groupi_g6110(csa_tree_add_24_21_groupi_n_1436 ,csa_tree_add_24_21_groupi_n_1302 ,csa_tree_add_24_21_groupi_n_1315);
  xnor csa_tree_add_24_21_groupi_g6111(csa_tree_add_24_21_groupi_n_1435 ,csa_tree_add_24_21_groupi_n_1311 ,csa_tree_add_24_21_groupi_n_1243);
  xnor csa_tree_add_24_21_groupi_g6112(csa_tree_add_24_21_groupi_n_1434 ,csa_tree_add_24_21_groupi_n_1185 ,csa_tree_add_24_21_groupi_n_1304);
  xor csa_tree_add_24_21_groupi_g6113(csa_tree_add_24_21_groupi_n_1433 ,csa_tree_add_24_21_groupi_n_1175 ,csa_tree_add_24_21_groupi_n_1319);
  xnor csa_tree_add_24_21_groupi_g6114(csa_tree_add_24_21_groupi_n_1432 ,csa_tree_add_24_21_groupi_n_1305 ,csa_tree_add_24_21_groupi_n_985);
  xnor csa_tree_add_24_21_groupi_g6115(csa_tree_add_24_21_groupi_n_1431 ,csa_tree_add_24_21_groupi_n_1306 ,csa_tree_add_24_21_groupi_n_967);
  xnor csa_tree_add_24_21_groupi_g6116(csa_tree_add_24_21_groupi_n_1473 ,csa_tree_add_24_21_groupi_n_918 ,csa_tree_add_24_21_groupi_n_1255);
  and csa_tree_add_24_21_groupi_g6117(csa_tree_add_24_21_groupi_n_1472 ,csa_tree_add_24_21_groupi_n_1289 ,csa_tree_add_24_21_groupi_n_1391);
  or csa_tree_add_24_21_groupi_g6118(csa_tree_add_24_21_groupi_n_1471 ,csa_tree_add_24_21_groupi_n_1301 ,csa_tree_add_24_21_groupi_n_1399);
  xnor csa_tree_add_24_21_groupi_g6119(csa_tree_add_24_21_groupi_n_1469 ,csa_tree_add_24_21_groupi_n_996 ,csa_tree_add_24_21_groupi_n_1258);
  xnor csa_tree_add_24_21_groupi_g6120(csa_tree_add_24_21_groupi_n_1467 ,csa_tree_add_24_21_groupi_n_1310 ,csa_tree_add_24_21_groupi_n_1131);
  xnor csa_tree_add_24_21_groupi_g6121(csa_tree_add_24_21_groupi_n_1465 ,csa_tree_add_24_21_groupi_n_1313 ,csa_tree_add_24_21_groupi_n_1135);
  xnor csa_tree_add_24_21_groupi_g6122(csa_tree_add_24_21_groupi_n_1464 ,csa_tree_add_24_21_groupi_n_1316 ,csa_tree_add_24_21_groupi_n_1256);
  xnor csa_tree_add_24_21_groupi_g6123(csa_tree_add_24_21_groupi_n_1463 ,csa_tree_add_24_21_groupi_n_1314 ,csa_tree_add_24_21_groupi_n_1142);
  xnor csa_tree_add_24_21_groupi_g6124(csa_tree_add_24_21_groupi_n_1461 ,csa_tree_add_24_21_groupi_n_934 ,csa_tree_add_24_21_groupi_n_1257);
  and csa_tree_add_24_21_groupi_g6125(csa_tree_add_24_21_groupi_n_1460 ,csa_tree_add_24_21_groupi_n_1266 ,csa_tree_add_24_21_groupi_n_1392);
  and csa_tree_add_24_21_groupi_g6126(csa_tree_add_24_21_groupi_n_1458 ,csa_tree_add_24_21_groupi_n_1276 ,csa_tree_add_24_21_groupi_n_1383);
  not csa_tree_add_24_21_groupi_g6127(csa_tree_add_24_21_groupi_n_1425 ,csa_tree_add_24_21_groupi_n_1426);
  not csa_tree_add_24_21_groupi_g6128(csa_tree_add_24_21_groupi_n_1424 ,csa_tree_add_24_21_groupi_n_1423);
  not csa_tree_add_24_21_groupi_g6129(csa_tree_add_24_21_groupi_n_1420 ,csa_tree_add_24_21_groupi_n_1421);
  not csa_tree_add_24_21_groupi_g6130(csa_tree_add_24_21_groupi_n_1419 ,csa_tree_add_24_21_groupi_n_1418);
  not csa_tree_add_24_21_groupi_g6131(csa_tree_add_24_21_groupi_n_1415 ,csa_tree_add_24_21_groupi_n_1416);
  not csa_tree_add_24_21_groupi_g6132(csa_tree_add_24_21_groupi_n_1413 ,csa_tree_add_24_21_groupi_n_1414);
  not csa_tree_add_24_21_groupi_g6133(csa_tree_add_24_21_groupi_n_1411 ,csa_tree_add_24_21_groupi_n_1412);
  not csa_tree_add_24_21_groupi_g6134(csa_tree_add_24_21_groupi_n_1409 ,csa_tree_add_24_21_groupi_n_1410);
  not csa_tree_add_24_21_groupi_g6135(csa_tree_add_24_21_groupi_n_1408 ,csa_tree_add_24_21_groupi_n_1407);
  not csa_tree_add_24_21_groupi_g6136(csa_tree_add_24_21_groupi_n_1405 ,csa_tree_add_24_21_groupi_n_1406);
  not csa_tree_add_24_21_groupi_g6137(csa_tree_add_24_21_groupi_n_1403 ,csa_tree_add_24_21_groupi_n_1404);
  not csa_tree_add_24_21_groupi_g6138(csa_tree_add_24_21_groupi_n_1401 ,csa_tree_add_24_21_groupi_n_1402);
  and csa_tree_add_24_21_groupi_g6139(csa_tree_add_24_21_groupi_n_1400 ,csa_tree_add_24_21_groupi_n_967 ,csa_tree_add_24_21_groupi_n_1306);
  and csa_tree_add_24_21_groupi_g6140(csa_tree_add_24_21_groupi_n_1399 ,csa_tree_add_24_21_groupi_n_1318 ,csa_tree_add_24_21_groupi_n_1291);
  or csa_tree_add_24_21_groupi_g6141(csa_tree_add_24_21_groupi_n_1398 ,csa_tree_add_24_21_groupi_n_1295 ,csa_tree_add_24_21_groupi_n_1308);
  or csa_tree_add_24_21_groupi_g6142(csa_tree_add_24_21_groupi_n_1397 ,csa_tree_add_24_21_groupi_n_1054 ,csa_tree_add_24_21_groupi_n_1310);
  or csa_tree_add_24_21_groupi_g6143(csa_tree_add_24_21_groupi_n_1396 ,csa_tree_add_24_21_groupi_n_1032 ,csa_tree_add_24_21_groupi_n_1314);
  or csa_tree_add_24_21_groupi_g6144(csa_tree_add_24_21_groupi_n_1395 ,csa_tree_add_24_21_groupi_n_1225 ,csa_tree_add_24_21_groupi_n_1316);
  or csa_tree_add_24_21_groupi_g6145(csa_tree_add_24_21_groupi_n_1394 ,csa_tree_add_24_21_groupi_n_1077 ,csa_tree_add_24_21_groupi_n_1313);
  nor csa_tree_add_24_21_groupi_g6146(csa_tree_add_24_21_groupi_n_1393 ,csa_tree_add_24_21_groupi_n_967 ,csa_tree_add_24_21_groupi_n_1306);
  or csa_tree_add_24_21_groupi_g6147(csa_tree_add_24_21_groupi_n_1392 ,csa_tree_add_24_21_groupi_n_1320 ,csa_tree_add_24_21_groupi_n_1290);
  or csa_tree_add_24_21_groupi_g6148(csa_tree_add_24_21_groupi_n_1391 ,csa_tree_add_24_21_groupi_n_1251 ,csa_tree_add_24_21_groupi_n_1294);
  or csa_tree_add_24_21_groupi_g6149(csa_tree_add_24_21_groupi_n_1390 ,csa_tree_add_24_21_groupi_n_985 ,csa_tree_add_24_21_groupi_n_1305);
  or csa_tree_add_24_21_groupi_g6150(csa_tree_add_24_21_groupi_n_1389 ,csa_tree_add_24_21_groupi_n_1184 ,csa_tree_add_24_21_groupi_n_1304);
  or csa_tree_add_24_21_groupi_g6151(csa_tree_add_24_21_groupi_n_1388 ,csa_tree_add_24_21_groupi_n_1249 ,csa_tree_add_24_21_groupi_n_1279);
  or csa_tree_add_24_21_groupi_g6152(csa_tree_add_24_21_groupi_n_1387 ,csa_tree_add_24_21_groupi_n_1300 ,csa_tree_add_24_21_groupi_n_1309);
  nor csa_tree_add_24_21_groupi_g6153(csa_tree_add_24_21_groupi_n_1386 ,csa_tree_add_24_21_groupi_n_1185 ,csa_tree_add_24_21_groupi_n_1303);
  or csa_tree_add_24_21_groupi_g6154(csa_tree_add_24_21_groupi_n_1385 ,csa_tree_add_24_21_groupi_n_1274 ,csa_tree_add_24_21_groupi_n_1281);
  and csa_tree_add_24_21_groupi_g6155(csa_tree_add_24_21_groupi_n_1384 ,csa_tree_add_24_21_groupi_n_985 ,csa_tree_add_24_21_groupi_n_1305);
  or csa_tree_add_24_21_groupi_g6156(csa_tree_add_24_21_groupi_n_1383 ,csa_tree_add_24_21_groupi_n_1267 ,csa_tree_add_24_21_groupi_n_1286);
  nor csa_tree_add_24_21_groupi_g6157(csa_tree_add_24_21_groupi_n_1382 ,csa_tree_add_24_21_groupi_n_1248 ,csa_tree_add_24_21_groupi_n_1280);
  or csa_tree_add_24_21_groupi_g6158(csa_tree_add_24_21_groupi_n_1381 ,csa_tree_add_24_21_groupi_n_1268 ,csa_tree_add_24_21_groupi_n_1282);
  and csa_tree_add_24_21_groupi_g6159(csa_tree_add_24_21_groupi_n_1380 ,csa_tree_add_24_21_groupi_n_1239 ,csa_tree_add_24_21_groupi_n_1277);
  or csa_tree_add_24_21_groupi_g6160(csa_tree_add_24_21_groupi_n_1379 ,csa_tree_add_24_21_groupi_n_1239 ,csa_tree_add_24_21_groupi_n_1277);
  and csa_tree_add_24_21_groupi_g6161(csa_tree_add_24_21_groupi_n_1430 ,csa_tree_add_24_21_groupi_n_1209 ,csa_tree_add_24_21_groupi_n_1260);
  and csa_tree_add_24_21_groupi_g6162(csa_tree_add_24_21_groupi_n_1429 ,csa_tree_add_24_21_groupi_n_1064 ,csa_tree_add_24_21_groupi_n_1271);
  and csa_tree_add_24_21_groupi_g6163(csa_tree_add_24_21_groupi_n_1428 ,csa_tree_add_24_21_groupi_n_1201 ,csa_tree_add_24_21_groupi_n_1262);
  and csa_tree_add_24_21_groupi_g6164(csa_tree_add_24_21_groupi_n_1427 ,csa_tree_add_24_21_groupi_n_1234 ,csa_tree_add_24_21_groupi_n_1265);
  and csa_tree_add_24_21_groupi_g6165(csa_tree_add_24_21_groupi_n_1426 ,csa_tree_add_24_21_groupi_n_1220 ,csa_tree_add_24_21_groupi_n_1259);
  or csa_tree_add_24_21_groupi_g6166(csa_tree_add_24_21_groupi_n_1423 ,csa_tree_add_24_21_groupi_n_1031 ,csa_tree_add_24_21_groupi_n_1299);
  and csa_tree_add_24_21_groupi_g6167(csa_tree_add_24_21_groupi_n_1422 ,csa_tree_add_24_21_groupi_n_1100 ,csa_tree_add_24_21_groupi_n_1269);
  or csa_tree_add_24_21_groupi_g6168(csa_tree_add_24_21_groupi_n_1421 ,csa_tree_add_24_21_groupi_n_1026 ,csa_tree_add_24_21_groupi_n_1261);
  and csa_tree_add_24_21_groupi_g6169(csa_tree_add_24_21_groupi_n_1418 ,csa_tree_add_24_21_groupi_n_1216 ,csa_tree_add_24_21_groupi_n_1293);
  and csa_tree_add_24_21_groupi_g6170(csa_tree_add_24_21_groupi_n_1417 ,csa_tree_add_24_21_groupi_n_851 ,csa_tree_add_24_21_groupi_n_1292);
  xnor csa_tree_add_24_21_groupi_g6171(csa_tree_add_24_21_groupi_n_1416 ,csa_tree_add_24_21_groupi_n_899 ,csa_tree_add_24_21_groupi_n_1162);
  xnor csa_tree_add_24_21_groupi_g6172(csa_tree_add_24_21_groupi_n_1414 ,csa_tree_add_24_21_groupi_n_1012 ,csa_tree_add_24_21_groupi_n_1161);
  xnor csa_tree_add_24_21_groupi_g6173(csa_tree_add_24_21_groupi_n_1412 ,csa_tree_add_24_21_groupi_n_977 ,csa_tree_add_24_21_groupi_n_1155);
  xnor csa_tree_add_24_21_groupi_g6174(csa_tree_add_24_21_groupi_n_1410 ,csa_tree_add_24_21_groupi_n_952 ,csa_tree_add_24_21_groupi_n_1144);
  xnor csa_tree_add_24_21_groupi_g6175(csa_tree_add_24_21_groupi_n_1407 ,csa_tree_add_24_21_groupi_n_1000 ,csa_tree_add_24_21_groupi_n_1152);
  xnor csa_tree_add_24_21_groupi_g6176(csa_tree_add_24_21_groupi_n_1406 ,csa_tree_add_24_21_groupi_n_1017 ,csa_tree_add_24_21_groupi_n_1156);
  xnor csa_tree_add_24_21_groupi_g6177(csa_tree_add_24_21_groupi_n_1404 ,csa_tree_add_24_21_groupi_n_1015 ,csa_tree_add_24_21_groupi_n_1154);
  and csa_tree_add_24_21_groupi_g6178(csa_tree_add_24_21_groupi_n_1402 ,csa_tree_add_24_21_groupi_n_1200 ,csa_tree_add_24_21_groupi_n_1298);
  not csa_tree_add_24_21_groupi_g6179(csa_tree_add_24_21_groupi_n_1374 ,csa_tree_add_24_21_groupi_n_1375);
  not csa_tree_add_24_21_groupi_g6180(csa_tree_add_24_21_groupi_n_1373 ,csa_tree_add_24_21_groupi_n_1372);
  not csa_tree_add_24_21_groupi_g6181(csa_tree_add_24_21_groupi_n_1370 ,csa_tree_add_24_21_groupi_n_1369);
  not csa_tree_add_24_21_groupi_g6182(csa_tree_add_24_21_groupi_n_1367 ,csa_tree_add_24_21_groupi_n_1368);
  not csa_tree_add_24_21_groupi_g6183(csa_tree_add_24_21_groupi_n_1364 ,csa_tree_add_24_21_groupi_n_1365);
  not csa_tree_add_24_21_groupi_g6184(csa_tree_add_24_21_groupi_n_1361 ,csa_tree_add_24_21_groupi_n_1362);
  not csa_tree_add_24_21_groupi_g6185(csa_tree_add_24_21_groupi_n_1359 ,csa_tree_add_24_21_groupi_n_1360);
  not csa_tree_add_24_21_groupi_g6186(csa_tree_add_24_21_groupi_n_1355 ,csa_tree_add_24_21_groupi_n_1356);
  not csa_tree_add_24_21_groupi_g6187(csa_tree_add_24_21_groupi_n_1353 ,csa_tree_add_24_21_groupi_n_1354);
  not csa_tree_add_24_21_groupi_g6188(csa_tree_add_24_21_groupi_n_1351 ,csa_tree_add_24_21_groupi_n_1352);
  not csa_tree_add_24_21_groupi_g6189(csa_tree_add_24_21_groupi_n_1346 ,csa_tree_add_24_21_groupi_n_1347);
  not csa_tree_add_24_21_groupi_g6190(csa_tree_add_24_21_groupi_n_1342 ,csa_tree_add_24_21_groupi_n_1343);
  not csa_tree_add_24_21_groupi_g6191(csa_tree_add_24_21_groupi_n_1339 ,csa_tree_add_24_21_groupi_n_1340);
  not csa_tree_add_24_21_groupi_g6192(csa_tree_add_24_21_groupi_n_1337 ,csa_tree_add_24_21_groupi_n_1338);
  not csa_tree_add_24_21_groupi_g6193(csa_tree_add_24_21_groupi_n_1335 ,csa_tree_add_24_21_groupi_n_1336);
  not csa_tree_add_24_21_groupi_g6194(csa_tree_add_24_21_groupi_n_1333 ,csa_tree_add_24_21_groupi_n_1334);
  xnor csa_tree_add_24_21_groupi_g6195(csa_tree_add_24_21_groupi_n_1332 ,csa_tree_add_24_21_groupi_n_1149 ,csa_tree_add_24_21_groupi_n_481);
  xnor csa_tree_add_24_21_groupi_g6196(csa_tree_add_24_21_groupi_n_1331 ,csa_tree_add_24_21_groupi_n_1240 ,csa_tree_add_24_21_groupi_n_1066);
  xnor csa_tree_add_24_21_groupi_g6197(csa_tree_add_24_21_groupi_n_1330 ,csa_tree_add_24_21_groupi_n_1121 ,csa_tree_add_24_21_groupi_n_1173);
  xnor csa_tree_add_24_21_groupi_g6198(csa_tree_add_24_21_groupi_n_1329 ,csa_tree_add_24_21_groupi_n_867 ,csa_tree_add_24_21_groupi_n_1171);
  xnor csa_tree_add_24_21_groupi_g6199(csa_tree_add_24_21_groupi_n_1328 ,csa_tree_add_24_21_groupi_n_1116 ,csa_tree_add_24_21_groupi_n_1189);
  xnor csa_tree_add_24_21_groupi_g6200(csa_tree_add_24_21_groupi_n_1327 ,csa_tree_add_24_21_groupi_n_983 ,csa_tree_add_24_21_groupi_n_1169);
  xnor csa_tree_add_24_21_groupi_g6201(csa_tree_add_24_21_groupi_n_1326 ,csa_tree_add_24_21_groupi_n_1118 ,csa_tree_add_24_21_groupi_n_1167);
  xnor csa_tree_add_24_21_groupi_g6202(csa_tree_add_24_21_groupi_n_1325 ,csa_tree_add_24_21_groupi_n_1186 ,csa_tree_add_24_21_groupi_n_1119);
  xnor csa_tree_add_24_21_groupi_g6203(csa_tree_add_24_21_groupi_n_1324 ,csa_tree_add_24_21_groupi_n_1250 ,csa_tree_add_24_21_groupi_n_935);
  xnor csa_tree_add_24_21_groupi_g6204(csa_tree_add_24_21_groupi_n_1323 ,csa_tree_add_24_21_groupi_n_688 ,csa_tree_add_24_21_groupi_n_1183);
  xnor csa_tree_add_24_21_groupi_g6205(csa_tree_add_24_21_groupi_n_1322 ,csa_tree_add_24_21_groupi_n_953 ,csa_tree_add_24_21_groupi_n_1244);
  xnor csa_tree_add_24_21_groupi_g6206(csa_tree_add_24_21_groupi_n_1378 ,csa_tree_add_24_21_groupi_n_915 ,csa_tree_add_24_21_groupi_n_1129);
  xnor csa_tree_add_24_21_groupi_g6207(csa_tree_add_24_21_groupi_n_1377 ,csa_tree_add_24_21_groupi_n_890 ,csa_tree_add_24_21_groupi_n_1133);
  xnor csa_tree_add_24_21_groupi_g6208(csa_tree_add_24_21_groupi_n_1376 ,csa_tree_add_24_21_groupi_n_937 ,csa_tree_add_24_21_groupi_n_1138);
  xnor csa_tree_add_24_21_groupi_g6209(csa_tree_add_24_21_groupi_n_1375 ,csa_tree_add_24_21_groupi_n_889 ,csa_tree_add_24_21_groupi_n_1158);
  xnor csa_tree_add_24_21_groupi_g6210(csa_tree_add_24_21_groupi_n_1372 ,csa_tree_add_24_21_groupi_n_1254 ,csa_tree_add_24_21_groupi_n_1021);
  xnor csa_tree_add_24_21_groupi_g6211(csa_tree_add_24_21_groupi_n_1371 ,csa_tree_add_24_21_groupi_n_900 ,csa_tree_add_24_21_groupi_n_1153);
  xnor csa_tree_add_24_21_groupi_g6212(csa_tree_add_24_21_groupi_n_1369 ,csa_tree_add_24_21_groupi_n_1252 ,csa_tree_add_24_21_groupi_n_1136);
  xnor csa_tree_add_24_21_groupi_g6213(csa_tree_add_24_21_groupi_n_1368 ,csa_tree_add_24_21_groupi_n_1192 ,csa_tree_add_24_21_groupi_n_1163);
  xnor csa_tree_add_24_21_groupi_g6214(csa_tree_add_24_21_groupi_n_1366 ,csa_tree_add_24_21_groupi_n_1069 ,csa_tree_add_24_21_groupi_n_1147);
  xnor csa_tree_add_24_21_groupi_g6215(csa_tree_add_24_21_groupi_n_1365 ,csa_tree_add_24_21_groupi_n_1067 ,csa_tree_add_24_21_groupi_n_1150);
  xnor csa_tree_add_24_21_groupi_g6216(csa_tree_add_24_21_groupi_n_1363 ,csa_tree_add_24_21_groupi_n_980 ,csa_tree_add_24_21_groupi_n_1146);
  xnor csa_tree_add_24_21_groupi_g6217(csa_tree_add_24_21_groupi_n_1362 ,csa_tree_add_24_21_groupi_n_1191 ,csa_tree_add_24_21_groupi_n_1159);
  xnor csa_tree_add_24_21_groupi_g6218(csa_tree_add_24_21_groupi_n_1360 ,csa_tree_add_24_21_groupi_n_901 ,csa_tree_add_24_21_groupi_n_1157);
  xnor csa_tree_add_24_21_groupi_g6219(csa_tree_add_24_21_groupi_n_1358 ,csa_tree_add_24_21_groupi_n_964 ,csa_tree_add_24_21_groupi_n_1127);
  xnor csa_tree_add_24_21_groupi_g6220(csa_tree_add_24_21_groupi_n_1357 ,csa_tree_add_24_21_groupi_n_1008 ,csa_tree_add_24_21_groupi_n_1126);
  xnor csa_tree_add_24_21_groupi_g6221(csa_tree_add_24_21_groupi_n_1356 ,csa_tree_add_24_21_groupi_n_1019 ,csa_tree_add_24_21_groupi_n_1125);
  xnor csa_tree_add_24_21_groupi_g6222(csa_tree_add_24_21_groupi_n_1354 ,csa_tree_add_24_21_groupi_n_929 ,csa_tree_add_24_21_groupi_n_1124);
  xnor csa_tree_add_24_21_groupi_g6223(csa_tree_add_24_21_groupi_n_1352 ,csa_tree_add_24_21_groupi_n_939 ,csa_tree_add_24_21_groupi_n_1128);
  xnor csa_tree_add_24_21_groupi_g6224(csa_tree_add_24_21_groupi_n_1350 ,csa_tree_add_24_21_groupi_n_1014 ,csa_tree_add_24_21_groupi_n_1132);
  xnor csa_tree_add_24_21_groupi_g6225(csa_tree_add_24_21_groupi_n_1349 ,csa_tree_add_24_21_groupi_n_1010 ,csa_tree_add_24_21_groupi_n_1137);
  xnor csa_tree_add_24_21_groupi_g6226(csa_tree_add_24_21_groupi_n_1348 ,csa_tree_add_24_21_groupi_n_912 ,csa_tree_add_24_21_groupi_n_1130);
  xnor csa_tree_add_24_21_groupi_g6227(csa_tree_add_24_21_groupi_n_1347 ,csa_tree_add_24_21_groupi_n_969 ,csa_tree_add_24_21_groupi_n_1140);
  xnor csa_tree_add_24_21_groupi_g6228(csa_tree_add_24_21_groupi_n_1345 ,csa_tree_add_24_21_groupi_n_1005 ,csa_tree_add_24_21_groupi_n_1141);
  xnor csa_tree_add_24_21_groupi_g6229(csa_tree_add_24_21_groupi_n_1344 ,csa_tree_add_24_21_groupi_n_970 ,csa_tree_add_24_21_groupi_n_1143);
  xnor csa_tree_add_24_21_groupi_g6230(csa_tree_add_24_21_groupi_n_1343 ,csa_tree_add_24_21_groupi_n_1194 ,csa_tree_add_24_21_groupi_n_1134);
  xnor csa_tree_add_24_21_groupi_g6231(csa_tree_add_24_21_groupi_n_1341 ,csa_tree_add_24_21_groupi_n_854 ,csa_tree_add_24_21_groupi_n_1145);
  xnor csa_tree_add_24_21_groupi_g6232(csa_tree_add_24_21_groupi_n_1340 ,csa_tree_add_24_21_groupi_n_895 ,csa_tree_add_24_21_groupi_n_1139);
  xnor csa_tree_add_24_21_groupi_g6233(csa_tree_add_24_21_groupi_n_1338 ,csa_tree_add_24_21_groupi_n_963 ,csa_tree_add_24_21_groupi_n_1148);
  xnor csa_tree_add_24_21_groupi_g6234(csa_tree_add_24_21_groupi_n_1336 ,csa_tree_add_24_21_groupi_n_948 ,csa_tree_add_24_21_groupi_n_1160);
  xnor csa_tree_add_24_21_groupi_g6235(csa_tree_add_24_21_groupi_n_1334 ,csa_tree_add_24_21_groupi_n_902 ,csa_tree_add_24_21_groupi_n_1151);
  not csa_tree_add_24_21_groupi_g6236(csa_tree_add_24_21_groupi_n_1303 ,csa_tree_add_24_21_groupi_n_1304);
  nor csa_tree_add_24_21_groupi_g6237(csa_tree_add_24_21_groupi_n_1301 ,csa_tree_add_24_21_groupi_n_983 ,csa_tree_add_24_21_groupi_n_1168);
  and csa_tree_add_24_21_groupi_g6238(csa_tree_add_24_21_groupi_n_1300 ,csa_tree_add_24_21_groupi_n_1066 ,csa_tree_add_24_21_groupi_n_1240);
  and csa_tree_add_24_21_groupi_g6239(csa_tree_add_24_21_groupi_n_1299 ,csa_tree_add_24_21_groupi_n_1099 ,csa_tree_add_24_21_groupi_n_1194);
  or csa_tree_add_24_21_groupi_g6240(csa_tree_add_24_21_groupi_n_1298 ,csa_tree_add_24_21_groupi_n_905 ,csa_tree_add_24_21_groupi_n_1237);
  or csa_tree_add_24_21_groupi_g6241(csa_tree_add_24_21_groupi_n_1297 ,csa_tree_add_24_21_groupi_n_1118 ,csa_tree_add_24_21_groupi_n_1166);
  or csa_tree_add_24_21_groupi_g6242(csa_tree_add_24_21_groupi_n_1296 ,csa_tree_add_24_21_groupi_n_1066 ,csa_tree_add_24_21_groupi_n_1240);
  nor csa_tree_add_24_21_groupi_g6243(csa_tree_add_24_21_groupi_n_1295 ,csa_tree_add_24_21_groupi_n_1117 ,csa_tree_add_24_21_groupi_n_1167);
  nor csa_tree_add_24_21_groupi_g6244(csa_tree_add_24_21_groupi_n_1294 ,csa_tree_add_24_21_groupi_n_687 ,csa_tree_add_24_21_groupi_n_1183);
  or csa_tree_add_24_21_groupi_g6245(csa_tree_add_24_21_groupi_n_1293 ,csa_tree_add_24_21_groupi_n_1190 ,csa_tree_add_24_21_groupi_n_1215);
  or csa_tree_add_24_21_groupi_g6246(csa_tree_add_24_21_groupi_n_1292 ,csa_tree_add_24_21_groupi_n_933 ,csa_tree_add_24_21_groupi_n_1254);
  or csa_tree_add_24_21_groupi_g6247(csa_tree_add_24_21_groupi_n_1291 ,csa_tree_add_24_21_groupi_n_982 ,csa_tree_add_24_21_groupi_n_1169);
  nor csa_tree_add_24_21_groupi_g6248(csa_tree_add_24_21_groupi_n_1290 ,csa_tree_add_24_21_groupi_n_867 ,csa_tree_add_24_21_groupi_n_1170);
  or csa_tree_add_24_21_groupi_g6249(csa_tree_add_24_21_groupi_n_1289 ,csa_tree_add_24_21_groupi_n_688 ,csa_tree_add_24_21_groupi_n_1182);
  and csa_tree_add_24_21_groupi_g6250(csa_tree_add_24_21_groupi_n_1321 ,csa_tree_add_24_21_groupi_n_1103 ,csa_tree_add_24_21_groupi_n_1218);
  and csa_tree_add_24_21_groupi_g6251(csa_tree_add_24_21_groupi_n_1320 ,csa_tree_add_24_21_groupi_n_1107 ,csa_tree_add_24_21_groupi_n_1196);
  and csa_tree_add_24_21_groupi_g6252(csa_tree_add_24_21_groupi_n_1319 ,csa_tree_add_24_21_groupi_n_1109 ,csa_tree_add_24_21_groupi_n_1210);
  or csa_tree_add_24_21_groupi_g6253(csa_tree_add_24_21_groupi_n_1318 ,csa_tree_add_24_21_groupi_n_1082 ,csa_tree_add_24_21_groupi_n_1224);
  and csa_tree_add_24_21_groupi_g6254(csa_tree_add_24_21_groupi_n_1317 ,csa_tree_add_24_21_groupi_n_1089 ,csa_tree_add_24_21_groupi_n_1229);
  and csa_tree_add_24_21_groupi_g6255(csa_tree_add_24_21_groupi_n_1316 ,csa_tree_add_24_21_groupi_n_1080 ,csa_tree_add_24_21_groupi_n_1223);
  and csa_tree_add_24_21_groupi_g6256(csa_tree_add_24_21_groupi_n_1315 ,csa_tree_add_24_21_groupi_n_1027 ,csa_tree_add_24_21_groupi_n_1230);
  and csa_tree_add_24_21_groupi_g6257(csa_tree_add_24_21_groupi_n_1314 ,csa_tree_add_24_21_groupi_n_1088 ,csa_tree_add_24_21_groupi_n_1227);
  and csa_tree_add_24_21_groupi_g6258(csa_tree_add_24_21_groupi_n_1313 ,csa_tree_add_24_21_groupi_n_1076 ,csa_tree_add_24_21_groupi_n_1221);
  and csa_tree_add_24_21_groupi_g6259(csa_tree_add_24_21_groupi_n_1312 ,csa_tree_add_24_21_groupi_n_1085 ,csa_tree_add_24_21_groupi_n_1228);
  and csa_tree_add_24_21_groupi_g6260(csa_tree_add_24_21_groupi_n_1311 ,csa_tree_add_24_21_groupi_n_1050 ,csa_tree_add_24_21_groupi_n_1219);
  and csa_tree_add_24_21_groupi_g6261(csa_tree_add_24_21_groupi_n_1310 ,csa_tree_add_24_21_groupi_n_1112 ,csa_tree_add_24_21_groupi_n_1232);
  and csa_tree_add_24_21_groupi_g6262(csa_tree_add_24_21_groupi_n_1309 ,csa_tree_add_24_21_groupi_n_1056 ,csa_tree_add_24_21_groupi_n_1207);
  and csa_tree_add_24_21_groupi_g6263(csa_tree_add_24_21_groupi_n_1308 ,csa_tree_add_24_21_groupi_n_1102 ,csa_tree_add_24_21_groupi_n_1235);
  and csa_tree_add_24_21_groupi_g6264(csa_tree_add_24_21_groupi_n_1307 ,csa_tree_add_24_21_groupi_n_1104 ,csa_tree_add_24_21_groupi_n_1231);
  and csa_tree_add_24_21_groupi_g6265(csa_tree_add_24_21_groupi_n_1306 ,csa_tree_add_24_21_groupi_n_1061 ,csa_tree_add_24_21_groupi_n_1206);
  and csa_tree_add_24_21_groupi_g6266(csa_tree_add_24_21_groupi_n_1305 ,csa_tree_add_24_21_groupi_n_1060 ,csa_tree_add_24_21_groupi_n_1211);
  and csa_tree_add_24_21_groupi_g6267(csa_tree_add_24_21_groupi_n_1304 ,csa_tree_add_24_21_groupi_n_1059 ,csa_tree_add_24_21_groupi_n_1238);
  and csa_tree_add_24_21_groupi_g6268(csa_tree_add_24_21_groupi_n_1302 ,csa_tree_add_24_21_groupi_n_1029 ,csa_tree_add_24_21_groupi_n_1233);
  not csa_tree_add_24_21_groupi_g6269(csa_tree_add_24_21_groupi_n_1279 ,csa_tree_add_24_21_groupi_n_1280);
  or csa_tree_add_24_21_groupi_g6270(csa_tree_add_24_21_groupi_n_1276 ,csa_tree_add_24_21_groupi_n_1121 ,csa_tree_add_24_21_groupi_n_1172);
  or csa_tree_add_24_21_groupi_g6271(csa_tree_add_24_21_groupi_n_1275 ,csa_tree_add_24_21_groupi_n_935 ,csa_tree_add_24_21_groupi_n_1250);
  and csa_tree_add_24_21_groupi_g6272(csa_tree_add_24_21_groupi_n_1274 ,csa_tree_add_24_21_groupi_n_935 ,csa_tree_add_24_21_groupi_n_1250);
  or csa_tree_add_24_21_groupi_g6273(csa_tree_add_24_21_groupi_n_1273 ,csa_tree_add_24_21_groupi_n_865 ,csa_tree_add_24_21_groupi_n_1178);
  nor csa_tree_add_24_21_groupi_g6274(csa_tree_add_24_21_groupi_n_1272 ,csa_tree_add_24_21_groupi_n_864 ,csa_tree_add_24_21_groupi_n_1179);
  or csa_tree_add_24_21_groupi_g6275(csa_tree_add_24_21_groupi_n_1271 ,csa_tree_add_24_21_groupi_n_1038 ,csa_tree_add_24_21_groupi_n_1193);
  or csa_tree_add_24_21_groupi_g6276(csa_tree_add_24_21_groupi_n_1270 ,csa_tree_add_24_21_groupi_n_1119 ,csa_tree_add_24_21_groupi_n_1186);
  or csa_tree_add_24_21_groupi_g6277(csa_tree_add_24_21_groupi_n_1269 ,csa_tree_add_24_21_groupi_n_1097 ,csa_tree_add_24_21_groupi_n_1191);
  and csa_tree_add_24_21_groupi_g6278(csa_tree_add_24_21_groupi_n_1268 ,csa_tree_add_24_21_groupi_n_1119 ,csa_tree_add_24_21_groupi_n_1186);
  nor csa_tree_add_24_21_groupi_g6279(csa_tree_add_24_21_groupi_n_1267 ,csa_tree_add_24_21_groupi_n_1120 ,csa_tree_add_24_21_groupi_n_1173);
  or csa_tree_add_24_21_groupi_g6280(csa_tree_add_24_21_groupi_n_1266 ,csa_tree_add_24_21_groupi_n_866 ,csa_tree_add_24_21_groupi_n_1171);
  or csa_tree_add_24_21_groupi_g6281(csa_tree_add_24_21_groupi_n_1265 ,csa_tree_add_24_21_groupi_n_919 ,csa_tree_add_24_21_groupi_n_1197);
  and csa_tree_add_24_21_groupi_g6282(csa_tree_add_24_21_groupi_n_1264 ,csa_tree_add_24_21_groupi_n_1244 ,csa_tree_add_24_21_groupi_n_953);
  or csa_tree_add_24_21_groupi_g6283(csa_tree_add_24_21_groupi_n_1263 ,csa_tree_add_24_21_groupi_n_1244 ,csa_tree_add_24_21_groupi_n_953);
  or csa_tree_add_24_21_groupi_g6284(csa_tree_add_24_21_groupi_n_1262 ,csa_tree_add_24_21_groupi_n_911 ,csa_tree_add_24_21_groupi_n_1203);
  nor csa_tree_add_24_21_groupi_g6285(csa_tree_add_24_21_groupi_n_1261 ,csa_tree_add_24_21_groupi_n_1252 ,csa_tree_add_24_21_groupi_n_1095);
  or csa_tree_add_24_21_groupi_g6286(csa_tree_add_24_21_groupi_n_1260 ,csa_tree_add_24_21_groupi_n_917 ,csa_tree_add_24_21_groupi_n_1208);
  or csa_tree_add_24_21_groupi_g6287(csa_tree_add_24_21_groupi_n_1259 ,csa_tree_add_24_21_groupi_n_918 ,csa_tree_add_24_21_groupi_n_1217);
  xnor csa_tree_add_24_21_groupi_g6288(csa_tree_add_24_21_groupi_n_1258 ,csa_tree_add_24_21_groupi_n_905 ,csa_tree_add_24_21_groupi_n_1070);
  xnor csa_tree_add_24_21_groupi_g6289(csa_tree_add_24_21_groupi_n_1257 ,csa_tree_add_24_21_groupi_n_917 ,csa_tree_add_24_21_groupi_n_1065);
  xnor csa_tree_add_24_21_groupi_g6290(csa_tree_add_24_21_groupi_n_1256 ,csa_tree_add_24_21_groupi_n_984 ,csa_tree_add_24_21_groupi_n_1114);
  xnor csa_tree_add_24_21_groupi_g6291(csa_tree_add_24_21_groupi_n_1255 ,csa_tree_add_24_21_groupi_n_882 ,csa_tree_add_24_21_groupi_n_1068);
  and csa_tree_add_24_21_groupi_g6292(csa_tree_add_24_21_groupi_n_1288 ,csa_tree_add_24_21_groupi_n_1023 ,csa_tree_add_24_21_groupi_n_1213);
  and csa_tree_add_24_21_groupi_g6293(csa_tree_add_24_21_groupi_n_1287 ,csa_tree_add_24_21_groupi_n_1046 ,csa_tree_add_24_21_groupi_n_1202);
  and csa_tree_add_24_21_groupi_g6294(csa_tree_add_24_21_groupi_n_1286 ,csa_tree_add_24_21_groupi_n_1024 ,csa_tree_add_24_21_groupi_n_1212);
  and csa_tree_add_24_21_groupi_g6295(csa_tree_add_24_21_groupi_n_1285 ,csa_tree_add_24_21_groupi_n_1053 ,csa_tree_add_24_21_groupi_n_1236);
  and csa_tree_add_24_21_groupi_g6296(csa_tree_add_24_21_groupi_n_1284 ,csa_tree_add_24_21_groupi_n_1086 ,csa_tree_add_24_21_groupi_n_1222);
  and csa_tree_add_24_21_groupi_g6297(csa_tree_add_24_21_groupi_n_1283 ,csa_tree_add_24_21_groupi_n_1093 ,csa_tree_add_24_21_groupi_n_1205);
  and csa_tree_add_24_21_groupi_g6298(csa_tree_add_24_21_groupi_n_1282 ,csa_tree_add_24_21_groupi_n_1079 ,csa_tree_add_24_21_groupi_n_1198);
  and csa_tree_add_24_21_groupi_g6299(csa_tree_add_24_21_groupi_n_1281 ,csa_tree_add_24_21_groupi_n_1048 ,csa_tree_add_24_21_groupi_n_1204);
  and csa_tree_add_24_21_groupi_g6300(csa_tree_add_24_21_groupi_n_1280 ,csa_tree_add_24_21_groupi_n_1043 ,csa_tree_add_24_21_groupi_n_1214);
  and csa_tree_add_24_21_groupi_g6301(csa_tree_add_24_21_groupi_n_1278 ,csa_tree_add_24_21_groupi_n_1037 ,csa_tree_add_24_21_groupi_n_1199);
  and csa_tree_add_24_21_groupi_g6302(csa_tree_add_24_21_groupi_n_1277 ,csa_tree_add_24_21_groupi_n_1113 ,csa_tree_add_24_21_groupi_n_1195);
  not csa_tree_add_24_21_groupi_g6303(csa_tree_add_24_21_groupi_n_1249 ,csa_tree_add_24_21_groupi_n_1248);
  not csa_tree_add_24_21_groupi_g6304(csa_tree_add_24_21_groupi_n_1246 ,csa_tree_add_24_21_groupi_n_1245);
  not csa_tree_add_24_21_groupi_g6305(csa_tree_add_24_21_groupi_n_1242 ,csa_tree_add_24_21_groupi_n_1241);
  or csa_tree_add_24_21_groupi_g6306(csa_tree_add_24_21_groupi_n_1238 ,csa_tree_add_24_21_groupi_n_1005 ,csa_tree_add_24_21_groupi_n_1057);
  and csa_tree_add_24_21_groupi_g6307(csa_tree_add_24_21_groupi_n_1237 ,csa_tree_add_24_21_groupi_n_1070 ,csa_tree_add_24_21_groupi_n_996);
  or csa_tree_add_24_21_groupi_g6308(csa_tree_add_24_21_groupi_n_1236 ,csa_tree_add_24_21_groupi_n_903 ,csa_tree_add_24_21_groupi_n_1045);
  or csa_tree_add_24_21_groupi_g6309(csa_tree_add_24_21_groupi_n_1235 ,csa_tree_add_24_21_groupi_n_1012 ,csa_tree_add_24_21_groupi_n_1087);
  or csa_tree_add_24_21_groupi_g6310(csa_tree_add_24_21_groupi_n_1234 ,csa_tree_add_24_21_groupi_n_1069 ,csa_tree_add_24_21_groupi_n_973);
  or csa_tree_add_24_21_groupi_g6311(csa_tree_add_24_21_groupi_n_1233 ,csa_tree_add_24_21_groupi_n_999 ,csa_tree_add_24_21_groupi_n_1062);
  or csa_tree_add_24_21_groupi_g6312(csa_tree_add_24_21_groupi_n_1232 ,csa_tree_add_24_21_groupi_n_1110 ,csa_tree_add_24_21_groupi_n_902);
  or csa_tree_add_24_21_groupi_g6313(csa_tree_add_24_21_groupi_n_1231 ,csa_tree_add_24_21_groupi_n_1019 ,csa_tree_add_24_21_groupi_n_1091);
  or csa_tree_add_24_21_groupi_g6314(csa_tree_add_24_21_groupi_n_1230 ,csa_tree_add_24_21_groupi_n_1016 ,csa_tree_add_24_21_groupi_n_1028);
  or csa_tree_add_24_21_groupi_g6315(csa_tree_add_24_21_groupi_n_1229 ,csa_tree_add_24_21_groupi_n_929 ,csa_tree_add_24_21_groupi_n_1090);
  or csa_tree_add_24_21_groupi_g6316(csa_tree_add_24_21_groupi_n_1228 ,csa_tree_add_24_21_groupi_n_1014 ,csa_tree_add_24_21_groupi_n_1084);
  or csa_tree_add_24_21_groupi_g6317(csa_tree_add_24_21_groupi_n_1227 ,csa_tree_add_24_21_groupi_n_1013 ,csa_tree_add_24_21_groupi_n_1083);
  or csa_tree_add_24_21_groupi_g6318(csa_tree_add_24_21_groupi_n_1226 ,csa_tree_add_24_21_groupi_n_984 ,csa_tree_add_24_21_groupi_n_1114);
  and csa_tree_add_24_21_groupi_g6319(csa_tree_add_24_21_groupi_n_1225 ,csa_tree_add_24_21_groupi_n_984 ,csa_tree_add_24_21_groupi_n_1114);
  nor csa_tree_add_24_21_groupi_g6320(csa_tree_add_24_21_groupi_n_1224 ,csa_tree_add_24_21_groupi_n_1081 ,csa_tree_add_24_21_groupi_n_910);
  or csa_tree_add_24_21_groupi_g6321(csa_tree_add_24_21_groupi_n_1223 ,csa_tree_add_24_21_groupi_n_1011 ,csa_tree_add_24_21_groupi_n_1075);
  or csa_tree_add_24_21_groupi_g6322(csa_tree_add_24_21_groupi_n_1222 ,csa_tree_add_24_21_groupi_n_895 ,csa_tree_add_24_21_groupi_n_1033);
  or csa_tree_add_24_21_groupi_g6323(csa_tree_add_24_21_groupi_n_1221 ,csa_tree_add_24_21_groupi_n_912 ,csa_tree_add_24_21_groupi_n_1073);
  or csa_tree_add_24_21_groupi_g6324(csa_tree_add_24_21_groupi_n_1220 ,csa_tree_add_24_21_groupi_n_1068 ,csa_tree_add_24_21_groupi_n_882);
  or csa_tree_add_24_21_groupi_g6325(csa_tree_add_24_21_groupi_n_1219 ,csa_tree_add_24_21_groupi_n_1010 ,csa_tree_add_24_21_groupi_n_1105);
  or csa_tree_add_24_21_groupi_g6326(csa_tree_add_24_21_groupi_n_1218 ,csa_tree_add_24_21_groupi_n_1009 ,csa_tree_add_24_21_groupi_n_1106);
  and csa_tree_add_24_21_groupi_g6327(csa_tree_add_24_21_groupi_n_1217 ,csa_tree_add_24_21_groupi_n_1068 ,csa_tree_add_24_21_groupi_n_882);
  or csa_tree_add_24_21_groupi_g6328(csa_tree_add_24_21_groupi_n_1216 ,csa_tree_add_24_21_groupi_n_1116 ,csa_tree_add_24_21_groupi_n_1122);
  nor csa_tree_add_24_21_groupi_g6329(csa_tree_add_24_21_groupi_n_1215 ,csa_tree_add_24_21_groupi_n_1115 ,csa_tree_add_24_21_groupi_n_1123);
  or csa_tree_add_24_21_groupi_g6330(csa_tree_add_24_21_groupi_n_1214 ,csa_tree_add_24_21_groupi_n_1008 ,csa_tree_add_24_21_groupi_n_1072);
  or csa_tree_add_24_21_groupi_g6331(csa_tree_add_24_21_groupi_n_1213 ,csa_tree_add_24_21_groupi_n_926 ,csa_tree_add_24_21_groupi_n_1094);
  or csa_tree_add_24_21_groupi_g6332(csa_tree_add_24_21_groupi_n_1212 ,csa_tree_add_24_21_groupi_n_899 ,csa_tree_add_24_21_groupi_n_1022);
  or csa_tree_add_24_21_groupi_g6333(csa_tree_add_24_21_groupi_n_1211 ,csa_tree_add_24_21_groupi_n_1003 ,csa_tree_add_24_21_groupi_n_1055);
  or csa_tree_add_24_21_groupi_g6334(csa_tree_add_24_21_groupi_n_1210 ,csa_tree_add_24_21_groupi_n_1111 ,csa_tree_add_24_21_groupi_n_901);
  or csa_tree_add_24_21_groupi_g6335(csa_tree_add_24_21_groupi_n_1209 ,csa_tree_add_24_21_groupi_n_1065 ,csa_tree_add_24_21_groupi_n_934);
  and csa_tree_add_24_21_groupi_g6336(csa_tree_add_24_21_groupi_n_1208 ,csa_tree_add_24_21_groupi_n_1065 ,csa_tree_add_24_21_groupi_n_934);
  or csa_tree_add_24_21_groupi_g6337(csa_tree_add_24_21_groupi_n_1207 ,csa_tree_add_24_21_groupi_n_1000 ,csa_tree_add_24_21_groupi_n_1051);
  or csa_tree_add_24_21_groupi_g6338(csa_tree_add_24_21_groupi_n_1206 ,csa_tree_add_24_21_groupi_n_1015 ,csa_tree_add_24_21_groupi_n_1047);
  or csa_tree_add_24_21_groupi_g6339(csa_tree_add_24_21_groupi_n_1205 ,csa_tree_add_24_21_groupi_n_913 ,csa_tree_add_24_21_groupi_n_1030);
  or csa_tree_add_24_21_groupi_g6340(csa_tree_add_24_21_groupi_n_1204 ,csa_tree_add_24_21_groupi_n_927 ,csa_tree_add_24_21_groupi_n_1044);
  and csa_tree_add_24_21_groupi_g6341(csa_tree_add_24_21_groupi_n_1203 ,csa_tree_add_24_21_groupi_n_1067 ,csa_tree_add_24_21_groupi_n_975);
  or csa_tree_add_24_21_groupi_g6342(csa_tree_add_24_21_groupi_n_1202 ,csa_tree_add_24_21_groupi_n_930 ,csa_tree_add_24_21_groupi_n_1041);
  or csa_tree_add_24_21_groupi_g6343(csa_tree_add_24_21_groupi_n_1201 ,csa_tree_add_24_21_groupi_n_1067 ,csa_tree_add_24_21_groupi_n_975);
  or csa_tree_add_24_21_groupi_g6344(csa_tree_add_24_21_groupi_n_1200 ,csa_tree_add_24_21_groupi_n_1070 ,csa_tree_add_24_21_groupi_n_996);
  or csa_tree_add_24_21_groupi_g6345(csa_tree_add_24_21_groupi_n_1199 ,csa_tree_add_24_21_groupi_n_915 ,csa_tree_add_24_21_groupi_n_1101);
  or csa_tree_add_24_21_groupi_g6346(csa_tree_add_24_21_groupi_n_1198 ,csa_tree_add_24_21_groupi_n_1017 ,csa_tree_add_24_21_groupi_n_1036);
  and csa_tree_add_24_21_groupi_g6347(csa_tree_add_24_21_groupi_n_1197 ,csa_tree_add_24_21_groupi_n_1069 ,csa_tree_add_24_21_groupi_n_973);
  or csa_tree_add_24_21_groupi_g6348(csa_tree_add_24_21_groupi_n_1196 ,csa_tree_add_24_21_groupi_n_1108 ,csa_tree_add_24_21_groupi_n_900);
  or csa_tree_add_24_21_groupi_g6349(csa_tree_add_24_21_groupi_n_1195 ,csa_tree_add_24_21_groupi_n_916 ,csa_tree_add_24_21_groupi_n_1034);
  and csa_tree_add_24_21_groupi_g6350(csa_tree_add_24_21_groupi_n_1254 ,csa_tree_add_24_21_groupi_n_373 ,csa_tree_add_24_21_groupi_n_1040);
  and csa_tree_add_24_21_groupi_g6351(csa_tree_add_24_21_groupi_n_1253 ,csa_tree_add_24_21_groupi_n_374 ,csa_tree_add_24_21_groupi_n_1042);
  and csa_tree_add_24_21_groupi_g6352(csa_tree_add_24_21_groupi_n_1252 ,csa_tree_add_24_21_groupi_n_841 ,csa_tree_add_24_21_groupi_n_1025);
  and csa_tree_add_24_21_groupi_g6353(csa_tree_add_24_21_groupi_n_1251 ,csa_tree_add_24_21_groupi_n_932 ,csa_tree_add_24_21_groupi_n_1096);
  and csa_tree_add_24_21_groupi_g6354(csa_tree_add_24_21_groupi_n_1250 ,csa_tree_add_24_21_groupi_n_838 ,csa_tree_add_24_21_groupi_n_1049);
  and csa_tree_add_24_21_groupi_g6355(csa_tree_add_24_21_groupi_n_1248 ,csa_tree_add_24_21_groupi_n_378 ,csa_tree_add_24_21_groupi_n_1039);
  or csa_tree_add_24_21_groupi_g6356(csa_tree_add_24_21_groupi_n_1247 ,csa_tree_add_24_21_groupi_n_383 ,csa_tree_add_24_21_groupi_n_1052);
  and csa_tree_add_24_21_groupi_g6357(csa_tree_add_24_21_groupi_n_1245 ,csa_tree_add_24_21_groupi_n_835 ,csa_tree_add_24_21_groupi_n_1098);
  and csa_tree_add_24_21_groupi_g6358(csa_tree_add_24_21_groupi_n_1244 ,csa_tree_add_24_21_groupi_n_836 ,csa_tree_add_24_21_groupi_n_1058);
  and csa_tree_add_24_21_groupi_g6359(csa_tree_add_24_21_groupi_n_1243 ,csa_tree_add_24_21_groupi_n_832 ,csa_tree_add_24_21_groupi_n_1071);
  and csa_tree_add_24_21_groupi_g6360(csa_tree_add_24_21_groupi_n_1241 ,csa_tree_add_24_21_groupi_n_379 ,csa_tree_add_24_21_groupi_n_1074);
  xnor csa_tree_add_24_21_groupi_g6361(csa_tree_add_24_21_groupi_n_1240 ,csa_tree_add_24_21_groupi_n_1020 ,in3[19]);
  and csa_tree_add_24_21_groupi_g6362(csa_tree_add_24_21_groupi_n_1239 ,csa_tree_add_24_21_groupi_n_840 ,csa_tree_add_24_21_groupi_n_1063);
  not csa_tree_add_24_21_groupi_g6363(csa_tree_add_24_21_groupi_n_1193 ,csa_tree_add_24_21_groupi_n_1192);
  not csa_tree_add_24_21_groupi_g6364(csa_tree_add_24_21_groupi_n_1190 ,csa_tree_add_24_21_groupi_n_1189);
  not csa_tree_add_24_21_groupi_g6365(csa_tree_add_24_21_groupi_n_1187 ,csa_tree_add_24_21_groupi_n_1188);
  not csa_tree_add_24_21_groupi_g6366(csa_tree_add_24_21_groupi_n_1184 ,csa_tree_add_24_21_groupi_n_1185);
  not csa_tree_add_24_21_groupi_g6367(csa_tree_add_24_21_groupi_n_1182 ,csa_tree_add_24_21_groupi_n_1183);
  not csa_tree_add_24_21_groupi_g6368(csa_tree_add_24_21_groupi_n_1180 ,csa_tree_add_24_21_groupi_n_1181);
  not csa_tree_add_24_21_groupi_g6369(csa_tree_add_24_21_groupi_n_1178 ,csa_tree_add_24_21_groupi_n_1179);
  not csa_tree_add_24_21_groupi_g6370(csa_tree_add_24_21_groupi_n_1176 ,csa_tree_add_24_21_groupi_n_1177);
  not csa_tree_add_24_21_groupi_g6371(csa_tree_add_24_21_groupi_n_1175 ,csa_tree_add_24_21_groupi_n_1174);
  not csa_tree_add_24_21_groupi_g6372(csa_tree_add_24_21_groupi_n_1172 ,csa_tree_add_24_21_groupi_n_1173);
  not csa_tree_add_24_21_groupi_g6373(csa_tree_add_24_21_groupi_n_1170 ,csa_tree_add_24_21_groupi_n_1171);
  not csa_tree_add_24_21_groupi_g6374(csa_tree_add_24_21_groupi_n_1168 ,csa_tree_add_24_21_groupi_n_1169);
  not csa_tree_add_24_21_groupi_g6375(csa_tree_add_24_21_groupi_n_1166 ,csa_tree_add_24_21_groupi_n_1167);
  not csa_tree_add_24_21_groupi_g6376(csa_tree_add_24_21_groupi_n_1164 ,csa_tree_add_24_21_groupi_n_1165);
  xnor csa_tree_add_24_21_groupi_g6377(csa_tree_add_24_21_groupi_n_1163 ,csa_tree_add_24_21_groupi_n_858 ,csa_tree_add_24_21_groupi_n_869);
  xnor csa_tree_add_24_21_groupi_g6378(csa_tree_add_24_21_groupi_n_1162 ,csa_tree_add_24_21_groupi_n_884 ,csa_tree_add_24_21_groupi_n_886);
  xnor csa_tree_add_24_21_groupi_g6379(csa_tree_add_24_21_groupi_n_1161 ,csa_tree_add_24_21_groupi_n_989 ,csa_tree_add_24_21_groupi_n_941);
  xnor csa_tree_add_24_21_groupi_g6380(csa_tree_add_24_21_groupi_n_1160 ,csa_tree_add_24_21_groupi_n_873 ,csa_tree_add_24_21_groupi_n_913);
  xnor csa_tree_add_24_21_groupi_g6381(csa_tree_add_24_21_groupi_n_1159 ,csa_tree_add_24_21_groupi_n_878 ,csa_tree_add_24_21_groupi_n_857);
  xor csa_tree_add_24_21_groupi_g6382(csa_tree_add_24_21_groupi_n_1158 ,csa_tree_add_24_21_groupi_n_1016 ,in3[20]);
  xnor csa_tree_add_24_21_groupi_g6383(csa_tree_add_24_21_groupi_n_1157 ,csa_tree_add_24_21_groupi_n_860 ,in3[24]);
  xnor csa_tree_add_24_21_groupi_g6384(csa_tree_add_24_21_groupi_n_1156 ,csa_tree_add_24_21_groupi_n_861 ,csa_tree_add_24_21_groupi_n_994);
  xnor csa_tree_add_24_21_groupi_g6385(csa_tree_add_24_21_groupi_n_1155 ,csa_tree_add_24_21_groupi_n_1011 ,csa_tree_add_24_21_groupi_n_979);
  xnor csa_tree_add_24_21_groupi_g6386(csa_tree_add_24_21_groupi_n_1154 ,csa_tree_add_24_21_groupi_n_961 ,csa_tree_add_24_21_groupi_n_955);
  xnor csa_tree_add_24_21_groupi_g6387(csa_tree_add_24_21_groupi_n_1153 ,csa_tree_add_24_21_groupi_n_945 ,in3[28]);
  xnor csa_tree_add_24_21_groupi_g6388(csa_tree_add_24_21_groupi_n_1152 ,csa_tree_add_24_21_groupi_n_947 ,csa_tree_add_24_21_groupi_n_943);
  xnor csa_tree_add_24_21_groupi_g6389(csa_tree_add_24_21_groupi_n_1151 ,csa_tree_add_24_21_groupi_n_959 ,in3[26]);
  xnor csa_tree_add_24_21_groupi_g6390(csa_tree_add_24_21_groupi_n_1150 ,csa_tree_add_24_21_groupi_n_975 ,csa_tree_add_24_21_groupi_n_911);
  xnor csa_tree_add_24_21_groupi_g6391(csa_tree_add_24_21_groupi_n_1149 ,csa_tree_add_24_21_groupi_n_759 ,csa_tree_add_24_21_groupi_n_922);
  xnor csa_tree_add_24_21_groupi_g6392(csa_tree_add_24_21_groupi_n_1148 ,csa_tree_add_24_21_groupi_n_916 ,csa_tree_add_24_21_groupi_n_872);
  xnor csa_tree_add_24_21_groupi_g6393(csa_tree_add_24_21_groupi_n_1147 ,csa_tree_add_24_21_groupi_n_973 ,csa_tree_add_24_21_groupi_n_919);
  xnor csa_tree_add_24_21_groupi_g6394(csa_tree_add_24_21_groupi_n_1146 ,csa_tree_add_24_21_groupi_n_910 ,in3[13]);
  xnor csa_tree_add_24_21_groupi_g6395(csa_tree_add_24_21_groupi_n_1145 ,csa_tree_add_24_21_groupi_n_855 ,csa_tree_add_24_21_groupi_n_930);
  xnor csa_tree_add_24_21_groupi_g6396(csa_tree_add_24_21_groupi_n_1144 ,csa_tree_add_24_21_groupi_n_993 ,csa_tree_add_24_21_groupi_n_1013);
  xnor csa_tree_add_24_21_groupi_g6397(csa_tree_add_24_21_groupi_n_1143 ,csa_tree_add_24_21_groupi_n_927 ,csa_tree_add_24_21_groupi_n_853);
  xnor csa_tree_add_24_21_groupi_g6398(csa_tree_add_24_21_groupi_n_1142 ,csa_tree_add_24_21_groupi_n_938 ,csa_tree_add_24_21_groupi_n_874);
  xnor csa_tree_add_24_21_groupi_g6399(csa_tree_add_24_21_groupi_n_1141 ,csa_tree_add_24_21_groupi_n_956 ,csa_tree_add_24_21_groupi_n_957);
  xnor csa_tree_add_24_21_groupi_g6400(csa_tree_add_24_21_groupi_n_1140 ,csa_tree_add_24_21_groupi_n_1009 ,csa_tree_add_24_21_groupi_n_966);
  xnor csa_tree_add_24_21_groupi_g6401(csa_tree_add_24_21_groupi_n_1139 ,csa_tree_add_24_21_groupi_n_965 ,csa_tree_add_24_21_groupi_n_995);
  xnor csa_tree_add_24_21_groupi_g6402(csa_tree_add_24_21_groupi_n_1138 ,csa_tree_add_24_21_groupi_n_871 ,csa_tree_add_24_21_groupi_n_903);
  xnor csa_tree_add_24_21_groupi_g6403(csa_tree_add_24_21_groupi_n_1137 ,csa_tree_add_24_21_groupi_n_968 ,csa_tree_add_24_21_groupi_n_852);
  xnor csa_tree_add_24_21_groupi_g6404(csa_tree_add_24_21_groupi_n_1136 ,csa_tree_add_24_21_groupi_n_879 ,csa_tree_add_24_21_groupi_n_868);
  xnor csa_tree_add_24_21_groupi_g6405(csa_tree_add_24_21_groupi_n_1135 ,csa_tree_add_24_21_groupi_n_972 ,csa_tree_add_24_21_groupi_n_974);
  xnor csa_tree_add_24_21_groupi_g6406(csa_tree_add_24_21_groupi_n_1134 ,csa_tree_add_24_21_groupi_n_998 ,csa_tree_add_24_21_groupi_n_876);
  xnor csa_tree_add_24_21_groupi_g6407(csa_tree_add_24_21_groupi_n_1133 ,csa_tree_add_24_21_groupi_n_926 ,csa_tree_add_24_21_groupi_n_888);
  xnor csa_tree_add_24_21_groupi_g6408(csa_tree_add_24_21_groupi_n_1132 ,csa_tree_add_24_21_groupi_n_990 ,csa_tree_add_24_21_groupi_n_991);
  xnor csa_tree_add_24_21_groupi_g6409(csa_tree_add_24_21_groupi_n_1131 ,csa_tree_add_24_21_groupi_n_887 ,csa_tree_add_24_21_groupi_n_892);
  xnor csa_tree_add_24_21_groupi_g6410(csa_tree_add_24_21_groupi_n_1130 ,csa_tree_add_24_21_groupi_n_881 ,csa_tree_add_24_21_groupi_n_971);
  xnor csa_tree_add_24_21_groupi_g6411(csa_tree_add_24_21_groupi_n_1129 ,csa_tree_add_24_21_groupi_n_863 ,csa_tree_add_24_21_groupi_n_880);
  xnor csa_tree_add_24_21_groupi_g6412(csa_tree_add_24_21_groupi_n_1128 ,csa_tree_add_24_21_groupi_n_999 ,csa_tree_add_24_21_groupi_n_986);
  xnor csa_tree_add_24_21_groupi_g6413(csa_tree_add_24_21_groupi_n_1127 ,csa_tree_add_24_21_groupi_n_1003 ,in3[22]);
  xnor csa_tree_add_24_21_groupi_g6414(csa_tree_add_24_21_groupi_n_1126 ,csa_tree_add_24_21_groupi_n_987 ,csa_tree_add_24_21_groupi_n_891);
  xnor csa_tree_add_24_21_groupi_g6415(csa_tree_add_24_21_groupi_n_1125 ,csa_tree_add_24_21_groupi_n_962 ,csa_tree_add_24_21_groupi_n_981);
  xnor csa_tree_add_24_21_groupi_g6416(csa_tree_add_24_21_groupi_n_1124 ,csa_tree_add_24_21_groupi_n_949 ,csa_tree_add_24_21_groupi_n_950);
  xnor csa_tree_add_24_21_groupi_g6417(csa_tree_add_24_21_groupi_n_1194 ,csa_tree_add_24_21_groupi_n_896 ,csa_tree_add_24_21_groupi_n_847);
  xnor csa_tree_add_24_21_groupi_g6418(csa_tree_add_24_21_groupi_n_1192 ,csa_tree_add_24_21_groupi_n_923 ,csa_tree_add_24_21_groupi_n_848);
  xnor csa_tree_add_24_21_groupi_g6419(csa_tree_add_24_21_groupi_n_1191 ,csa_tree_add_24_21_groupi_n_898 ,csa_tree_add_24_21_groupi_n_389);
  xnor csa_tree_add_24_21_groupi_g6420(csa_tree_add_24_21_groupi_n_1189 ,csa_tree_add_24_21_groupi_n_920 ,in3[15]);
  xnor csa_tree_add_24_21_groupi_g6421(csa_tree_add_24_21_groupi_n_1188 ,csa_tree_add_24_21_groupi_n_1018 ,csa_tree_add_24_21_groupi_n_1001);
  xnor csa_tree_add_24_21_groupi_g6422(csa_tree_add_24_21_groupi_n_1186 ,csa_tree_add_24_21_groupi_n_1006 ,in3[18]);
  xnor csa_tree_add_24_21_groupi_g6423(csa_tree_add_24_21_groupi_n_1185 ,csa_tree_add_24_21_groupi_n_914 ,csa_tree_add_24_21_groupi_n_846);
  xnor csa_tree_add_24_21_groupi_g6424(csa_tree_add_24_21_groupi_n_1183 ,csa_tree_add_24_21_groupi_n_906 ,csa_tree_add_24_21_groupi_n_845);
  xnor csa_tree_add_24_21_groupi_g6425(csa_tree_add_24_21_groupi_n_1181 ,csa_tree_add_24_21_groupi_n_907 ,csa_tree_add_24_21_groupi_n_849);
  xnor csa_tree_add_24_21_groupi_g6426(csa_tree_add_24_21_groupi_n_1179 ,csa_tree_add_24_21_groupi_n_1004 ,csa_tree_add_24_21_groupi_n_850);
  xnor csa_tree_add_24_21_groupi_g6427(csa_tree_add_24_21_groupi_n_1177 ,csa_tree_add_24_21_groupi_n_893 ,csa_tree_add_24_21_groupi_n_391);
  xnor csa_tree_add_24_21_groupi_g6428(csa_tree_add_24_21_groupi_n_1174 ,csa_tree_add_24_21_groupi_n_897 ,csa_tree_add_24_21_groupi_n_388);
  xnor csa_tree_add_24_21_groupi_g6429(csa_tree_add_24_21_groupi_n_1173 ,csa_tree_add_24_21_groupi_n_904 ,in3[17]);
  xnor csa_tree_add_24_21_groupi_g6430(csa_tree_add_24_21_groupi_n_1171 ,csa_tree_add_24_21_groupi_n_894 ,csa_tree_add_24_21_groupi_n_392);
  xnor csa_tree_add_24_21_groupi_g6431(csa_tree_add_24_21_groupi_n_1169 ,csa_tree_add_24_21_groupi_n_908 ,in3[14]);
  xnor csa_tree_add_24_21_groupi_g6432(csa_tree_add_24_21_groupi_n_1167 ,csa_tree_add_24_21_groupi_n_924 ,in3[16]);
  xnor csa_tree_add_24_21_groupi_g6433(csa_tree_add_24_21_groupi_n_1165 ,csa_tree_add_24_21_groupi_n_928 ,csa_tree_add_24_21_groupi_n_390);
  not csa_tree_add_24_21_groupi_g6434(csa_tree_add_24_21_groupi_n_1122 ,csa_tree_add_24_21_groupi_n_1123);
  not csa_tree_add_24_21_groupi_g6435(csa_tree_add_24_21_groupi_n_1121 ,csa_tree_add_24_21_groupi_n_1120);
  not csa_tree_add_24_21_groupi_g6436(csa_tree_add_24_21_groupi_n_1118 ,csa_tree_add_24_21_groupi_n_1117);
  not csa_tree_add_24_21_groupi_g6437(csa_tree_add_24_21_groupi_n_1116 ,csa_tree_add_24_21_groupi_n_1115);
  or csa_tree_add_24_21_groupi_g6438(csa_tree_add_24_21_groupi_n_1113 ,csa_tree_add_24_21_groupi_n_963 ,csa_tree_add_24_21_groupi_n_872);
  or csa_tree_add_24_21_groupi_g6439(csa_tree_add_24_21_groupi_n_1112 ,in3[26] ,csa_tree_add_24_21_groupi_n_958);
  nor csa_tree_add_24_21_groupi_g6440(csa_tree_add_24_21_groupi_n_1111 ,csa_tree_add_24_21_groupi_n_349 ,csa_tree_add_24_21_groupi_n_860);
  nor csa_tree_add_24_21_groupi_g6441(csa_tree_add_24_21_groupi_n_1110 ,csa_tree_add_24_21_groupi_n_348 ,csa_tree_add_24_21_groupi_n_959);
  or csa_tree_add_24_21_groupi_g6442(csa_tree_add_24_21_groupi_n_1109 ,in3[24] ,csa_tree_add_24_21_groupi_n_859);
  nor csa_tree_add_24_21_groupi_g6443(csa_tree_add_24_21_groupi_n_1108 ,csa_tree_add_24_21_groupi_n_328 ,csa_tree_add_24_21_groupi_n_945);
  or csa_tree_add_24_21_groupi_g6444(csa_tree_add_24_21_groupi_n_1107 ,in3[28] ,csa_tree_add_24_21_groupi_n_944);
  and csa_tree_add_24_21_groupi_g6445(csa_tree_add_24_21_groupi_n_1106 ,csa_tree_add_24_21_groupi_n_969 ,csa_tree_add_24_21_groupi_n_966);
  and csa_tree_add_24_21_groupi_g6446(csa_tree_add_24_21_groupi_n_1105 ,csa_tree_add_24_21_groupi_n_852 ,csa_tree_add_24_21_groupi_n_968);
  or csa_tree_add_24_21_groupi_g6447(csa_tree_add_24_21_groupi_n_1104 ,csa_tree_add_24_21_groupi_n_981 ,csa_tree_add_24_21_groupi_n_962);
  or csa_tree_add_24_21_groupi_g6448(csa_tree_add_24_21_groupi_n_1103 ,csa_tree_add_24_21_groupi_n_969 ,csa_tree_add_24_21_groupi_n_966);
  or csa_tree_add_24_21_groupi_g6449(csa_tree_add_24_21_groupi_n_1102 ,csa_tree_add_24_21_groupi_n_988 ,csa_tree_add_24_21_groupi_n_941);
  and csa_tree_add_24_21_groupi_g6450(csa_tree_add_24_21_groupi_n_1101 ,csa_tree_add_24_21_groupi_n_880 ,csa_tree_add_24_21_groupi_n_863);
  or csa_tree_add_24_21_groupi_g6451(csa_tree_add_24_21_groupi_n_1100 ,csa_tree_add_24_21_groupi_n_877 ,csa_tree_add_24_21_groupi_n_857);
  or csa_tree_add_24_21_groupi_g6452(csa_tree_add_24_21_groupi_n_1099 ,csa_tree_add_24_21_groupi_n_875 ,csa_tree_add_24_21_groupi_n_997);
  or csa_tree_add_24_21_groupi_g6453(csa_tree_add_24_21_groupi_n_1098 ,csa_tree_add_24_21_groupi_n_834 ,csa_tree_add_24_21_groupi_n_906);
  nor csa_tree_add_24_21_groupi_g6454(csa_tree_add_24_21_groupi_n_1097 ,csa_tree_add_24_21_groupi_n_878 ,csa_tree_add_24_21_groupi_n_856);
  or csa_tree_add_24_21_groupi_g6455(csa_tree_add_24_21_groupi_n_1096 ,csa_tree_add_24_21_groupi_n_931 ,csa_tree_add_24_21_groupi_n_922);
  and csa_tree_add_24_21_groupi_g6456(csa_tree_add_24_21_groupi_n_1095 ,csa_tree_add_24_21_groupi_n_868 ,csa_tree_add_24_21_groupi_n_879);
  and csa_tree_add_24_21_groupi_g6457(csa_tree_add_24_21_groupi_n_1094 ,csa_tree_add_24_21_groupi_n_888 ,csa_tree_add_24_21_groupi_n_890);
  or csa_tree_add_24_21_groupi_g6458(csa_tree_add_24_21_groupi_n_1093 ,csa_tree_add_24_21_groupi_n_948 ,csa_tree_add_24_21_groupi_n_873);
  or csa_tree_add_24_21_groupi_g6459(csa_tree_add_24_21_groupi_n_1092 ,csa_tree_add_24_21_groupi_n_874 ,csa_tree_add_24_21_groupi_n_938);
  and csa_tree_add_24_21_groupi_g6460(csa_tree_add_24_21_groupi_n_1091 ,csa_tree_add_24_21_groupi_n_981 ,csa_tree_add_24_21_groupi_n_962);
  and csa_tree_add_24_21_groupi_g6461(csa_tree_add_24_21_groupi_n_1090 ,csa_tree_add_24_21_groupi_n_950 ,csa_tree_add_24_21_groupi_n_949);
  or csa_tree_add_24_21_groupi_g6462(csa_tree_add_24_21_groupi_n_1089 ,csa_tree_add_24_21_groupi_n_950 ,csa_tree_add_24_21_groupi_n_949);
  or csa_tree_add_24_21_groupi_g6463(csa_tree_add_24_21_groupi_n_1088 ,csa_tree_add_24_21_groupi_n_951 ,csa_tree_add_24_21_groupi_n_993);
  nor csa_tree_add_24_21_groupi_g6464(csa_tree_add_24_21_groupi_n_1087 ,csa_tree_add_24_21_groupi_n_989 ,csa_tree_add_24_21_groupi_n_940);
  or csa_tree_add_24_21_groupi_g6465(csa_tree_add_24_21_groupi_n_1086 ,csa_tree_add_24_21_groupi_n_995 ,csa_tree_add_24_21_groupi_n_965);
  or csa_tree_add_24_21_groupi_g6466(csa_tree_add_24_21_groupi_n_1085 ,csa_tree_add_24_21_groupi_n_991 ,csa_tree_add_24_21_groupi_n_990);
  and csa_tree_add_24_21_groupi_g6467(csa_tree_add_24_21_groupi_n_1084 ,csa_tree_add_24_21_groupi_n_991 ,csa_tree_add_24_21_groupi_n_990);
  nor csa_tree_add_24_21_groupi_g6468(csa_tree_add_24_21_groupi_n_1083 ,csa_tree_add_24_21_groupi_n_952 ,csa_tree_add_24_21_groupi_n_992);
  and csa_tree_add_24_21_groupi_g6469(csa_tree_add_24_21_groupi_n_1082 ,in3[13] ,csa_tree_add_24_21_groupi_n_980);
  nor csa_tree_add_24_21_groupi_g6470(csa_tree_add_24_21_groupi_n_1081 ,in3[13] ,csa_tree_add_24_21_groupi_n_980);
  or csa_tree_add_24_21_groupi_g6471(csa_tree_add_24_21_groupi_n_1080 ,csa_tree_add_24_21_groupi_n_978 ,csa_tree_add_24_21_groupi_n_977);
  or csa_tree_add_24_21_groupi_g6472(csa_tree_add_24_21_groupi_n_1079 ,csa_tree_add_24_21_groupi_n_862 ,csa_tree_add_24_21_groupi_n_994);
  or csa_tree_add_24_21_groupi_g6473(csa_tree_add_24_21_groupi_n_1078 ,csa_tree_add_24_21_groupi_n_974 ,csa_tree_add_24_21_groupi_n_972);
  and csa_tree_add_24_21_groupi_g6474(csa_tree_add_24_21_groupi_n_1077 ,csa_tree_add_24_21_groupi_n_974 ,csa_tree_add_24_21_groupi_n_972);
  or csa_tree_add_24_21_groupi_g6475(csa_tree_add_24_21_groupi_n_1076 ,csa_tree_add_24_21_groupi_n_971 ,csa_tree_add_24_21_groupi_n_881);
  nor csa_tree_add_24_21_groupi_g6476(csa_tree_add_24_21_groupi_n_1075 ,csa_tree_add_24_21_groupi_n_979 ,csa_tree_add_24_21_groupi_n_976);
  or csa_tree_add_24_21_groupi_g6477(csa_tree_add_24_21_groupi_n_1074 ,csa_tree_add_24_21_groupi_n_385 ,csa_tree_add_24_21_groupi_n_893);
  and csa_tree_add_24_21_groupi_g6478(csa_tree_add_24_21_groupi_n_1073 ,csa_tree_add_24_21_groupi_n_971 ,csa_tree_add_24_21_groupi_n_881);
  and csa_tree_add_24_21_groupi_g6479(csa_tree_add_24_21_groupi_n_1072 ,csa_tree_add_24_21_groupi_n_891 ,csa_tree_add_24_21_groupi_n_987);
  or csa_tree_add_24_21_groupi_g6480(csa_tree_add_24_21_groupi_n_1071 ,csa_tree_add_24_21_groupi_n_833 ,csa_tree_add_24_21_groupi_n_914);
  and csa_tree_add_24_21_groupi_g6481(csa_tree_add_24_21_groupi_n_1123 ,csa_tree_add_24_21_groupi_n_1018 ,csa_tree_add_24_21_groupi_n_1002);
  and csa_tree_add_24_21_groupi_g6482(csa_tree_add_24_21_groupi_n_1120 ,in3[16] ,csa_tree_add_24_21_groupi_n_925);
  or csa_tree_add_24_21_groupi_g6483(csa_tree_add_24_21_groupi_n_1119 ,csa_tree_add_24_21_groupi_n_340 ,csa_tree_add_24_21_groupi_n_904);
  and csa_tree_add_24_21_groupi_g6484(csa_tree_add_24_21_groupi_n_1117 ,in3[15] ,csa_tree_add_24_21_groupi_n_921);
  and csa_tree_add_24_21_groupi_g6485(csa_tree_add_24_21_groupi_n_1115 ,in3[14] ,csa_tree_add_24_21_groupi_n_909);
  and csa_tree_add_24_21_groupi_g6486(csa_tree_add_24_21_groupi_n_1114 ,csa_tree_add_24_21_groupi_n_363 ,csa_tree_add_24_21_groupi_n_1020);
  or csa_tree_add_24_21_groupi_g6487(csa_tree_add_24_21_groupi_n_1064 ,csa_tree_add_24_21_groupi_n_869 ,csa_tree_add_24_21_groupi_n_858);
  or csa_tree_add_24_21_groupi_g6488(csa_tree_add_24_21_groupi_n_1063 ,csa_tree_add_24_21_groupi_n_839 ,csa_tree_add_24_21_groupi_n_1004);
  and csa_tree_add_24_21_groupi_g6489(csa_tree_add_24_21_groupi_n_1062 ,csa_tree_add_24_21_groupi_n_939 ,csa_tree_add_24_21_groupi_n_986);
  or csa_tree_add_24_21_groupi_g6490(csa_tree_add_24_21_groupi_n_1061 ,csa_tree_add_24_21_groupi_n_960 ,csa_tree_add_24_21_groupi_n_955);
  or csa_tree_add_24_21_groupi_g6491(csa_tree_add_24_21_groupi_n_1060 ,in3[22] ,csa_tree_add_24_21_groupi_n_964);
  or csa_tree_add_24_21_groupi_g6492(csa_tree_add_24_21_groupi_n_1059 ,csa_tree_add_24_21_groupi_n_957 ,csa_tree_add_24_21_groupi_n_956);
  or csa_tree_add_24_21_groupi_g6493(csa_tree_add_24_21_groupi_n_1058 ,csa_tree_add_24_21_groupi_n_806 ,csa_tree_add_24_21_groupi_n_896);
  and csa_tree_add_24_21_groupi_g6494(csa_tree_add_24_21_groupi_n_1057 ,csa_tree_add_24_21_groupi_n_957 ,csa_tree_add_24_21_groupi_n_956);
  or csa_tree_add_24_21_groupi_g6495(csa_tree_add_24_21_groupi_n_1056 ,csa_tree_add_24_21_groupi_n_946 ,csa_tree_add_24_21_groupi_n_943);
  and csa_tree_add_24_21_groupi_g6496(csa_tree_add_24_21_groupi_n_1055 ,in3[22] ,csa_tree_add_24_21_groupi_n_964);
  and csa_tree_add_24_21_groupi_g6497(csa_tree_add_24_21_groupi_n_1054 ,csa_tree_add_24_21_groupi_n_892 ,csa_tree_add_24_21_groupi_n_887);
  or csa_tree_add_24_21_groupi_g6498(csa_tree_add_24_21_groupi_n_1053 ,csa_tree_add_24_21_groupi_n_870 ,csa_tree_add_24_21_groupi_n_937);
  and csa_tree_add_24_21_groupi_g6499(csa_tree_add_24_21_groupi_n_1052 ,csa_tree_add_24_21_groupi_n_368 ,csa_tree_add_24_21_groupi_n_928);
  nor csa_tree_add_24_21_groupi_g6500(csa_tree_add_24_21_groupi_n_1051 ,csa_tree_add_24_21_groupi_n_947 ,csa_tree_add_24_21_groupi_n_942);
  or csa_tree_add_24_21_groupi_g6501(csa_tree_add_24_21_groupi_n_1050 ,csa_tree_add_24_21_groupi_n_852 ,csa_tree_add_24_21_groupi_n_968);
  or csa_tree_add_24_21_groupi_g6502(csa_tree_add_24_21_groupi_n_1049 ,csa_tree_add_24_21_groupi_n_842 ,csa_tree_add_24_21_groupi_n_923);
  or csa_tree_add_24_21_groupi_g6503(csa_tree_add_24_21_groupi_n_1048 ,csa_tree_add_24_21_groupi_n_853 ,csa_tree_add_24_21_groupi_n_970);
  nor csa_tree_add_24_21_groupi_g6504(csa_tree_add_24_21_groupi_n_1047 ,csa_tree_add_24_21_groupi_n_961 ,csa_tree_add_24_21_groupi_n_954);
  or csa_tree_add_24_21_groupi_g6505(csa_tree_add_24_21_groupi_n_1046 ,csa_tree_add_24_21_groupi_n_854 ,csa_tree_add_24_21_groupi_n_855);
  nor csa_tree_add_24_21_groupi_g6506(csa_tree_add_24_21_groupi_n_1045 ,csa_tree_add_24_21_groupi_n_871 ,csa_tree_add_24_21_groupi_n_936);
  and csa_tree_add_24_21_groupi_g6507(csa_tree_add_24_21_groupi_n_1044 ,csa_tree_add_24_21_groupi_n_853 ,csa_tree_add_24_21_groupi_n_970);
  or csa_tree_add_24_21_groupi_g6508(csa_tree_add_24_21_groupi_n_1043 ,csa_tree_add_24_21_groupi_n_891 ,csa_tree_add_24_21_groupi_n_987);
  or csa_tree_add_24_21_groupi_g6509(csa_tree_add_24_21_groupi_n_1042 ,csa_tree_add_24_21_groupi_n_370 ,csa_tree_add_24_21_groupi_n_897);
  and csa_tree_add_24_21_groupi_g6510(csa_tree_add_24_21_groupi_n_1041 ,csa_tree_add_24_21_groupi_n_854 ,csa_tree_add_24_21_groupi_n_855);
  or csa_tree_add_24_21_groupi_g6511(csa_tree_add_24_21_groupi_n_1040 ,csa_tree_add_24_21_groupi_n_377 ,csa_tree_add_24_21_groupi_n_894);
  or csa_tree_add_24_21_groupi_g6512(csa_tree_add_24_21_groupi_n_1039 ,csa_tree_add_24_21_groupi_n_366 ,csa_tree_add_24_21_groupi_n_898);
  and csa_tree_add_24_21_groupi_g6513(csa_tree_add_24_21_groupi_n_1038 ,csa_tree_add_24_21_groupi_n_869 ,csa_tree_add_24_21_groupi_n_858);
  or csa_tree_add_24_21_groupi_g6514(csa_tree_add_24_21_groupi_n_1037 ,csa_tree_add_24_21_groupi_n_880 ,csa_tree_add_24_21_groupi_n_863);
  and csa_tree_add_24_21_groupi_g6515(csa_tree_add_24_21_groupi_n_1036 ,csa_tree_add_24_21_groupi_n_862 ,csa_tree_add_24_21_groupi_n_994);
  or csa_tree_add_24_21_groupi_g6516(csa_tree_add_24_21_groupi_n_1035 ,csa_tree_add_24_21_groupi_n_892 ,csa_tree_add_24_21_groupi_n_887);
  and csa_tree_add_24_21_groupi_g6517(csa_tree_add_24_21_groupi_n_1034 ,csa_tree_add_24_21_groupi_n_963 ,csa_tree_add_24_21_groupi_n_872);
  and csa_tree_add_24_21_groupi_g6518(csa_tree_add_24_21_groupi_n_1033 ,csa_tree_add_24_21_groupi_n_995 ,csa_tree_add_24_21_groupi_n_965);
  and csa_tree_add_24_21_groupi_g6519(csa_tree_add_24_21_groupi_n_1032 ,csa_tree_add_24_21_groupi_n_874 ,csa_tree_add_24_21_groupi_n_938);
  nor csa_tree_add_24_21_groupi_g6520(csa_tree_add_24_21_groupi_n_1031 ,csa_tree_add_24_21_groupi_n_876 ,csa_tree_add_24_21_groupi_n_998);
  and csa_tree_add_24_21_groupi_g6521(csa_tree_add_24_21_groupi_n_1030 ,csa_tree_add_24_21_groupi_n_948 ,csa_tree_add_24_21_groupi_n_873);
  or csa_tree_add_24_21_groupi_g6522(csa_tree_add_24_21_groupi_n_1029 ,csa_tree_add_24_21_groupi_n_939 ,csa_tree_add_24_21_groupi_n_986);
  and csa_tree_add_24_21_groupi_g6523(csa_tree_add_24_21_groupi_n_1028 ,in3[20] ,csa_tree_add_24_21_groupi_n_889);
  or csa_tree_add_24_21_groupi_g6524(csa_tree_add_24_21_groupi_n_1027 ,in3[20] ,csa_tree_add_24_21_groupi_n_889);
  nor csa_tree_add_24_21_groupi_g6525(csa_tree_add_24_21_groupi_n_1026 ,csa_tree_add_24_21_groupi_n_868 ,csa_tree_add_24_21_groupi_n_879);
  or csa_tree_add_24_21_groupi_g6526(csa_tree_add_24_21_groupi_n_1025 ,csa_tree_add_24_21_groupi_n_837 ,csa_tree_add_24_21_groupi_n_907);
  or csa_tree_add_24_21_groupi_g6527(csa_tree_add_24_21_groupi_n_1024 ,csa_tree_add_24_21_groupi_n_883 ,csa_tree_add_24_21_groupi_n_886);
  or csa_tree_add_24_21_groupi_g6528(csa_tree_add_24_21_groupi_n_1023 ,csa_tree_add_24_21_groupi_n_888 ,csa_tree_add_24_21_groupi_n_890);
  nor csa_tree_add_24_21_groupi_g6529(csa_tree_add_24_21_groupi_n_1022 ,csa_tree_add_24_21_groupi_n_884 ,csa_tree_add_24_21_groupi_n_885);
  xnor csa_tree_add_24_21_groupi_g6530(csa_tree_add_24_21_groupi_n_1021 ,csa_tree_add_24_21_groupi_n_844 ,in3[30]);
  xnor csa_tree_add_24_21_groupi_g6531(csa_tree_add_24_21_groupi_n_1070 ,csa_tree_add_24_21_groupi_n_768 ,in3[3]);
  xnor csa_tree_add_24_21_groupi_g6532(csa_tree_add_24_21_groupi_n_1069 ,csa_tree_add_24_21_groupi_n_766 ,in3[9]);
  xnor csa_tree_add_24_21_groupi_g6533(csa_tree_add_24_21_groupi_n_1068 ,csa_tree_add_24_21_groupi_n_764 ,in3[5]);
  xnor csa_tree_add_24_21_groupi_g6534(csa_tree_add_24_21_groupi_n_1067 ,csa_tree_add_24_21_groupi_n_760 ,in3[7]);
  or csa_tree_add_24_21_groupi_g6535(csa_tree_add_24_21_groupi_n_1066 ,csa_tree_add_24_21_groupi_n_341 ,csa_tree_add_24_21_groupi_n_1007);
  xnor csa_tree_add_24_21_groupi_g6536(csa_tree_add_24_21_groupi_n_1065 ,csa_tree_add_24_21_groupi_n_762 ,in3[11]);
  not csa_tree_add_24_21_groupi_g6537(csa_tree_add_24_21_groupi_n_1007 ,csa_tree_add_24_21_groupi_n_1006);
  not csa_tree_add_24_21_groupi_g6538(csa_tree_add_24_21_groupi_n_1002 ,csa_tree_add_24_21_groupi_n_1001);
  not csa_tree_add_24_21_groupi_g6539(csa_tree_add_24_21_groupi_n_997 ,csa_tree_add_24_21_groupi_n_998);
  not csa_tree_add_24_21_groupi_g6540(csa_tree_add_24_21_groupi_n_992 ,csa_tree_add_24_21_groupi_n_993);
  not csa_tree_add_24_21_groupi_g6541(csa_tree_add_24_21_groupi_n_988 ,csa_tree_add_24_21_groupi_n_989);
  not csa_tree_add_24_21_groupi_g6542(csa_tree_add_24_21_groupi_n_982 ,csa_tree_add_24_21_groupi_n_983);
  not csa_tree_add_24_21_groupi_g6543(csa_tree_add_24_21_groupi_n_978 ,csa_tree_add_24_21_groupi_n_979);
  not csa_tree_add_24_21_groupi_g6544(csa_tree_add_24_21_groupi_n_976 ,csa_tree_add_24_21_groupi_n_977);
  not csa_tree_add_24_21_groupi_g6545(csa_tree_add_24_21_groupi_n_960 ,csa_tree_add_24_21_groupi_n_961);
  not csa_tree_add_24_21_groupi_g6546(csa_tree_add_24_21_groupi_n_958 ,csa_tree_add_24_21_groupi_n_959);
  not csa_tree_add_24_21_groupi_g6547(csa_tree_add_24_21_groupi_n_954 ,csa_tree_add_24_21_groupi_n_955);
  not csa_tree_add_24_21_groupi_g6548(csa_tree_add_24_21_groupi_n_951 ,csa_tree_add_24_21_groupi_n_952);
  not csa_tree_add_24_21_groupi_g6549(csa_tree_add_24_21_groupi_n_946 ,csa_tree_add_24_21_groupi_n_947);
  not csa_tree_add_24_21_groupi_g6550(csa_tree_add_24_21_groupi_n_944 ,csa_tree_add_24_21_groupi_n_945);
  not csa_tree_add_24_21_groupi_g6551(csa_tree_add_24_21_groupi_n_942 ,csa_tree_add_24_21_groupi_n_943);
  not csa_tree_add_24_21_groupi_g6552(csa_tree_add_24_21_groupi_n_940 ,csa_tree_add_24_21_groupi_n_941);
  not csa_tree_add_24_21_groupi_g6553(csa_tree_add_24_21_groupi_n_936 ,csa_tree_add_24_21_groupi_n_937);
  and csa_tree_add_24_21_groupi_g6554(csa_tree_add_24_21_groupi_n_933 ,in3[30] ,csa_tree_add_24_21_groupi_n_844);
  or csa_tree_add_24_21_groupi_g6555(csa_tree_add_24_21_groupi_n_932 ,csa_tree_add_24_21_groupi_n_257 ,csa_tree_add_24_21_groupi_n_758);
  nor csa_tree_add_24_21_groupi_g6556(csa_tree_add_24_21_groupi_n_931 ,csa_tree_add_24_21_groupi_n_320 ,csa_tree_add_24_21_groupi_n_759);
  and csa_tree_add_24_21_groupi_g6557(csa_tree_add_24_21_groupi_n_1020 ,csa_tree_add_24_21_groupi_n_640 ,csa_tree_add_24_21_groupi_n_744);
  and csa_tree_add_24_21_groupi_g6558(csa_tree_add_24_21_groupi_n_1019 ,csa_tree_add_24_21_groupi_n_650 ,csa_tree_add_24_21_groupi_n_813);
  or csa_tree_add_24_21_groupi_g6559(csa_tree_add_24_21_groupi_n_1018 ,csa_tree_add_24_21_groupi_n_679 ,csa_tree_add_24_21_groupi_n_829);
  and csa_tree_add_24_21_groupi_g6560(csa_tree_add_24_21_groupi_n_1017 ,csa_tree_add_24_21_groupi_n_627 ,csa_tree_add_24_21_groupi_n_701);
  and csa_tree_add_24_21_groupi_g6561(csa_tree_add_24_21_groupi_n_1016 ,csa_tree_add_24_21_groupi_n_671 ,csa_tree_add_24_21_groupi_n_818);
  and csa_tree_add_24_21_groupi_g6562(csa_tree_add_24_21_groupi_n_1015 ,csa_tree_add_24_21_groupi_n_617 ,csa_tree_add_24_21_groupi_n_733);
  and csa_tree_add_24_21_groupi_g6563(csa_tree_add_24_21_groupi_n_1014 ,csa_tree_add_24_21_groupi_n_559 ,csa_tree_add_24_21_groupi_n_746);
  and csa_tree_add_24_21_groupi_g6564(csa_tree_add_24_21_groupi_n_1013 ,csa_tree_add_24_21_groupi_n_565 ,csa_tree_add_24_21_groupi_n_810);
  and csa_tree_add_24_21_groupi_g6565(csa_tree_add_24_21_groupi_n_1012 ,csa_tree_add_24_21_groupi_n_572 ,csa_tree_add_24_21_groupi_n_719);
  or csa_tree_add_24_21_groupi_g6566(csa_tree_add_24_21_groupi_n_1011 ,csa_tree_add_24_21_groupi_n_375 ,csa_tree_add_24_21_groupi_n_689);
  and csa_tree_add_24_21_groupi_g6567(csa_tree_add_24_21_groupi_n_1010 ,csa_tree_add_24_21_groupi_n_624 ,csa_tree_add_24_21_groupi_n_736);
  and csa_tree_add_24_21_groupi_g6568(csa_tree_add_24_21_groupi_n_1009 ,csa_tree_add_24_21_groupi_n_634 ,csa_tree_add_24_21_groupi_n_738);
  and csa_tree_add_24_21_groupi_g6569(csa_tree_add_24_21_groupi_n_1008 ,csa_tree_add_24_21_groupi_n_663 ,csa_tree_add_24_21_groupi_n_700);
  or csa_tree_add_24_21_groupi_g6570(csa_tree_add_24_21_groupi_n_1006 ,csa_tree_add_24_21_groupi_n_375 ,csa_tree_add_24_21_groupi_n_789);
  and csa_tree_add_24_21_groupi_g6571(csa_tree_add_24_21_groupi_n_1005 ,csa_tree_add_24_21_groupi_n_626 ,csa_tree_add_24_21_groupi_n_778);
  and csa_tree_add_24_21_groupi_g6572(csa_tree_add_24_21_groupi_n_1004 ,csa_tree_add_24_21_groupi_n_569 ,csa_tree_add_24_21_groupi_n_727);
  and csa_tree_add_24_21_groupi_g6573(csa_tree_add_24_21_groupi_n_1003 ,csa_tree_add_24_21_groupi_n_649 ,csa_tree_add_24_21_groupi_n_739);
  and csa_tree_add_24_21_groupi_g6574(csa_tree_add_24_21_groupi_n_1001 ,csa_tree_add_24_21_groupi_n_629 ,csa_tree_add_24_21_groupi_n_720);
  and csa_tree_add_24_21_groupi_g6575(csa_tree_add_24_21_groupi_n_1000 ,csa_tree_add_24_21_groupi_n_567 ,csa_tree_add_24_21_groupi_n_724);
  and csa_tree_add_24_21_groupi_g6576(csa_tree_add_24_21_groupi_n_999 ,csa_tree_add_24_21_groupi_n_651 ,csa_tree_add_24_21_groupi_n_770);
  and csa_tree_add_24_21_groupi_g6577(csa_tree_add_24_21_groupi_n_998 ,csa_tree_add_24_21_groupi_n_655 ,csa_tree_add_24_21_groupi_n_777);
  and csa_tree_add_24_21_groupi_g6578(csa_tree_add_24_21_groupi_n_996 ,csa_tree_add_24_21_groupi_n_562 ,csa_tree_add_24_21_groupi_n_776);
  and csa_tree_add_24_21_groupi_g6579(csa_tree_add_24_21_groupi_n_995 ,csa_tree_add_24_21_groupi_n_654 ,csa_tree_add_24_21_groupi_n_817);
  and csa_tree_add_24_21_groupi_g6580(csa_tree_add_24_21_groupi_n_994 ,csa_tree_add_24_21_groupi_n_631 ,csa_tree_add_24_21_groupi_n_716);
  and csa_tree_add_24_21_groupi_g6581(csa_tree_add_24_21_groupi_n_993 ,csa_tree_add_24_21_groupi_n_643 ,csa_tree_add_24_21_groupi_n_750);
  and csa_tree_add_24_21_groupi_g6582(csa_tree_add_24_21_groupi_n_991 ,csa_tree_add_24_21_groupi_n_581 ,csa_tree_add_24_21_groupi_n_748);
  and csa_tree_add_24_21_groupi_g6583(csa_tree_add_24_21_groupi_n_990 ,csa_tree_add_24_21_groupi_n_642 ,csa_tree_add_24_21_groupi_n_747);
  or csa_tree_add_24_21_groupi_g6584(csa_tree_add_24_21_groupi_n_989 ,csa_tree_add_24_21_groupi_n_675 ,csa_tree_add_24_21_groupi_n_830);
  and csa_tree_add_24_21_groupi_g6585(csa_tree_add_24_21_groupi_n_987 ,csa_tree_add_24_21_groupi_n_571 ,csa_tree_add_24_21_groupi_n_702);
  and csa_tree_add_24_21_groupi_g6586(csa_tree_add_24_21_groupi_n_986 ,csa_tree_add_24_21_groupi_n_653 ,csa_tree_add_24_21_groupi_n_753);
  and csa_tree_add_24_21_groupi_g6587(csa_tree_add_24_21_groupi_n_985 ,csa_tree_add_24_21_groupi_n_646 ,csa_tree_add_24_21_groupi_n_732);
  and csa_tree_add_24_21_groupi_g6588(csa_tree_add_24_21_groupi_n_984 ,csa_tree_add_24_21_groupi_n_568 ,csa_tree_add_24_21_groupi_n_745);
  and csa_tree_add_24_21_groupi_g6589(csa_tree_add_24_21_groupi_n_983 ,csa_tree_add_24_21_groupi_n_641 ,csa_tree_add_24_21_groupi_n_809);
  and csa_tree_add_24_21_groupi_g6590(csa_tree_add_24_21_groupi_n_981 ,csa_tree_add_24_21_groupi_n_639 ,csa_tree_add_24_21_groupi_n_734);
  or csa_tree_add_24_21_groupi_g6591(csa_tree_add_24_21_groupi_n_980 ,csa_tree_add_24_21_groupi_n_676 ,csa_tree_add_24_21_groupi_n_694);
  or csa_tree_add_24_21_groupi_g6592(csa_tree_add_24_21_groupi_n_979 ,csa_tree_add_24_21_groupi_n_678 ,csa_tree_add_24_21_groupi_n_825);
  and csa_tree_add_24_21_groupi_g6593(csa_tree_add_24_21_groupi_n_977 ,csa_tree_add_24_21_groupi_n_556 ,csa_tree_add_24_21_groupi_n_743);
  and csa_tree_add_24_21_groupi_g6594(csa_tree_add_24_21_groupi_n_975 ,csa_tree_add_24_21_groupi_n_652 ,csa_tree_add_24_21_groupi_n_708);
  and csa_tree_add_24_21_groupi_g6595(csa_tree_add_24_21_groupi_n_974 ,csa_tree_add_24_21_groupi_n_580 ,csa_tree_add_24_21_groupi_n_797);
  and csa_tree_add_24_21_groupi_g6596(csa_tree_add_24_21_groupi_n_973 ,csa_tree_add_24_21_groupi_n_657 ,csa_tree_add_24_21_groupi_n_728);
  and csa_tree_add_24_21_groupi_g6597(csa_tree_add_24_21_groupi_n_972 ,csa_tree_add_24_21_groupi_n_549 ,csa_tree_add_24_21_groupi_n_742);
  and csa_tree_add_24_21_groupi_g6598(csa_tree_add_24_21_groupi_n_971 ,csa_tree_add_24_21_groupi_n_558 ,csa_tree_add_24_21_groupi_n_741);
  and csa_tree_add_24_21_groupi_g6599(csa_tree_add_24_21_groupi_n_970 ,csa_tree_add_24_21_groupi_n_570 ,csa_tree_add_24_21_groupi_n_699);
  and csa_tree_add_24_21_groupi_g6600(csa_tree_add_24_21_groupi_n_969 ,csa_tree_add_24_21_groupi_n_633 ,csa_tree_add_24_21_groupi_n_807);
  and csa_tree_add_24_21_groupi_g6601(csa_tree_add_24_21_groupi_n_968 ,csa_tree_add_24_21_groupi_n_632 ,csa_tree_add_24_21_groupi_n_737);
  and csa_tree_add_24_21_groupi_g6602(csa_tree_add_24_21_groupi_n_967 ,csa_tree_add_24_21_groupi_n_619 ,csa_tree_add_24_21_groupi_n_843);
  and csa_tree_add_24_21_groupi_g6603(csa_tree_add_24_21_groupi_n_966 ,csa_tree_add_24_21_groupi_n_620 ,csa_tree_add_24_21_groupi_n_735);
  and csa_tree_add_24_21_groupi_g6604(csa_tree_add_24_21_groupi_n_965 ,csa_tree_add_24_21_groupi_n_621 ,csa_tree_add_24_21_groupi_n_752);
  and csa_tree_add_24_21_groupi_g6605(csa_tree_add_24_21_groupi_n_964 ,csa_tree_add_24_21_groupi_n_644 ,csa_tree_add_24_21_groupi_n_802);
  or csa_tree_add_24_21_groupi_g6606(csa_tree_add_24_21_groupi_n_963 ,csa_tree_add_24_21_groupi_n_362 ,csa_tree_add_24_21_groupi_n_761);
  and csa_tree_add_24_21_groupi_g6607(csa_tree_add_24_21_groupi_n_962 ,csa_tree_add_24_21_groupi_n_659 ,csa_tree_add_24_21_groupi_n_754);
  or csa_tree_add_24_21_groupi_g6608(csa_tree_add_24_21_groupi_n_961 ,csa_tree_add_24_21_groupi_n_684 ,csa_tree_add_24_21_groupi_n_823);
  or csa_tree_add_24_21_groupi_g6609(csa_tree_add_24_21_groupi_n_959 ,csa_tree_add_24_21_groupi_n_682 ,csa_tree_add_24_21_groupi_n_822);
  and csa_tree_add_24_21_groupi_g6610(csa_tree_add_24_21_groupi_n_957 ,csa_tree_add_24_21_groupi_n_618 ,csa_tree_add_24_21_groupi_n_731);
  and csa_tree_add_24_21_groupi_g6611(csa_tree_add_24_21_groupi_n_956 ,csa_tree_add_24_21_groupi_n_551 ,csa_tree_add_24_21_groupi_n_697);
  and csa_tree_add_24_21_groupi_g6612(csa_tree_add_24_21_groupi_n_955 ,csa_tree_add_24_21_groupi_n_664 ,csa_tree_add_24_21_groupi_n_805);
  and csa_tree_add_24_21_groupi_g6613(csa_tree_add_24_21_groupi_n_953 ,csa_tree_add_24_21_groupi_n_622 ,csa_tree_add_24_21_groupi_n_696);
  or csa_tree_add_24_21_groupi_g6614(csa_tree_add_24_21_groupi_n_952 ,csa_tree_add_24_21_groupi_n_681 ,csa_tree_add_24_21_groupi_n_826);
  and csa_tree_add_24_21_groupi_g6615(csa_tree_add_24_21_groupi_n_950 ,csa_tree_add_24_21_groupi_n_636 ,csa_tree_add_24_21_groupi_n_755);
  and csa_tree_add_24_21_groupi_g6616(csa_tree_add_24_21_groupi_n_949 ,csa_tree_add_24_21_groupi_n_685 ,csa_tree_add_24_21_groupi_n_757);
  and csa_tree_add_24_21_groupi_g6617(csa_tree_add_24_21_groupi_n_948 ,csa_tree_add_24_21_groupi_n_635 ,csa_tree_add_24_21_groupi_n_800);
  or csa_tree_add_24_21_groupi_g6618(csa_tree_add_24_21_groupi_n_947 ,csa_tree_add_24_21_groupi_n_680 ,csa_tree_add_24_21_groupi_n_831);
  or csa_tree_add_24_21_groupi_g6619(csa_tree_add_24_21_groupi_n_945 ,csa_tree_add_24_21_groupi_n_677 ,csa_tree_add_24_21_groupi_n_827);
  and csa_tree_add_24_21_groupi_g6620(csa_tree_add_24_21_groupi_n_943 ,csa_tree_add_24_21_groupi_n_637 ,csa_tree_add_24_21_groupi_n_729);
  and csa_tree_add_24_21_groupi_g6621(csa_tree_add_24_21_groupi_n_941 ,csa_tree_add_24_21_groupi_n_564 ,csa_tree_add_24_21_groupi_n_751);
  and csa_tree_add_24_21_groupi_g6622(csa_tree_add_24_21_groupi_n_939 ,csa_tree_add_24_21_groupi_n_665 ,csa_tree_add_24_21_groupi_n_812);
  and csa_tree_add_24_21_groupi_g6623(csa_tree_add_24_21_groupi_n_938 ,csa_tree_add_24_21_groupi_n_647 ,csa_tree_add_24_21_groupi_n_749);
  and csa_tree_add_24_21_groupi_g6624(csa_tree_add_24_21_groupi_n_937 ,csa_tree_add_24_21_groupi_n_576 ,csa_tree_add_24_21_groupi_n_775);
  and csa_tree_add_24_21_groupi_g6625(csa_tree_add_24_21_groupi_n_935 ,csa_tree_add_24_21_groupi_n_662 ,csa_tree_add_24_21_groupi_n_804);
  and csa_tree_add_24_21_groupi_g6626(csa_tree_add_24_21_groupi_n_934 ,csa_tree_add_24_21_groupi_n_582 ,csa_tree_add_24_21_groupi_n_710);
  not csa_tree_add_24_21_groupi_g6627(csa_tree_add_24_21_groupi_n_925 ,csa_tree_add_24_21_groupi_n_924);
  not csa_tree_add_24_21_groupi_g6628(csa_tree_add_24_21_groupi_n_921 ,csa_tree_add_24_21_groupi_n_920);
  not csa_tree_add_24_21_groupi_g6629(csa_tree_add_24_21_groupi_n_909 ,csa_tree_add_24_21_groupi_n_908);
  not csa_tree_add_24_21_groupi_g6630(csa_tree_add_24_21_groupi_n_885 ,csa_tree_add_24_21_groupi_n_886);
  not csa_tree_add_24_21_groupi_g6631(csa_tree_add_24_21_groupi_n_883 ,csa_tree_add_24_21_groupi_n_884);
  not csa_tree_add_24_21_groupi_g6632(csa_tree_add_24_21_groupi_n_877 ,csa_tree_add_24_21_groupi_n_878);
  not csa_tree_add_24_21_groupi_g6633(csa_tree_add_24_21_groupi_n_875 ,csa_tree_add_24_21_groupi_n_876);
  not csa_tree_add_24_21_groupi_g6634(csa_tree_add_24_21_groupi_n_870 ,csa_tree_add_24_21_groupi_n_871);
  not csa_tree_add_24_21_groupi_g6635(csa_tree_add_24_21_groupi_n_866 ,csa_tree_add_24_21_groupi_n_867);
  not csa_tree_add_24_21_groupi_g6636(csa_tree_add_24_21_groupi_n_864 ,csa_tree_add_24_21_groupi_n_865);
  not csa_tree_add_24_21_groupi_g6637(csa_tree_add_24_21_groupi_n_862 ,csa_tree_add_24_21_groupi_n_861);
  not csa_tree_add_24_21_groupi_g6638(csa_tree_add_24_21_groupi_n_859 ,csa_tree_add_24_21_groupi_n_860);
  not csa_tree_add_24_21_groupi_g6639(csa_tree_add_24_21_groupi_n_856 ,csa_tree_add_24_21_groupi_n_857);
  or csa_tree_add_24_21_groupi_g6640(csa_tree_add_24_21_groupi_n_851 ,in3[30] ,csa_tree_add_24_21_groupi_n_844);
  xnor csa_tree_add_24_21_groupi_g6641(csa_tree_add_24_21_groupi_n_850 ,csa_tree_add_24_21_groupi_n_603 ,in3[8]);
  xnor csa_tree_add_24_21_groupi_g6642(csa_tree_add_24_21_groupi_n_849 ,csa_tree_add_24_21_groupi_n_601 ,in3[6]);
  xnor csa_tree_add_24_21_groupi_g6643(csa_tree_add_24_21_groupi_n_848 ,csa_tree_add_24_21_groupi_n_597 ,in3[10]);
  xnor csa_tree_add_24_21_groupi_g6644(csa_tree_add_24_21_groupi_n_847 ,csa_tree_add_24_21_groupi_n_605 ,in3[4]);
  xnor csa_tree_add_24_21_groupi_g6645(csa_tree_add_24_21_groupi_n_846 ,csa_tree_add_24_21_groupi_n_599 ,in3[12]);
  xnor csa_tree_add_24_21_groupi_g6646(csa_tree_add_24_21_groupi_n_845 ,csa_tree_add_24_21_groupi_n_595 ,in3[2]);
  and csa_tree_add_24_21_groupi_g6647(csa_tree_add_24_21_groupi_n_930 ,csa_tree_add_24_21_groupi_n_574 ,csa_tree_add_24_21_groupi_n_721);
  and csa_tree_add_24_21_groupi_g6648(csa_tree_add_24_21_groupi_n_929 ,csa_tree_add_24_21_groupi_n_548 ,csa_tree_add_24_21_groupi_n_711);
  or csa_tree_add_24_21_groupi_g6649(csa_tree_add_24_21_groupi_n_928 ,csa_tree_add_24_21_groupi_n_668 ,csa_tree_add_24_21_groupi_n_820);
  and csa_tree_add_24_21_groupi_g6650(csa_tree_add_24_21_groupi_n_927 ,csa_tree_add_24_21_groupi_n_578 ,csa_tree_add_24_21_groupi_n_723);
  and csa_tree_add_24_21_groupi_g6651(csa_tree_add_24_21_groupi_n_926 ,csa_tree_add_24_21_groupi_n_531 ,csa_tree_add_24_21_groupi_n_781);
  and csa_tree_add_24_21_groupi_g6652(csa_tree_add_24_21_groupi_n_924 ,csa_tree_add_24_21_groupi_n_547 ,csa_tree_add_24_21_groupi_n_782);
  and csa_tree_add_24_21_groupi_g6653(csa_tree_add_24_21_groupi_n_923 ,csa_tree_add_24_21_groupi_n_566 ,csa_tree_add_24_21_groupi_n_726);
  and csa_tree_add_24_21_groupi_g6654(csa_tree_add_24_21_groupi_n_922 ,csa_tree_add_24_21_groupi_n_541 ,csa_tree_add_24_21_groupi_n_795);
  and csa_tree_add_24_21_groupi_g6655(csa_tree_add_24_21_groupi_n_920 ,csa_tree_add_24_21_groupi_n_544 ,csa_tree_add_24_21_groupi_n_788);
  and csa_tree_add_24_21_groupi_g6656(csa_tree_add_24_21_groupi_n_919 ,csa_tree_add_24_21_groupi_n_661 ,csa_tree_add_24_21_groupi_n_714);
  and csa_tree_add_24_21_groupi_g6657(csa_tree_add_24_21_groupi_n_918 ,csa_tree_add_24_21_groupi_n_536 ,csa_tree_add_24_21_groupi_n_779);
  and csa_tree_add_24_21_groupi_g6658(csa_tree_add_24_21_groupi_n_917 ,csa_tree_add_24_21_groupi_n_542 ,csa_tree_add_24_21_groupi_n_785);
  and csa_tree_add_24_21_groupi_g6659(csa_tree_add_24_21_groupi_n_916 ,csa_tree_add_24_21_groupi_n_561 ,csa_tree_add_24_21_groupi_n_712);
  and csa_tree_add_24_21_groupi_g6660(csa_tree_add_24_21_groupi_n_915 ,csa_tree_add_24_21_groupi_n_533 ,csa_tree_add_24_21_groupi_n_780);
  and csa_tree_add_24_21_groupi_g6661(csa_tree_add_24_21_groupi_n_914 ,csa_tree_add_24_21_groupi_n_538 ,csa_tree_add_24_21_groupi_n_791);
  and csa_tree_add_24_21_groupi_g6662(csa_tree_add_24_21_groupi_n_913 ,csa_tree_add_24_21_groupi_n_553 ,csa_tree_add_24_21_groupi_n_704);
  and csa_tree_add_24_21_groupi_g6663(csa_tree_add_24_21_groupi_n_912 ,csa_tree_add_24_21_groupi_n_573 ,csa_tree_add_24_21_groupi_n_808);
  and csa_tree_add_24_21_groupi_g6664(csa_tree_add_24_21_groupi_n_911 ,csa_tree_add_24_21_groupi_n_660 ,csa_tree_add_24_21_groupi_n_707);
  and csa_tree_add_24_21_groupi_g6665(csa_tree_add_24_21_groupi_n_910 ,csa_tree_add_24_21_groupi_n_540 ,csa_tree_add_24_21_groupi_n_792);
  and csa_tree_add_24_21_groupi_g6666(csa_tree_add_24_21_groupi_n_908 ,csa_tree_add_24_21_groupi_n_537 ,csa_tree_add_24_21_groupi_n_793);
  and csa_tree_add_24_21_groupi_g6667(csa_tree_add_24_21_groupi_n_907 ,csa_tree_add_24_21_groupi_n_563 ,csa_tree_add_24_21_groupi_n_705);
  and csa_tree_add_24_21_groupi_g6668(csa_tree_add_24_21_groupi_n_906 ,csa_tree_add_24_21_groupi_n_545 ,csa_tree_add_24_21_groupi_n_794);
  and csa_tree_add_24_21_groupi_g6669(csa_tree_add_24_21_groupi_n_905 ,csa_tree_add_24_21_groupi_n_535 ,csa_tree_add_24_21_groupi_n_790);
  and csa_tree_add_24_21_groupi_g6670(csa_tree_add_24_21_groupi_n_904 ,csa_tree_add_24_21_groupi_n_539 ,csa_tree_add_24_21_groupi_n_786);
  and csa_tree_add_24_21_groupi_g6671(csa_tree_add_24_21_groupi_n_903 ,csa_tree_add_24_21_groupi_n_609 ,csa_tree_add_24_21_groupi_n_730);
  and csa_tree_add_24_21_groupi_g6672(csa_tree_add_24_21_groupi_n_902 ,csa_tree_add_24_21_groupi_n_613 ,csa_tree_add_24_21_groupi_n_771);
  and csa_tree_add_24_21_groupi_g6673(csa_tree_add_24_21_groupi_n_901 ,csa_tree_add_24_21_groupi_n_611 ,csa_tree_add_24_21_groupi_n_773);
  and csa_tree_add_24_21_groupi_g6674(csa_tree_add_24_21_groupi_n_900 ,csa_tree_add_24_21_groupi_n_615 ,csa_tree_add_24_21_groupi_n_803);
  and csa_tree_add_24_21_groupi_g6675(csa_tree_add_24_21_groupi_n_899 ,csa_tree_add_24_21_groupi_n_554 ,csa_tree_add_24_21_groupi_n_772);
  or csa_tree_add_24_21_groupi_g6676(csa_tree_add_24_21_groupi_n_898 ,csa_tree_add_24_21_groupi_n_606 ,csa_tree_add_24_21_groupi_n_695);
  or csa_tree_add_24_21_groupi_g6677(csa_tree_add_24_21_groupi_n_897 ,csa_tree_add_24_21_groupi_n_610 ,csa_tree_add_24_21_groupi_n_691);
  or csa_tree_add_24_21_groupi_g6678(csa_tree_add_24_21_groupi_n_896 ,csa_tree_add_24_21_groupi_n_336 ,csa_tree_add_24_21_groupi_n_769);
  and csa_tree_add_24_21_groupi_g6679(csa_tree_add_24_21_groupi_n_895 ,csa_tree_add_24_21_groupi_n_583 ,csa_tree_add_24_21_groupi_n_798);
  or csa_tree_add_24_21_groupi_g6680(csa_tree_add_24_21_groupi_n_894 ,csa_tree_add_24_21_groupi_n_614 ,csa_tree_add_24_21_groupi_n_690);
  or csa_tree_add_24_21_groupi_g6681(csa_tree_add_24_21_groupi_n_893 ,csa_tree_add_24_21_groupi_n_608 ,csa_tree_add_24_21_groupi_n_692);
  or csa_tree_add_24_21_groupi_g6682(csa_tree_add_24_21_groupi_n_892 ,csa_tree_add_24_21_groupi_n_612 ,csa_tree_add_24_21_groupi_n_693);
  and csa_tree_add_24_21_groupi_g6683(csa_tree_add_24_21_groupi_n_891 ,csa_tree_add_24_21_groupi_n_645 ,csa_tree_add_24_21_groupi_n_713);
  and csa_tree_add_24_21_groupi_g6684(csa_tree_add_24_21_groupi_n_890 ,csa_tree_add_24_21_groupi_n_550 ,csa_tree_add_24_21_groupi_n_709);
  and csa_tree_add_24_21_groupi_g6685(csa_tree_add_24_21_groupi_n_889 ,csa_tree_add_24_21_groupi_n_607 ,csa_tree_add_24_21_groupi_n_756);
  or csa_tree_add_24_21_groupi_g6686(csa_tree_add_24_21_groupi_n_888 ,csa_tree_add_24_21_groupi_n_361 ,csa_tree_add_24_21_groupi_n_765);
  and csa_tree_add_24_21_groupi_g6687(csa_tree_add_24_21_groupi_n_887 ,csa_tree_add_24_21_groupi_n_656 ,csa_tree_add_24_21_groupi_n_799);
  and csa_tree_add_24_21_groupi_g6688(csa_tree_add_24_21_groupi_n_886 ,csa_tree_add_24_21_groupi_n_625 ,csa_tree_add_24_21_groupi_n_703);
  or csa_tree_add_24_21_groupi_g6689(csa_tree_add_24_21_groupi_n_884 ,csa_tree_add_24_21_groupi_n_670 ,csa_tree_add_24_21_groupi_n_819);
  and csa_tree_add_24_21_groupi_g6690(csa_tree_add_24_21_groupi_n_882 ,csa_tree_add_24_21_groupi_n_648 ,csa_tree_add_24_21_groupi_n_698);
  and csa_tree_add_24_21_groupi_g6691(csa_tree_add_24_21_groupi_n_881 ,csa_tree_add_24_21_groupi_n_555 ,csa_tree_add_24_21_groupi_n_740);
  and csa_tree_add_24_21_groupi_g6692(csa_tree_add_24_21_groupi_n_880 ,csa_tree_add_24_21_groupi_n_557 ,csa_tree_add_24_21_groupi_n_718);
  and csa_tree_add_24_21_groupi_g6693(csa_tree_add_24_21_groupi_n_879 ,csa_tree_add_24_21_groupi_n_552 ,csa_tree_add_24_21_groupi_n_706);
  or csa_tree_add_24_21_groupi_g6694(csa_tree_add_24_21_groupi_n_878 ,csa_tree_add_24_21_groupi_n_672 ,csa_tree_add_24_21_groupi_n_828);
  and csa_tree_add_24_21_groupi_g6695(csa_tree_add_24_21_groupi_n_876 ,csa_tree_add_24_21_groupi_n_546 ,csa_tree_add_24_21_groupi_n_796);
  and csa_tree_add_24_21_groupi_g6696(csa_tree_add_24_21_groupi_n_874 ,csa_tree_add_24_21_groupi_n_623 ,csa_tree_add_24_21_groupi_n_814);
  and csa_tree_add_24_21_groupi_g6697(csa_tree_add_24_21_groupi_n_873 ,csa_tree_add_24_21_groupi_n_560 ,csa_tree_add_24_21_groupi_n_715);
  and csa_tree_add_24_21_groupi_g6698(csa_tree_add_24_21_groupi_n_872 ,csa_tree_add_24_21_groupi_n_584 ,csa_tree_add_24_21_groupi_n_725);
  or csa_tree_add_24_21_groupi_g6699(csa_tree_add_24_21_groupi_n_871 ,csa_tree_add_24_21_groupi_n_674 ,csa_tree_add_24_21_groupi_n_821);
  and csa_tree_add_24_21_groupi_g6700(csa_tree_add_24_21_groupi_n_869 ,csa_tree_add_24_21_groupi_n_534 ,csa_tree_add_24_21_groupi_n_787);
  and csa_tree_add_24_21_groupi_g6701(csa_tree_add_24_21_groupi_n_868 ,csa_tree_add_24_21_groupi_n_543 ,csa_tree_add_24_21_groupi_n_783);
  or csa_tree_add_24_21_groupi_g6702(csa_tree_add_24_21_groupi_n_867 ,csa_tree_add_24_21_groupi_n_669 ,csa_tree_add_24_21_groupi_n_816);
  and csa_tree_add_24_21_groupi_g6703(csa_tree_add_24_21_groupi_n_865 ,csa_tree_add_24_21_groupi_n_532 ,csa_tree_add_24_21_groupi_n_784);
  and csa_tree_add_24_21_groupi_g6704(csa_tree_add_24_21_groupi_n_863 ,csa_tree_add_24_21_groupi_n_666 ,csa_tree_add_24_21_groupi_n_717);
  or csa_tree_add_24_21_groupi_g6705(csa_tree_add_24_21_groupi_n_861 ,csa_tree_add_24_21_groupi_n_683 ,csa_tree_add_24_21_groupi_n_815);
  or csa_tree_add_24_21_groupi_g6706(csa_tree_add_24_21_groupi_n_860 ,csa_tree_add_24_21_groupi_n_673 ,csa_tree_add_24_21_groupi_n_824);
  and csa_tree_add_24_21_groupi_g6707(csa_tree_add_24_21_groupi_n_858 ,csa_tree_add_24_21_groupi_n_628 ,csa_tree_add_24_21_groupi_n_774);
  and csa_tree_add_24_21_groupi_g6708(csa_tree_add_24_21_groupi_n_857 ,csa_tree_add_24_21_groupi_n_658 ,csa_tree_add_24_21_groupi_n_811);
  and csa_tree_add_24_21_groupi_g6709(csa_tree_add_24_21_groupi_n_855 ,csa_tree_add_24_21_groupi_n_577 ,csa_tree_add_24_21_groupi_n_722);
  and csa_tree_add_24_21_groupi_g6710(csa_tree_add_24_21_groupi_n_854 ,csa_tree_add_24_21_groupi_n_579 ,csa_tree_add_24_21_groupi_n_801);
  or csa_tree_add_24_21_groupi_g6711(csa_tree_add_24_21_groupi_n_853 ,csa_tree_add_24_21_groupi_n_338 ,csa_tree_add_24_21_groupi_n_767);
  or csa_tree_add_24_21_groupi_g6712(csa_tree_add_24_21_groupi_n_852 ,csa_tree_add_24_21_groupi_n_360 ,csa_tree_add_24_21_groupi_n_763);
  or csa_tree_add_24_21_groupi_g6713(csa_tree_add_24_21_groupi_n_843 ,csa_tree_add_24_21_groupi_n_416 ,csa_tree_add_24_21_groupi_n_80);
  nor csa_tree_add_24_21_groupi_g6714(csa_tree_add_24_21_groupi_n_842 ,in3[10] ,csa_tree_add_24_21_groupi_n_596);
  or csa_tree_add_24_21_groupi_g6715(csa_tree_add_24_21_groupi_n_841 ,csa_tree_add_24_21_groupi_n_357 ,csa_tree_add_24_21_groupi_n_601);
  or csa_tree_add_24_21_groupi_g6716(csa_tree_add_24_21_groupi_n_840 ,csa_tree_add_24_21_groupi_n_359 ,csa_tree_add_24_21_groupi_n_603);
  nor csa_tree_add_24_21_groupi_g6717(csa_tree_add_24_21_groupi_n_839 ,in3[8] ,csa_tree_add_24_21_groupi_n_602);
  or csa_tree_add_24_21_groupi_g6718(csa_tree_add_24_21_groupi_n_838 ,csa_tree_add_24_21_groupi_n_356 ,csa_tree_add_24_21_groupi_n_597);
  nor csa_tree_add_24_21_groupi_g6719(csa_tree_add_24_21_groupi_n_837 ,in3[6] ,csa_tree_add_24_21_groupi_n_600);
  or csa_tree_add_24_21_groupi_g6720(csa_tree_add_24_21_groupi_n_836 ,csa_tree_add_24_21_groupi_n_333 ,csa_tree_add_24_21_groupi_n_605);
  or csa_tree_add_24_21_groupi_g6721(csa_tree_add_24_21_groupi_n_835 ,csa_tree_add_24_21_groupi_n_358 ,csa_tree_add_24_21_groupi_n_595);
  nor csa_tree_add_24_21_groupi_g6722(csa_tree_add_24_21_groupi_n_834 ,in3[2] ,csa_tree_add_24_21_groupi_n_594);
  nor csa_tree_add_24_21_groupi_g6723(csa_tree_add_24_21_groupi_n_833 ,in3[12] ,csa_tree_add_24_21_groupi_n_598);
  or csa_tree_add_24_21_groupi_g6724(csa_tree_add_24_21_groupi_n_832 ,csa_tree_add_24_21_groupi_n_334 ,csa_tree_add_24_21_groupi_n_599);
  and csa_tree_add_24_21_groupi_g6725(csa_tree_add_24_21_groupi_n_831 ,in2[5] ,csa_tree_add_24_21_groupi_n_281);
  and csa_tree_add_24_21_groupi_g6726(csa_tree_add_24_21_groupi_n_830 ,in2[2] ,csa_tree_add_24_21_groupi_n_281);
  and csa_tree_add_24_21_groupi_g6727(csa_tree_add_24_21_groupi_n_829 ,in2[1] ,csa_tree_add_24_21_groupi_n_277);
  and csa_tree_add_24_21_groupi_g6728(csa_tree_add_24_21_groupi_n_828 ,in2[8] ,csa_tree_add_24_21_groupi_n_277);
  and csa_tree_add_24_21_groupi_g6729(csa_tree_add_24_21_groupi_n_827 ,in2[15] ,csa_tree_add_24_21_groupi_n_281);
  and csa_tree_add_24_21_groupi_g6730(csa_tree_add_24_21_groupi_n_826 ,in2[10] ,csa_tree_add_24_21_groupi_n_281);
  and csa_tree_add_24_21_groupi_g6731(csa_tree_add_24_21_groupi_n_825 ,in2[6] ,csa_tree_add_24_21_groupi_n_281);
  and csa_tree_add_24_21_groupi_g6732(csa_tree_add_24_21_groupi_n_824 ,in2[11] ,csa_tree_add_24_21_groupi_n_281);
  and csa_tree_add_24_21_groupi_g6733(csa_tree_add_24_21_groupi_n_823 ,in2[12] ,csa_tree_add_24_21_groupi_n_281);
  and csa_tree_add_24_21_groupi_g6734(csa_tree_add_24_21_groupi_n_822 ,in2[13] ,csa_tree_add_24_21_groupi_n_278);
  and csa_tree_add_24_21_groupi_g6735(csa_tree_add_24_21_groupi_n_821 ,in2[9] ,csa_tree_add_24_21_groupi_n_278);
  and csa_tree_add_24_21_groupi_g6736(csa_tree_add_24_21_groupi_n_820 ,in2[14] ,csa_tree_add_24_21_groupi_n_254);
  and csa_tree_add_24_21_groupi_g6737(csa_tree_add_24_21_groupi_n_819 ,in2[3] ,csa_tree_add_24_21_groupi_n_254);
  or csa_tree_add_24_21_groupi_g6738(csa_tree_add_24_21_groupi_n_818 ,csa_tree_add_24_21_groupi_n_346 ,csa_tree_add_24_21_groupi_n_279);
  or csa_tree_add_24_21_groupi_g6739(csa_tree_add_24_21_groupi_n_817 ,csa_tree_add_24_21_groupi_n_524 ,csa_tree_add_24_21_groupi_n_77);
  and csa_tree_add_24_21_groupi_g6740(csa_tree_add_24_21_groupi_n_816 ,in2[16] ,csa_tree_add_24_21_groupi_n_281);
  and csa_tree_add_24_21_groupi_g6741(csa_tree_add_24_21_groupi_n_815 ,in2[4] ,csa_tree_add_24_21_groupi_n_281);
  or csa_tree_add_24_21_groupi_g6742(csa_tree_add_24_21_groupi_n_814 ,csa_tree_add_24_21_groupi_n_423 ,csa_tree_add_24_21_groupi_n_220);
  or csa_tree_add_24_21_groupi_g6743(csa_tree_add_24_21_groupi_n_813 ,csa_tree_add_24_21_groupi_n_419 ,csa_tree_add_24_21_groupi_n_220);
  or csa_tree_add_24_21_groupi_g6744(csa_tree_add_24_21_groupi_n_812 ,csa_tree_add_24_21_groupi_n_408 ,csa_tree_add_24_21_groupi_n_220);
  or csa_tree_add_24_21_groupi_g6745(csa_tree_add_24_21_groupi_n_811 ,csa_tree_add_24_21_groupi_n_410 ,csa_tree_add_24_21_groupi_n_57);
  or csa_tree_add_24_21_groupi_g6746(csa_tree_add_24_21_groupi_n_810 ,csa_tree_add_24_21_groupi_n_420 ,csa_tree_add_24_21_groupi_n_57);
  or csa_tree_add_24_21_groupi_g6747(csa_tree_add_24_21_groupi_n_809 ,csa_tree_add_24_21_groupi_n_417 ,csa_tree_add_24_21_groupi_n_57);
  or csa_tree_add_24_21_groupi_g6748(csa_tree_add_24_21_groupi_n_808 ,csa_tree_add_24_21_groupi_n_414 ,csa_tree_add_24_21_groupi_n_39);
  or csa_tree_add_24_21_groupi_g6749(csa_tree_add_24_21_groupi_n_807 ,csa_tree_add_24_21_groupi_n_413 ,csa_tree_add_24_21_groupi_n_57);
  nor csa_tree_add_24_21_groupi_g6750(csa_tree_add_24_21_groupi_n_806 ,in3[4] ,csa_tree_add_24_21_groupi_n_604);
  or csa_tree_add_24_21_groupi_g6751(csa_tree_add_24_21_groupi_n_805 ,csa_tree_add_24_21_groupi_n_412 ,csa_tree_add_24_21_groupi_n_81);
  or csa_tree_add_24_21_groupi_g6752(csa_tree_add_24_21_groupi_n_804 ,csa_tree_add_24_21_groupi_n_393 ,csa_tree_add_24_21_groupi_n_57);
  or csa_tree_add_24_21_groupi_g6753(csa_tree_add_24_21_groupi_n_803 ,csa_tree_add_24_21_groupi_n_422 ,csa_tree_add_24_21_groupi_n_57);
  or csa_tree_add_24_21_groupi_g6754(csa_tree_add_24_21_groupi_n_802 ,csa_tree_add_24_21_groupi_n_425 ,csa_tree_add_24_21_groupi_n_39);
  or csa_tree_add_24_21_groupi_g6755(csa_tree_add_24_21_groupi_n_801 ,csa_tree_add_24_21_groupi_n_409 ,csa_tree_add_24_21_groupi_n_57);
  or csa_tree_add_24_21_groupi_g6756(csa_tree_add_24_21_groupi_n_800 ,csa_tree_add_24_21_groupi_n_424 ,csa_tree_add_24_21_groupi_n_80);
  or csa_tree_add_24_21_groupi_g6757(csa_tree_add_24_21_groupi_n_799 ,csa_tree_add_24_21_groupi_n_407 ,csa_tree_add_24_21_groupi_n_57);
  or csa_tree_add_24_21_groupi_g6758(csa_tree_add_24_21_groupi_n_798 ,csa_tree_add_24_21_groupi_n_411 ,csa_tree_add_24_21_groupi_n_57);
  or csa_tree_add_24_21_groupi_g6759(csa_tree_add_24_21_groupi_n_797 ,csa_tree_add_24_21_groupi_n_418 ,csa_tree_add_24_21_groupi_n_57);
  or csa_tree_add_24_21_groupi_g6760(csa_tree_add_24_21_groupi_n_796 ,csa_tree_add_24_21_groupi_n_430 ,csa_tree_add_24_21_groupi_n_69);
  or csa_tree_add_24_21_groupi_g6761(csa_tree_add_24_21_groupi_n_795 ,csa_tree_add_24_21_groupi_n_395 ,csa_tree_add_24_21_groupi_n_3);
  or csa_tree_add_24_21_groupi_g6762(csa_tree_add_24_21_groupi_n_794 ,csa_tree_add_24_21_groupi_n_440 ,csa_tree_add_24_21_groupi_n_69);
  or csa_tree_add_24_21_groupi_g6763(csa_tree_add_24_21_groupi_n_793 ,csa_tree_add_24_21_groupi_n_438 ,csa_tree_add_24_21_groupi_n_69);
  or csa_tree_add_24_21_groupi_g6764(csa_tree_add_24_21_groupi_n_792 ,csa_tree_add_24_21_groupi_n_434 ,csa_tree_add_24_21_groupi_n_69);
  or csa_tree_add_24_21_groupi_g6765(csa_tree_add_24_21_groupi_n_791 ,csa_tree_add_24_21_groupi_n_431 ,csa_tree_add_24_21_groupi_n_119);
  or csa_tree_add_24_21_groupi_g6766(csa_tree_add_24_21_groupi_n_790 ,csa_tree_add_24_21_groupi_n_439 ,csa_tree_add_24_21_groupi_n_69);
  nor csa_tree_add_24_21_groupi_g6767(csa_tree_add_24_21_groupi_n_789 ,csa_tree_add_24_21_groupi_n_214 ,csa_tree_add_24_21_groupi_n_437);
  or csa_tree_add_24_21_groupi_g6768(csa_tree_add_24_21_groupi_n_788 ,csa_tree_add_24_21_groupi_n_432 ,csa_tree_add_24_21_groupi_n_120);
  or csa_tree_add_24_21_groupi_g6769(csa_tree_add_24_21_groupi_n_787 ,csa_tree_add_24_21_groupi_n_429 ,csa_tree_add_24_21_groupi_n_69);
  or csa_tree_add_24_21_groupi_g6770(csa_tree_add_24_21_groupi_n_786 ,csa_tree_add_24_21_groupi_n_442 ,csa_tree_add_24_21_groupi_n_214);
  or csa_tree_add_24_21_groupi_g6771(csa_tree_add_24_21_groupi_n_785 ,csa_tree_add_24_21_groupi_n_436 ,csa_tree_add_24_21_groupi_n_69);
  or csa_tree_add_24_21_groupi_g6772(csa_tree_add_24_21_groupi_n_784 ,csa_tree_add_24_21_groupi_n_426 ,csa_tree_add_24_21_groupi_n_3);
  or csa_tree_add_24_21_groupi_g6773(csa_tree_add_24_21_groupi_n_783 ,csa_tree_add_24_21_groupi_n_428 ,csa_tree_add_24_21_groupi_n_69);
  or csa_tree_add_24_21_groupi_g6774(csa_tree_add_24_21_groupi_n_782 ,csa_tree_add_24_21_groupi_n_421 ,csa_tree_add_24_21_groupi_n_214);
  or csa_tree_add_24_21_groupi_g6775(csa_tree_add_24_21_groupi_n_781 ,csa_tree_add_24_21_groupi_n_427 ,csa_tree_add_24_21_groupi_n_119);
  or csa_tree_add_24_21_groupi_g6776(csa_tree_add_24_21_groupi_n_780 ,csa_tree_add_24_21_groupi_n_443 ,csa_tree_add_24_21_groupi_n_69);
  or csa_tree_add_24_21_groupi_g6777(csa_tree_add_24_21_groupi_n_779 ,csa_tree_add_24_21_groupi_n_435 ,csa_tree_add_24_21_groupi_n_69);
  or csa_tree_add_24_21_groupi_g6778(csa_tree_add_24_21_groupi_n_778 ,csa_tree_add_24_21_groupi_n_452 ,csa_tree_add_24_21_groupi_n_205);
  or csa_tree_add_24_21_groupi_g6779(csa_tree_add_24_21_groupi_n_777 ,csa_tree_add_24_21_groupi_n_495 ,csa_tree_add_24_21_groupi_n_211);
  or csa_tree_add_24_21_groupi_g6780(csa_tree_add_24_21_groupi_n_776 ,csa_tree_add_24_21_groupi_n_465 ,csa_tree_add_24_21_groupi_n_86);
  or csa_tree_add_24_21_groupi_g6781(csa_tree_add_24_21_groupi_n_775 ,csa_tree_add_24_21_groupi_n_497 ,csa_tree_add_24_21_groupi_n_217);
  or csa_tree_add_24_21_groupi_g6782(csa_tree_add_24_21_groupi_n_774 ,csa_tree_add_24_21_groupi_n_485 ,csa_tree_add_24_21_groupi_n_205);
  or csa_tree_add_24_21_groupi_g6783(csa_tree_add_24_21_groupi_n_773 ,csa_tree_add_24_21_groupi_n_459 ,csa_tree_add_24_21_groupi_n_75);
  or csa_tree_add_24_21_groupi_g6784(csa_tree_add_24_21_groupi_n_772 ,csa_tree_add_24_21_groupi_n_522 ,csa_tree_add_24_21_groupi_n_74);
  or csa_tree_add_24_21_groupi_g6785(csa_tree_add_24_21_groupi_n_771 ,csa_tree_add_24_21_groupi_n_529 ,csa_tree_add_24_21_groupi_n_205);
  or csa_tree_add_24_21_groupi_g6786(csa_tree_add_24_21_groupi_n_770 ,csa_tree_add_24_21_groupi_n_513 ,csa_tree_add_24_21_groupi_n_74);
  or csa_tree_add_24_21_groupi_g6787(csa_tree_add_24_21_groupi_n_844 ,csa_tree_add_24_21_groupi_n_327 ,csa_tree_add_24_21_groupi_n_279);
  not csa_tree_add_24_21_groupi_g6788(csa_tree_add_24_21_groupi_n_769 ,csa_tree_add_24_21_groupi_n_768);
  not csa_tree_add_24_21_groupi_g6789(csa_tree_add_24_21_groupi_n_767 ,csa_tree_add_24_21_groupi_n_766);
  not csa_tree_add_24_21_groupi_g6790(csa_tree_add_24_21_groupi_n_765 ,csa_tree_add_24_21_groupi_n_764);
  not csa_tree_add_24_21_groupi_g6791(csa_tree_add_24_21_groupi_n_763 ,csa_tree_add_24_21_groupi_n_762);
  not csa_tree_add_24_21_groupi_g6792(csa_tree_add_24_21_groupi_n_761 ,csa_tree_add_24_21_groupi_n_760);
  not csa_tree_add_24_21_groupi_g6793(csa_tree_add_24_21_groupi_n_758 ,csa_tree_add_24_21_groupi_n_759);
  or csa_tree_add_24_21_groupi_g6794(csa_tree_add_24_21_groupi_n_757 ,csa_tree_add_24_21_groupi_n_528 ,csa_tree_add_24_21_groupi_n_85);
  or csa_tree_add_24_21_groupi_g6795(csa_tree_add_24_21_groupi_n_756 ,csa_tree_add_24_21_groupi_n_489 ,csa_tree_add_24_21_groupi_n_85);
  or csa_tree_add_24_21_groupi_g6796(csa_tree_add_24_21_groupi_n_755 ,csa_tree_add_24_21_groupi_n_519 ,csa_tree_add_24_21_groupi_n_63);
  or csa_tree_add_24_21_groupi_g6797(csa_tree_add_24_21_groupi_n_754 ,csa_tree_add_24_21_groupi_n_446 ,csa_tree_add_24_21_groupi_n_60);
  or csa_tree_add_24_21_groupi_g6798(csa_tree_add_24_21_groupi_n_753 ,csa_tree_add_24_21_groupi_n_520 ,csa_tree_add_24_21_groupi_n_66);
  or csa_tree_add_24_21_groupi_g6799(csa_tree_add_24_21_groupi_n_752 ,csa_tree_add_24_21_groupi_n_487 ,csa_tree_add_24_21_groupi_n_60);
  or csa_tree_add_24_21_groupi_g6800(csa_tree_add_24_21_groupi_n_751 ,csa_tree_add_24_21_groupi_n_527 ,csa_tree_add_24_21_groupi_n_91);
  or csa_tree_add_24_21_groupi_g6801(csa_tree_add_24_21_groupi_n_750 ,csa_tree_add_24_21_groupi_n_510 ,csa_tree_add_24_21_groupi_n_66);
  or csa_tree_add_24_21_groupi_g6802(csa_tree_add_24_21_groupi_n_749 ,csa_tree_add_24_21_groupi_n_516 ,csa_tree_add_24_21_groupi_n_66);
  or csa_tree_add_24_21_groupi_g6803(csa_tree_add_24_21_groupi_n_748 ,csa_tree_add_24_21_groupi_n_512 ,csa_tree_add_24_21_groupi_n_63);
  or csa_tree_add_24_21_groupi_g6804(csa_tree_add_24_21_groupi_n_747 ,csa_tree_add_24_21_groupi_n_515 ,csa_tree_add_24_21_groupi_n_208);
  or csa_tree_add_24_21_groupi_g6805(csa_tree_add_24_21_groupi_n_746 ,csa_tree_add_24_21_groupi_n_457 ,csa_tree_add_24_21_groupi_n_60);
  or csa_tree_add_24_21_groupi_g6806(csa_tree_add_24_21_groupi_n_745 ,csa_tree_add_24_21_groupi_n_498 ,csa_tree_add_24_21_groupi_n_208);
  or csa_tree_add_24_21_groupi_g6807(csa_tree_add_24_21_groupi_n_744 ,csa_tree_add_24_21_groupi_n_500 ,csa_tree_add_24_21_groupi_n_208);
  or csa_tree_add_24_21_groupi_g6808(csa_tree_add_24_21_groupi_n_743 ,csa_tree_add_24_21_groupi_n_505 ,csa_tree_add_24_21_groupi_n_63);
  or csa_tree_add_24_21_groupi_g6809(csa_tree_add_24_21_groupi_n_742 ,csa_tree_add_24_21_groupi_n_445 ,csa_tree_add_24_21_groupi_n_41);
  or csa_tree_add_24_21_groupi_g6810(csa_tree_add_24_21_groupi_n_741 ,csa_tree_add_24_21_groupi_n_503 ,csa_tree_add_24_21_groupi_n_66);
  or csa_tree_add_24_21_groupi_g6811(csa_tree_add_24_21_groupi_n_740 ,csa_tree_add_24_21_groupi_n_458 ,csa_tree_add_24_21_groupi_n_60);
  or csa_tree_add_24_21_groupi_g6812(csa_tree_add_24_21_groupi_n_739 ,csa_tree_add_24_21_groupi_n_509 ,csa_tree_add_24_21_groupi_n_78);
  or csa_tree_add_24_21_groupi_g6813(csa_tree_add_24_21_groupi_n_738 ,csa_tree_add_24_21_groupi_n_499 ,csa_tree_add_24_21_groupi_n_34);
  or csa_tree_add_24_21_groupi_g6814(csa_tree_add_24_21_groupi_n_737 ,csa_tree_add_24_21_groupi_n_491 ,csa_tree_add_24_21_groupi_n_72);
  or csa_tree_add_24_21_groupi_g6815(csa_tree_add_24_21_groupi_n_736 ,csa_tree_add_24_21_groupi_n_496 ,csa_tree_add_24_21_groupi_n_63);
  or csa_tree_add_24_21_groupi_g6816(csa_tree_add_24_21_groupi_n_735 ,csa_tree_add_24_21_groupi_n_453 ,csa_tree_add_24_21_groupi_n_66);
  or csa_tree_add_24_21_groupi_g6817(csa_tree_add_24_21_groupi_n_734 ,csa_tree_add_24_21_groupi_n_517 ,csa_tree_add_24_21_groupi_n_66);
  or csa_tree_add_24_21_groupi_g6818(csa_tree_add_24_21_groupi_n_733 ,csa_tree_add_24_21_groupi_n_483 ,csa_tree_add_24_21_groupi_n_41);
  or csa_tree_add_24_21_groupi_g6819(csa_tree_add_24_21_groupi_n_732 ,csa_tree_add_24_21_groupi_n_514 ,csa_tree_add_24_21_groupi_n_43);
  or csa_tree_add_24_21_groupi_g6820(csa_tree_add_24_21_groupi_n_731 ,csa_tree_add_24_21_groupi_n_493 ,csa_tree_add_24_21_groupi_n_217);
  or csa_tree_add_24_21_groupi_g6821(csa_tree_add_24_21_groupi_n_730 ,csa_tree_add_24_21_groupi_n_502 ,csa_tree_add_24_21_groupi_n_72);
  or csa_tree_add_24_21_groupi_g6822(csa_tree_add_24_21_groupi_n_729 ,csa_tree_add_24_21_groupi_n_433 ,csa_tree_add_24_21_groupi_n_72);
  or csa_tree_add_24_21_groupi_g6823(csa_tree_add_24_21_groupi_n_728 ,csa_tree_add_24_21_groupi_n_507 ,csa_tree_add_24_21_groupi_n_30);
  or csa_tree_add_24_21_groupi_g6824(csa_tree_add_24_21_groupi_n_727 ,csa_tree_add_24_21_groupi_n_494 ,csa_tree_add_24_21_groupi_n_72);
  or csa_tree_add_24_21_groupi_g6825(csa_tree_add_24_21_groupi_n_726 ,csa_tree_add_24_21_groupi_n_525 ,csa_tree_add_24_21_groupi_n_92);
  or csa_tree_add_24_21_groupi_g6826(csa_tree_add_24_21_groupi_n_725 ,csa_tree_add_24_21_groupi_n_530 ,csa_tree_add_24_21_groupi_n_63);
  or csa_tree_add_24_21_groupi_g6827(csa_tree_add_24_21_groupi_n_724 ,csa_tree_add_24_21_groupi_n_511 ,csa_tree_add_24_21_groupi_n_63);
  or csa_tree_add_24_21_groupi_g6828(csa_tree_add_24_21_groupi_n_723 ,csa_tree_add_24_21_groupi_n_441 ,csa_tree_add_24_21_groupi_n_63);
  or csa_tree_add_24_21_groupi_g6829(csa_tree_add_24_21_groupi_n_722 ,csa_tree_add_24_21_groupi_n_448 ,csa_tree_add_24_21_groupi_n_211);
  or csa_tree_add_24_21_groupi_g6830(csa_tree_add_24_21_groupi_n_721 ,csa_tree_add_24_21_groupi_n_455 ,csa_tree_add_24_21_groupi_n_66);
  or csa_tree_add_24_21_groupi_g6831(csa_tree_add_24_21_groupi_n_720 ,csa_tree_add_24_21_groupi_n_449 ,csa_tree_add_24_21_groupi_n_72);
  or csa_tree_add_24_21_groupi_g6832(csa_tree_add_24_21_groupi_n_719 ,csa_tree_add_24_21_groupi_n_454 ,csa_tree_add_24_21_groupi_n_43);
  or csa_tree_add_24_21_groupi_g6833(csa_tree_add_24_21_groupi_n_718 ,csa_tree_add_24_21_groupi_n_394 ,csa_tree_add_24_21_groupi_n_77);
  or csa_tree_add_24_21_groupi_g6834(csa_tree_add_24_21_groupi_n_717 ,csa_tree_add_24_21_groupi_n_488 ,csa_tree_add_24_21_groupi_n_60);
  or csa_tree_add_24_21_groupi_g6835(csa_tree_add_24_21_groupi_n_716 ,csa_tree_add_24_21_groupi_n_521 ,csa_tree_add_24_21_groupi_n_72);
  or csa_tree_add_24_21_groupi_g6836(csa_tree_add_24_21_groupi_n_715 ,csa_tree_add_24_21_groupi_n_486 ,csa_tree_add_24_21_groupi_n_60);
  or csa_tree_add_24_21_groupi_g6837(csa_tree_add_24_21_groupi_n_714 ,csa_tree_add_24_21_groupi_n_447 ,csa_tree_add_24_21_groupi_n_217);
  or csa_tree_add_24_21_groupi_g6838(csa_tree_add_24_21_groupi_n_713 ,csa_tree_add_24_21_groupi_n_506 ,csa_tree_add_24_21_groupi_n_66);
  or csa_tree_add_24_21_groupi_g6839(csa_tree_add_24_21_groupi_n_712 ,csa_tree_add_24_21_groupi_n_484 ,csa_tree_add_24_21_groupi_n_60);
  or csa_tree_add_24_21_groupi_g6840(csa_tree_add_24_21_groupi_n_711 ,csa_tree_add_24_21_groupi_n_501 ,csa_tree_add_24_21_groupi_n_66);
  or csa_tree_add_24_21_groupi_g6841(csa_tree_add_24_21_groupi_n_710 ,csa_tree_add_24_21_groupi_n_490 ,csa_tree_add_24_21_groupi_n_30);
  or csa_tree_add_24_21_groupi_g6842(csa_tree_add_24_21_groupi_n_709 ,csa_tree_add_24_21_groupi_n_450 ,csa_tree_add_24_21_groupi_n_34);
  or csa_tree_add_24_21_groupi_g6843(csa_tree_add_24_21_groupi_n_708 ,csa_tree_add_24_21_groupi_n_523 ,csa_tree_add_24_21_groupi_n_72);
  or csa_tree_add_24_21_groupi_g6844(csa_tree_add_24_21_groupi_n_707 ,csa_tree_add_24_21_groupi_n_464 ,csa_tree_add_24_21_groupi_n_63);
  or csa_tree_add_24_21_groupi_g6845(csa_tree_add_24_21_groupi_n_706 ,csa_tree_add_24_21_groupi_n_451 ,csa_tree_add_24_21_groupi_n_211);
  or csa_tree_add_24_21_groupi_g6846(csa_tree_add_24_21_groupi_n_705 ,csa_tree_add_24_21_groupi_n_444 ,csa_tree_add_24_21_groupi_n_91);
  or csa_tree_add_24_21_groupi_g6847(csa_tree_add_24_21_groupi_n_704 ,csa_tree_add_24_21_groupi_n_518 ,csa_tree_add_24_21_groupi_n_66);
  or csa_tree_add_24_21_groupi_g6848(csa_tree_add_24_21_groupi_n_703 ,csa_tree_add_24_21_groupi_n_504 ,csa_tree_add_24_21_groupi_n_72);
  or csa_tree_add_24_21_groupi_g6849(csa_tree_add_24_21_groupi_n_702 ,csa_tree_add_24_21_groupi_n_456 ,csa_tree_add_24_21_groupi_n_63);
  or csa_tree_add_24_21_groupi_g6850(csa_tree_add_24_21_groupi_n_701 ,csa_tree_add_24_21_groupi_n_415 ,csa_tree_add_24_21_groupi_n_63);
  or csa_tree_add_24_21_groupi_g6851(csa_tree_add_24_21_groupi_n_700 ,csa_tree_add_24_21_groupi_n_526 ,csa_tree_add_24_21_groupi_n_72);
  or csa_tree_add_24_21_groupi_g6852(csa_tree_add_24_21_groupi_n_699 ,csa_tree_add_24_21_groupi_n_460 ,csa_tree_add_24_21_groupi_n_60);
  or csa_tree_add_24_21_groupi_g6853(csa_tree_add_24_21_groupi_n_698 ,csa_tree_add_24_21_groupi_n_466 ,csa_tree_add_24_21_groupi_n_72);
  or csa_tree_add_24_21_groupi_g6854(csa_tree_add_24_21_groupi_n_697 ,csa_tree_add_24_21_groupi_n_492 ,csa_tree_add_24_21_groupi_n_60);
  or csa_tree_add_24_21_groupi_g6855(csa_tree_add_24_21_groupi_n_696 ,csa_tree_add_24_21_groupi_n_508 ,csa_tree_add_24_21_groupi_n_60);
  nor csa_tree_add_24_21_groupi_g6856(csa_tree_add_24_21_groupi_n_695 ,csa_tree_add_24_21_groupi_n_60 ,csa_tree_add_22_22_n_102);
  nor csa_tree_add_24_21_groupi_g6857(csa_tree_add_24_21_groupi_n_694 ,csa_tree_add_24_21_groupi_n_325 ,csa_tree_add_24_21_groupi_n_279);
  nor csa_tree_add_24_21_groupi_g6858(csa_tree_add_24_21_groupi_n_693 ,csa_tree_add_24_21_groupi_n_66 ,csa_tree_add_22_22_n_103);
  nor csa_tree_add_24_21_groupi_g6859(csa_tree_add_24_21_groupi_n_692 ,csa_tree_add_24_21_groupi_n_72 ,csa_tree_add_22_22_n_114);
  nor csa_tree_add_24_21_groupi_g6860(csa_tree_add_24_21_groupi_n_691 ,csa_tree_add_24_21_groupi_n_63 ,csa_tree_add_22_22_n_100);
  nor csa_tree_add_24_21_groupi_g6861(csa_tree_add_24_21_groupi_n_690 ,csa_tree_add_24_21_groupi_n_57 ,csa_tree_add_22_22_n_118);
  nor csa_tree_add_24_21_groupi_g6862(csa_tree_add_24_21_groupi_n_689 ,csa_tree_add_24_21_groupi_n_69 ,csa_tree_add_22_22_n_101);
  and csa_tree_add_24_21_groupi_g6863(csa_tree_add_24_21_groupi_n_768 ,in1[3] ,csa_tree_add_24_21_groupi_n_630);
  and csa_tree_add_24_21_groupi_g6864(csa_tree_add_24_21_groupi_n_766 ,in1[9] ,csa_tree_add_24_21_groupi_n_575);
  and csa_tree_add_24_21_groupi_g6865(csa_tree_add_24_21_groupi_n_764 ,in1[5] ,csa_tree_add_24_21_groupi_n_667);
  and csa_tree_add_24_21_groupi_g6866(csa_tree_add_24_21_groupi_n_762 ,in1[11] ,csa_tree_add_24_21_groupi_n_616);
  and csa_tree_add_24_21_groupi_g6867(csa_tree_add_24_21_groupi_n_760 ,in1[7] ,csa_tree_add_24_21_groupi_n_638);
  xnor csa_tree_add_24_21_groupi_g6868(csa_tree_add_24_21_groupi_n_759 ,csa_tree_add_24_21_groupi_n_482 ,in3[1]);
  not csa_tree_add_24_21_groupi_g6869(csa_tree_add_24_21_groupi_n_687 ,csa_tree_add_24_21_groupi_n_688);
  or csa_tree_add_24_21_groupi_g6870(csa_tree_add_24_21_groupi_n_685 ,csa_tree_add_24_21_groupi_n_269 ,csa_tree_add_24_21_groupi_n_446);
  and csa_tree_add_24_21_groupi_g6871(csa_tree_add_24_21_groupi_n_684 ,in2[13] ,csa_tree_add_24_21_groupi_n_293);
  and csa_tree_add_24_21_groupi_g6872(csa_tree_add_24_21_groupi_n_683 ,in2[5] ,csa_tree_add_24_21_groupi_n_293);
  and csa_tree_add_24_21_groupi_g6873(csa_tree_add_24_21_groupi_n_682 ,in2[14] ,csa_tree_add_24_21_groupi_n_293);
  and csa_tree_add_24_21_groupi_g6874(csa_tree_add_24_21_groupi_n_681 ,in2[11] ,csa_tree_add_24_21_groupi_n_404);
  and csa_tree_add_24_21_groupi_g6875(csa_tree_add_24_21_groupi_n_680 ,in2[6] ,csa_tree_add_24_21_groupi_n_293);
  and csa_tree_add_24_21_groupi_g6876(csa_tree_add_24_21_groupi_n_679 ,in2[2] ,csa_tree_add_24_21_groupi_n_404);
  nor csa_tree_add_24_21_groupi_g6877(csa_tree_add_24_21_groupi_n_678 ,csa_tree_add_24_21_groupi_n_346 ,csa_tree_add_24_21_groupi_n_200);
  and csa_tree_add_24_21_groupi_g6878(csa_tree_add_24_21_groupi_n_677 ,in2[16] ,csa_tree_add_24_21_groupi_n_293);
  and csa_tree_add_24_21_groupi_g6879(csa_tree_add_24_21_groupi_n_676 ,in2[1] ,csa_tree_add_24_21_groupi_n_404);
  and csa_tree_add_24_21_groupi_g6880(csa_tree_add_24_21_groupi_n_675 ,in2[3] ,csa_tree_add_24_21_groupi_n_293);
  and csa_tree_add_24_21_groupi_g6881(csa_tree_add_24_21_groupi_n_674 ,in2[10] ,csa_tree_add_24_21_groupi_n_293);
  and csa_tree_add_24_21_groupi_g6882(csa_tree_add_24_21_groupi_n_673 ,in2[12] ,csa_tree_add_24_21_groupi_n_293);
  and csa_tree_add_24_21_groupi_g6883(csa_tree_add_24_21_groupi_n_672 ,in2[9] ,csa_tree_add_24_21_groupi_n_293);
  or csa_tree_add_24_21_groupi_g6884(csa_tree_add_24_21_groupi_n_671 ,csa_tree_add_24_21_groupi_n_347 ,csa_tree_add_24_21_groupi_n_200);
  and csa_tree_add_24_21_groupi_g6885(csa_tree_add_24_21_groupi_n_670 ,in2[4] ,csa_tree_add_24_21_groupi_n_293);
  nor csa_tree_add_24_21_groupi_g6886(csa_tree_add_24_21_groupi_n_669 ,csa_tree_add_24_21_groupi_n_327 ,csa_tree_add_24_21_groupi_n_200);
  and csa_tree_add_24_21_groupi_g6887(csa_tree_add_24_21_groupi_n_668 ,in2[15] ,csa_tree_add_24_21_groupi_n_293);
  or csa_tree_add_24_21_groupi_g6888(csa_tree_add_24_21_groupi_n_667 ,csa_tree_add_24_21_groupi_n_381 ,csa_tree_add_24_21_groupi_n_471);
  or csa_tree_add_24_21_groupi_g6889(csa_tree_add_24_21_groupi_n_666 ,csa_tree_add_24_21_groupi_n_269 ,csa_tree_add_24_21_groupi_n_460);
  or csa_tree_add_24_21_groupi_g6890(csa_tree_add_24_21_groupi_n_665 ,csa_tree_add_24_21_groupi_n_266 ,csa_tree_add_24_21_groupi_n_410);
  or csa_tree_add_24_21_groupi_g6891(csa_tree_add_24_21_groupi_n_664 ,csa_tree_add_24_21_groupi_n_266 ,csa_tree_add_24_21_groupi_n_416);
  or csa_tree_add_24_21_groupi_g6892(csa_tree_add_24_21_groupi_n_663 ,csa_tree_add_24_21_groupi_n_260 ,csa_tree_add_24_21_groupi_n_502);
  or csa_tree_add_24_21_groupi_g6893(csa_tree_add_24_21_groupi_n_662 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_414);
  or csa_tree_add_24_21_groupi_g6894(csa_tree_add_24_21_groupi_n_661 ,csa_tree_add_24_21_groupi_n_263 ,csa_tree_add_24_21_groupi_n_441);
  or csa_tree_add_24_21_groupi_g6895(csa_tree_add_24_21_groupi_n_660 ,csa_tree_add_24_21_groupi_n_263 ,csa_tree_add_24_21_groupi_n_530);
  or csa_tree_add_24_21_groupi_g6896(csa_tree_add_24_21_groupi_n_659 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_487);
  or csa_tree_add_24_21_groupi_g6897(csa_tree_add_24_21_groupi_n_658 ,csa_tree_add_24_21_groupi_n_266 ,csa_tree_add_24_21_groupi_n_425);
  or csa_tree_add_24_21_groupi_g6898(csa_tree_add_24_21_groupi_n_657 ,csa_tree_add_24_21_groupi_n_260 ,csa_tree_add_24_21_groupi_n_525);
  or csa_tree_add_24_21_groupi_g6899(csa_tree_add_24_21_groupi_n_656 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_422);
  or csa_tree_add_24_21_groupi_g6900(csa_tree_add_24_21_groupi_n_655 ,csa_tree_add_24_21_groupi_n_269 ,csa_tree_add_24_21_groupi_n_508);
  or csa_tree_add_24_21_groupi_g6901(csa_tree_add_24_21_groupi_n_654 ,csa_tree_add_24_21_groupi_n_272 ,csa_tree_add_24_21_groupi_n_518);
  or csa_tree_add_24_21_groupi_g6902(csa_tree_add_24_21_groupi_n_653 ,csa_tree_add_24_21_groupi_n_272 ,csa_tree_add_24_21_groupi_n_506);
  or csa_tree_add_24_21_groupi_g6903(csa_tree_add_24_21_groupi_n_652 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_494);
  or csa_tree_add_24_21_groupi_g6904(csa_tree_add_24_21_groupi_n_651 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_456);
  or csa_tree_add_24_21_groupi_g6905(csa_tree_add_24_21_groupi_n_650 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_411);
  or csa_tree_add_24_21_groupi_g6906(csa_tree_add_24_21_groupi_n_649 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_510);
  or csa_tree_add_24_21_groupi_g6907(csa_tree_add_24_21_groupi_n_648 ,csa_tree_add_24_21_groupi_n_260 ,csa_tree_add_24_21_groupi_n_444);
  or csa_tree_add_24_21_groupi_g6908(csa_tree_add_24_21_groupi_n_647 ,csa_tree_add_24_21_groupi_n_272 ,csa_tree_add_24_21_groupi_n_483);
  or csa_tree_add_24_21_groupi_g6909(csa_tree_add_24_21_groupi_n_646 ,csa_tree_add_24_21_groupi_n_263 ,csa_tree_add_24_21_groupi_n_459);
  or csa_tree_add_24_21_groupi_g6910(csa_tree_add_24_21_groupi_n_645 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_509);
  or csa_tree_add_24_21_groupi_g6911(csa_tree_add_24_21_groupi_n_644 ,csa_tree_add_24_21_groupi_n_266 ,csa_tree_add_24_21_groupi_n_420);
  or csa_tree_add_24_21_groupi_g6912(csa_tree_add_24_21_groupi_n_643 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_516);
  or csa_tree_add_24_21_groupi_g6913(csa_tree_add_24_21_groupi_n_642 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_449);
  or csa_tree_add_24_21_groupi_g6914(csa_tree_add_24_21_groupi_n_641 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_419);
  or csa_tree_add_24_21_groupi_g6915(csa_tree_add_24_21_groupi_n_640 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_498);
  or csa_tree_add_24_21_groupi_g6916(csa_tree_add_24_21_groupi_n_639 ,csa_tree_add_24_21_groupi_n_272 ,csa_tree_add_24_21_groupi_n_524);
  or csa_tree_add_24_21_groupi_g6917(csa_tree_add_24_21_groupi_n_638 ,csa_tree_add_24_21_groupi_n_367 ,csa_tree_add_24_21_groupi_n_472);
  or csa_tree_add_24_21_groupi_g6918(csa_tree_add_24_21_groupi_n_637 ,csa_tree_add_24_21_groupi_n_260 ,csa_tree_add_24_21_groupi_n_500);
  or csa_tree_add_24_21_groupi_g6919(csa_tree_add_24_21_groupi_n_636 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_454);
  or csa_tree_add_24_21_groupi_g6920(csa_tree_add_24_21_groupi_n_635 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_409);
  or csa_tree_add_24_21_groupi_g6921(csa_tree_add_24_21_groupi_n_634 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_489);
  or csa_tree_add_24_21_groupi_g6922(csa_tree_add_24_21_groupi_n_633 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_408);
  or csa_tree_add_24_21_groupi_g6923(csa_tree_add_24_21_groupi_n_632 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_515);
  or csa_tree_add_24_21_groupi_g6924(csa_tree_add_24_21_groupi_n_631 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_433);
  or csa_tree_add_24_21_groupi_g6925(csa_tree_add_24_21_groupi_n_630 ,csa_tree_add_24_21_groupi_n_384 ,csa_tree_add_24_21_groupi_n_473);
  or csa_tree_add_24_21_groupi_g6926(csa_tree_add_24_21_groupi_n_629 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_527);
  or csa_tree_add_24_21_groupi_g6927(csa_tree_add_24_21_groupi_n_628 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_452);
  or csa_tree_add_24_21_groupi_g6928(csa_tree_add_24_21_groupi_n_627 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_511);
  or csa_tree_add_24_21_groupi_g6929(csa_tree_add_24_21_groupi_n_626 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_503);
  or csa_tree_add_24_21_groupi_g6930(csa_tree_add_24_21_groupi_n_625 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_521);
  or csa_tree_add_24_21_groupi_g6931(csa_tree_add_24_21_groupi_n_624 ,csa_tree_add_24_21_groupi_n_263 ,csa_tree_add_24_21_groupi_n_512);
  or csa_tree_add_24_21_groupi_g6932(csa_tree_add_24_21_groupi_n_623 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_412);
  or csa_tree_add_24_21_groupi_g6933(csa_tree_add_24_21_groupi_n_622 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_450);
  or csa_tree_add_24_21_groupi_g6934(csa_tree_add_24_21_groupi_n_621 ,csa_tree_add_24_21_groupi_n_269 ,csa_tree_add_24_21_groupi_n_486);
  or csa_tree_add_24_21_groupi_g6935(csa_tree_add_24_21_groupi_n_620 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_520);
  or csa_tree_add_24_21_groupi_g6936(csa_tree_add_24_21_groupi_n_619 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_407);
  or csa_tree_add_24_21_groupi_g6937(csa_tree_add_24_21_groupi_n_618 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_496);
  or csa_tree_add_24_21_groupi_g6938(csa_tree_add_24_21_groupi_n_617 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_529);
  or csa_tree_add_24_21_groupi_g6939(csa_tree_add_24_21_groupi_n_616 ,csa_tree_add_24_21_groupi_n_380 ,csa_tree_add_24_21_groupi_n_470);
  or csa_tree_add_24_21_groupi_g6940(csa_tree_add_24_21_groupi_n_688 ,csa_tree_add_24_21_groupi_n_337 ,csa_tree_add_24_21_groupi_n_482);
  or csa_tree_add_24_21_groupi_g6941(csa_tree_add_24_21_groupi_n_686 ,in1[0] ,csa_tree_add_24_21_groupi_n_468);
  not csa_tree_add_24_21_groupi_g6942(csa_tree_add_24_21_groupi_n_615 ,csa_tree_add_24_21_groupi_n_614);
  not csa_tree_add_24_21_groupi_g6943(csa_tree_add_24_21_groupi_n_613 ,csa_tree_add_24_21_groupi_n_612);
  not csa_tree_add_24_21_groupi_g6944(csa_tree_add_24_21_groupi_n_611 ,csa_tree_add_24_21_groupi_n_610);
  not csa_tree_add_24_21_groupi_g6945(csa_tree_add_24_21_groupi_n_609 ,csa_tree_add_24_21_groupi_n_608);
  not csa_tree_add_24_21_groupi_g6946(csa_tree_add_24_21_groupi_n_607 ,csa_tree_add_24_21_groupi_n_606);
  not csa_tree_add_24_21_groupi_g6947(csa_tree_add_24_21_groupi_n_605 ,csa_tree_add_24_21_groupi_n_604);
  not csa_tree_add_24_21_groupi_g6948(csa_tree_add_24_21_groupi_n_603 ,csa_tree_add_24_21_groupi_n_602);
  not csa_tree_add_24_21_groupi_g6949(csa_tree_add_24_21_groupi_n_601 ,csa_tree_add_24_21_groupi_n_600);
  not csa_tree_add_24_21_groupi_g6950(csa_tree_add_24_21_groupi_n_599 ,csa_tree_add_24_21_groupi_n_598);
  not csa_tree_add_24_21_groupi_g6951(csa_tree_add_24_21_groupi_n_597 ,csa_tree_add_24_21_groupi_n_596);
  not csa_tree_add_24_21_groupi_g6952(csa_tree_add_24_21_groupi_n_595 ,csa_tree_add_24_21_groupi_n_594);
  not csa_tree_add_24_21_groupi_g6953(csa_tree_add_24_21_groupi_n_593 ,csa_tree_add_24_21_groupi_n_592);
  and csa_tree_add_24_21_groupi_g6957(csa_tree_add_24_21_groupi_n_585 ,csa_tree_add_24_21_groupi_n_461 ,csa_tree_add_24_21_groupi_n_481);
  or csa_tree_add_24_21_groupi_g6958(csa_tree_add_24_21_groupi_n_584 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_447);
  or csa_tree_add_24_21_groupi_g6959(csa_tree_add_24_21_groupi_n_583 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_424);
  or csa_tree_add_24_21_groupi_g6960(csa_tree_add_24_21_groupi_n_582 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_491);
  or csa_tree_add_24_21_groupi_g6961(csa_tree_add_24_21_groupi_n_581 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_519);
  or csa_tree_add_24_21_groupi_g6962(csa_tree_add_24_21_groupi_n_580 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_417);
  or csa_tree_add_24_21_groupi_g6963(csa_tree_add_24_21_groupi_n_579 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_413);
  or csa_tree_add_24_21_groupi_g6964(csa_tree_add_24_21_groupi_n_578 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_493);
  or csa_tree_add_24_21_groupi_g6965(csa_tree_add_24_21_groupi_n_577 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_499);
  or csa_tree_add_24_21_groupi_g6966(csa_tree_add_24_21_groupi_n_576 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_514);
  or csa_tree_add_24_21_groupi_g6967(csa_tree_add_24_21_groupi_n_575 ,csa_tree_add_24_21_groupi_n_382 ,csa_tree_add_24_21_groupi_n_469);
  or csa_tree_add_24_21_groupi_g6968(csa_tree_add_24_21_groupi_n_574 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_453);
  or csa_tree_add_24_21_groupi_g6969(csa_tree_add_24_21_groupi_n_573 ,csa_tree_add_24_21_groupi_n_266 ,csa_tree_add_24_21_groupi_n_418);
  or csa_tree_add_24_21_groupi_g6970(csa_tree_add_24_21_groupi_n_572 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_522);
  or csa_tree_add_24_21_groupi_g6971(csa_tree_add_24_21_groupi_n_571 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_497);
  or csa_tree_add_24_21_groupi_g6972(csa_tree_add_24_21_groupi_n_570 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_492);
  or csa_tree_add_24_21_groupi_g6973(csa_tree_add_24_21_groupi_n_569 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_507);
  or csa_tree_add_24_21_groupi_g6974(csa_tree_add_24_21_groupi_n_568 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_526);
  or csa_tree_add_24_21_groupi_g6975(csa_tree_add_24_21_groupi_n_567 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_505);
  or csa_tree_add_24_21_groupi_g6976(csa_tree_add_24_21_groupi_n_566 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_490);
  or csa_tree_add_24_21_groupi_g6977(csa_tree_add_24_21_groupi_n_565 ,csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_423);
  or csa_tree_add_24_21_groupi_g6978(csa_tree_add_24_21_groupi_n_564 ,csa_tree_add_24_21_groupi_n_260 ,csa_tree_add_24_21_groupi_n_504);
  or csa_tree_add_24_21_groupi_g6979(csa_tree_add_24_21_groupi_n_563 ,csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_523);
  or csa_tree_add_24_21_groupi_g6980(csa_tree_add_24_21_groupi_n_562 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_495);
  or csa_tree_add_24_21_groupi_g6981(csa_tree_add_24_21_groupi_n_561 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_488);
  or csa_tree_add_24_21_groupi_g6982(csa_tree_add_24_21_groupi_n_560 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_448);
  or csa_tree_add_24_21_groupi_g6983(csa_tree_add_24_21_groupi_n_559 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_528);
  or csa_tree_add_24_21_groupi_g6984(csa_tree_add_24_21_groupi_n_558 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_445);
  or csa_tree_add_24_21_groupi_g6985(csa_tree_add_24_21_groupi_n_557 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_485);
  or csa_tree_add_24_21_groupi_g6986(csa_tree_add_24_21_groupi_n_556 ,csa_tree_add_24_21_groupi_n_263 ,csa_tree_add_24_21_groupi_n_513);
  or csa_tree_add_24_21_groupi_g6987(csa_tree_add_24_21_groupi_n_555 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_457);
  or csa_tree_add_24_21_groupi_g6988(csa_tree_add_24_21_groupi_n_554 ,csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_415);
  or csa_tree_add_24_21_groupi_g6989(csa_tree_add_24_21_groupi_n_553 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_455);
  or csa_tree_add_24_21_groupi_g6990(csa_tree_add_24_21_groupi_n_552 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_484);
  or csa_tree_add_24_21_groupi_g6991(csa_tree_add_24_21_groupi_n_551 ,csa_tree_add_24_21_groupi_n_269 ,csa_tree_add_24_21_groupi_n_458);
  or csa_tree_add_24_21_groupi_g6992(csa_tree_add_24_21_groupi_n_550 ,csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_451);
  or csa_tree_add_24_21_groupi_g6993(csa_tree_add_24_21_groupi_n_549 ,csa_tree_add_24_21_groupi_n_272 ,csa_tree_add_24_21_groupi_n_501);
  or csa_tree_add_24_21_groupi_g6994(csa_tree_add_24_21_groupi_n_548 ,csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_517);
  or csa_tree_add_24_21_groupi_g6995(csa_tree_add_24_21_groupi_n_547 ,csa_tree_add_24_21_groupi_n_54 ,csa_tree_add_24_21_groupi_n_442);
  or csa_tree_add_24_21_groupi_g6996(csa_tree_add_24_21_groupi_n_546 ,csa_tree_add_22_22_n_86 ,csa_tree_add_24_21_groupi_n_435);
  or csa_tree_add_24_21_groupi_g6997(csa_tree_add_24_21_groupi_n_545 ,csa_tree_add_22_22_n_86 ,csa_tree_add_24_21_groupi_n_439);
  or csa_tree_add_24_21_groupi_g6998(csa_tree_add_24_21_groupi_n_544 ,csa_tree_add_24_21_groupi_n_54 ,csa_tree_add_24_21_groupi_n_421);
  or csa_tree_add_24_21_groupi_g6999(csa_tree_add_24_21_groupi_n_543 ,csa_tree_add_22_22_n_86 ,csa_tree_add_24_21_groupi_n_426);
  or csa_tree_add_24_21_groupi_g7000(csa_tree_add_24_21_groupi_n_542 ,csa_tree_add_24_21_groupi_n_54 ,csa_tree_add_24_21_groupi_n_431);
  or csa_tree_add_24_21_groupi_g7001(csa_tree_add_24_21_groupi_n_541 ,csa_tree_add_22_22_n_86 ,csa_tree_add_24_21_groupi_n_440);
  or csa_tree_add_24_21_groupi_g7002(csa_tree_add_24_21_groupi_n_540 ,csa_tree_add_24_21_groupi_n_54 ,csa_tree_add_24_21_groupi_n_438);
  or csa_tree_add_24_21_groupi_g7003(csa_tree_add_24_21_groupi_n_539 ,csa_tree_add_24_21_groupi_n_54 ,csa_tree_add_24_21_groupi_n_437);
  or csa_tree_add_24_21_groupi_g7004(csa_tree_add_24_21_groupi_n_538 ,csa_tree_add_24_21_groupi_n_54 ,csa_tree_add_24_21_groupi_n_434);
  or csa_tree_add_24_21_groupi_g7005(csa_tree_add_24_21_groupi_n_537 ,csa_tree_add_22_22_n_86 ,csa_tree_add_24_21_groupi_n_432);
  or csa_tree_add_24_21_groupi_g7006(csa_tree_add_24_21_groupi_n_536 ,csa_tree_add_24_21_groupi_n_54 ,csa_tree_add_24_21_groupi_n_427);
  or csa_tree_add_24_21_groupi_g7007(csa_tree_add_24_21_groupi_n_535 ,csa_tree_add_22_22_n_86 ,csa_tree_add_24_21_groupi_n_430);
  or csa_tree_add_24_21_groupi_g7008(csa_tree_add_24_21_groupi_n_534 ,csa_tree_add_24_21_groupi_n_54 ,csa_tree_add_24_21_groupi_n_436);
  or csa_tree_add_24_21_groupi_g7009(csa_tree_add_24_21_groupi_n_533 ,csa_tree_add_22_22_n_86 ,csa_tree_add_24_21_groupi_n_429);
  or csa_tree_add_24_21_groupi_g7010(csa_tree_add_24_21_groupi_n_532 ,csa_tree_add_24_21_groupi_n_54 ,csa_tree_add_24_21_groupi_n_443);
  or csa_tree_add_24_21_groupi_g7011(csa_tree_add_24_21_groupi_n_531 ,csa_tree_add_24_21_groupi_n_54 ,csa_tree_add_24_21_groupi_n_428);
  and csa_tree_add_24_21_groupi_g7012(csa_tree_add_24_21_groupi_n_614 ,in1[11] ,csa_tree_add_24_21_groupi_n_264);
  and csa_tree_add_24_21_groupi_g7013(csa_tree_add_24_21_groupi_n_612 ,in1[9] ,csa_tree_add_24_21_groupi_n_270);
  and csa_tree_add_24_21_groupi_g7014(csa_tree_add_24_21_groupi_n_610 ,in1[7] ,csa_tree_add_24_21_groupi_n_261);
  and csa_tree_add_24_21_groupi_g7015(csa_tree_add_24_21_groupi_n_608 ,in1[5] ,csa_tree_add_24_21_groupi_n_258);
  and csa_tree_add_24_21_groupi_g7016(csa_tree_add_24_21_groupi_n_606 ,in1[3] ,csa_tree_add_24_21_groupi_n_267);
  and csa_tree_add_24_21_groupi_g7017(csa_tree_add_24_21_groupi_n_604 ,in2[0] ,csa_tree_add_24_21_groupi_n_258);
  and csa_tree_add_24_21_groupi_g7018(csa_tree_add_24_21_groupi_n_602 ,in2[0] ,csa_tree_add_24_21_groupi_n_270);
  and csa_tree_add_24_21_groupi_g7019(csa_tree_add_24_21_groupi_n_600 ,in2[0] ,csa_tree_add_24_21_groupi_n_261);
  and csa_tree_add_24_21_groupi_g7020(csa_tree_add_24_21_groupi_n_598 ,in2[0] ,csa_tree_add_24_21_groupi_n_293);
  and csa_tree_add_24_21_groupi_g7021(csa_tree_add_24_21_groupi_n_596 ,in2[0] ,csa_tree_add_24_21_groupi_n_264);
  and csa_tree_add_24_21_groupi_g7022(csa_tree_add_24_21_groupi_n_594 ,in2[0] ,csa_tree_add_24_21_groupi_n_267);
  or csa_tree_add_24_21_groupi_g7023(csa_tree_add_24_21_groupi_n_592 ,csa_tree_add_22_22_n_117 ,csa_tree_add_24_21_groupi_n_404);
  or csa_tree_add_24_21_groupi_g7024(csa_tree_add_24_21_groupi_n_590 ,csa_tree_add_24_21_groupi_n_474 ,csa_tree_add_24_21_groupi_n_267);
  or csa_tree_add_24_21_groupi_g7025(csa_tree_add_24_21_groupi_n_589 ,csa_tree_add_24_21_groupi_n_462 ,csa_tree_add_24_21_groupi_n_258);
  or csa_tree_add_24_21_groupi_g7026(csa_tree_add_24_21_groupi_n_588 ,csa_tree_add_24_21_groupi_n_467 ,csa_tree_add_24_21_groupi_n_270);
  or csa_tree_add_24_21_groupi_g7027(csa_tree_add_24_21_groupi_n_587 ,csa_tree_add_24_21_groupi_n_396 ,csa_tree_add_24_21_groupi_n_264);
  or csa_tree_add_24_21_groupi_g7028(csa_tree_add_24_21_groupi_n_586 ,csa_tree_add_24_21_groupi_n_463 ,csa_tree_add_24_21_groupi_n_261);
  xnor csa_tree_add_24_21_groupi_g7039(csa_tree_add_24_21_groupi_n_474 ,in1[3] ,in1[2]);
  and csa_tree_add_24_21_groupi_g7040(csa_tree_add_24_21_groupi_n_473 ,csa_tree_add_24_21_groupi_n_173 ,csa_tree_add_24_21_groupi_n_369);
  and csa_tree_add_24_21_groupi_g7041(csa_tree_add_24_21_groupi_n_472 ,csa_tree_add_24_21_groupi_n_173 ,csa_tree_add_24_21_groupi_n_372);
  and csa_tree_add_24_21_groupi_g7042(csa_tree_add_24_21_groupi_n_471 ,csa_tree_add_24_21_groupi_n_173 ,csa_tree_add_24_21_groupi_n_371);
  and csa_tree_add_24_21_groupi_g7043(csa_tree_add_24_21_groupi_n_470 ,csa_tree_add_24_21_groupi_n_173 ,csa_tree_add_24_21_groupi_n_364);
  and csa_tree_add_24_21_groupi_g7044(csa_tree_add_24_21_groupi_n_469 ,csa_tree_add_24_21_groupi_n_173 ,csa_tree_add_24_21_groupi_n_365);
  xnor csa_tree_add_24_21_groupi_g7046(csa_tree_add_24_21_groupi_n_467 ,in1[9] ,in1[8]);
  xnor csa_tree_add_24_21_groupi_g7047(csa_tree_add_24_21_groupi_n_466 ,in1[5] ,in2[0]);
  xnor csa_tree_add_24_21_groupi_g7048(csa_tree_add_24_21_groupi_n_465 ,in1[3] ,in2[0]);
  xnor csa_tree_add_24_21_groupi_g7049(csa_tree_add_24_21_groupi_n_464 ,in1[7] ,in2[0]);
  xnor csa_tree_add_24_21_groupi_g7050(csa_tree_add_24_21_groupi_n_463 ,in1[7] ,in1[6]);
  xnor csa_tree_add_24_21_groupi_g7051(csa_tree_add_24_21_groupi_n_462 ,in1[5] ,in1[4]);
  or csa_tree_add_24_21_groupi_g7052(csa_tree_add_24_21_groupi_n_461 ,in3[0] ,csa_tree_add_24_21_groupi_n_387);
  xnor csa_tree_add_24_21_groupi_g7053(csa_tree_add_24_21_groupi_n_530 ,in1[7] ,in2[1]);
  xnor csa_tree_add_24_21_groupi_g7054(csa_tree_add_24_21_groupi_n_529 ,in1[9] ,in2[17]);
  xnor csa_tree_add_24_21_groupi_g7055(csa_tree_add_24_21_groupi_n_528 ,in1[3] ,in2[11]);
  xnor csa_tree_add_24_21_groupi_g7056(csa_tree_add_24_21_groupi_n_527 ,in1[5] ,in2[10]);
  xnor csa_tree_add_24_21_groupi_g7057(csa_tree_add_24_21_groupi_n_526 ,in1[5] ,in2[16]);
  xnor csa_tree_add_24_21_groupi_g7058(csa_tree_add_24_21_groupi_n_525 ,in1[5] ,in2[5]);
  xnor csa_tree_add_24_21_groupi_g7059(csa_tree_add_24_21_groupi_n_524 ,in1[9] ,in2[7]);
  xnor csa_tree_add_24_21_groupi_g7060(csa_tree_add_24_21_groupi_n_523 ,in1[5] ,in2[2]);
  xnor csa_tree_add_24_21_groupi_g7061(csa_tree_add_24_21_groupi_n_522 ,in1[7] ,in2[9]);
  xnor csa_tree_add_24_21_groupi_g7062(csa_tree_add_24_21_groupi_n_521 ,in1[5] ,in2[12]);
  xnor csa_tree_add_24_21_groupi_g7063(csa_tree_add_24_21_groupi_n_520 ,in1[9] ,in2[11]);
  xnor csa_tree_add_24_21_groupi_g7064(csa_tree_add_24_21_groupi_n_519 ,in1[7] ,in2[7]);
  xnor csa_tree_add_24_21_groupi_g7065(csa_tree_add_24_21_groupi_n_518 ,in1[9] ,in2[8]);
  xnor csa_tree_add_24_21_groupi_g7066(csa_tree_add_24_21_groupi_n_517 ,in1[9] ,in2[6]);
  xnor csa_tree_add_24_21_groupi_g7067(csa_tree_add_24_21_groupi_n_516 ,in1[9] ,in2[15]);
  xnor csa_tree_add_24_21_groupi_g7068(csa_tree_add_24_21_groupi_n_515 ,in1[5] ,in2[8]);
  xnor csa_tree_add_24_21_groupi_g7069(csa_tree_add_24_21_groupi_n_514 ,in1[7] ,in2[16]);
  xnor csa_tree_add_24_21_groupi_g7070(csa_tree_add_24_21_groupi_n_513 ,in1[7] ,in2[13]);
  xnor csa_tree_add_24_21_groupi_g7071(csa_tree_add_24_21_groupi_n_512 ,in1[7] ,in2[6]);
  xnor csa_tree_add_24_21_groupi_g7072(csa_tree_add_24_21_groupi_n_511 ,in1[7] ,in2[11]);
  xnor csa_tree_add_24_21_groupi_g7073(csa_tree_add_24_21_groupi_n_510 ,in1[9] ,in2[14]);
  xnor csa_tree_add_24_21_groupi_g7074(csa_tree_add_24_21_groupi_n_509 ,in1[9] ,in2[13]);
  xnor csa_tree_add_24_21_groupi_g7075(csa_tree_add_24_21_groupi_n_508 ,in1[3] ,in2[2]);
  xnor csa_tree_add_24_21_groupi_g7076(csa_tree_add_24_21_groupi_n_507 ,in1[5] ,in2[4]);
  xnor csa_tree_add_24_21_groupi_g7077(csa_tree_add_24_21_groupi_n_506 ,in1[9] ,in2[12]);
  xnor csa_tree_add_24_21_groupi_g7078(csa_tree_add_24_21_groupi_n_505 ,in1[7] ,in2[12]);
  xnor csa_tree_add_24_21_groupi_g7079(csa_tree_add_24_21_groupi_n_504 ,in1[5] ,in2[11]);
  xnor csa_tree_add_24_21_groupi_g7080(csa_tree_add_24_21_groupi_n_503 ,in1[9] ,in2[3]);
  xnor csa_tree_add_24_21_groupi_g7081(csa_tree_add_24_21_groupi_n_502 ,in1[5] ,in2[17]);
  xnor csa_tree_add_24_21_groupi_g7082(csa_tree_add_24_21_groupi_n_501 ,in1[9] ,in2[5]);
  xnor csa_tree_add_24_21_groupi_g7083(csa_tree_add_24_21_groupi_n_500 ,in1[5] ,in2[14]);
  xnor csa_tree_add_24_21_groupi_g7084(csa_tree_add_24_21_groupi_n_499 ,in1[3] ,in2[16]);
  xnor csa_tree_add_24_21_groupi_g7085(csa_tree_add_24_21_groupi_n_498 ,in1[5] ,in2[15]);
  xnor csa_tree_add_24_21_groupi_g7086(csa_tree_add_24_21_groupi_n_497 ,in1[7] ,in2[15]);
  xnor csa_tree_add_24_21_groupi_g7087(csa_tree_add_24_21_groupi_n_496 ,in1[7] ,in2[5]);
  xnor csa_tree_add_24_21_groupi_g7088(csa_tree_add_24_21_groupi_n_495 ,in1[3] ,in2[1]);
  xnor csa_tree_add_24_21_groupi_g7089(csa_tree_add_24_21_groupi_n_494 ,in1[5] ,in2[3]);
  xnor csa_tree_add_24_21_groupi_g7090(csa_tree_add_24_21_groupi_n_493 ,in1[7] ,in2[4]);
  xnor csa_tree_add_24_21_groupi_g7091(csa_tree_add_24_21_groupi_n_492 ,in1[3] ,in2[8]);
  xnor csa_tree_add_24_21_groupi_g7092(csa_tree_add_24_21_groupi_n_491 ,in1[5] ,in2[7]);
  xnor csa_tree_add_24_21_groupi_g7093(csa_tree_add_24_21_groupi_n_490 ,in1[5] ,in2[6]);
  xnor csa_tree_add_24_21_groupi_g7094(csa_tree_add_24_21_groupi_n_489 ,in1[3] ,in2[17]);
  xnor csa_tree_add_24_21_groupi_g7095(csa_tree_add_24_21_groupi_n_488 ,in1[3] ,in2[6]);
  xnor csa_tree_add_24_21_groupi_g7096(csa_tree_add_24_21_groupi_n_487 ,in1[3] ,in2[13]);
  xnor csa_tree_add_24_21_groupi_g7097(csa_tree_add_24_21_groupi_n_486 ,in1[3] ,in2[14]);
  xnor csa_tree_add_24_21_groupi_g7098(csa_tree_add_24_21_groupi_n_485 ,in1[9] ,in2[1]);
  xnor csa_tree_add_24_21_groupi_g7099(csa_tree_add_24_21_groupi_n_484 ,in1[3] ,in2[5]);
  xnor csa_tree_add_24_21_groupi_g7100(csa_tree_add_24_21_groupi_n_483 ,in1[9] ,in2[16]);
  or csa_tree_add_24_21_groupi_g7101(csa_tree_add_24_21_groupi_n_482 ,csa_tree_add_22_22_n_82 ,csa_tree_add_24_21_groupi_n_387);
  or csa_tree_add_24_21_groupi_g7102(csa_tree_add_24_21_groupi_n_481 ,csa_tree_add_24_21_groupi_n_342 ,csa_tree_add_24_21_groupi_n_386);
  xnor csa_tree_add_24_21_groupi_g7103(csa_tree_add_24_21_groupi_n_479 ,csa_tree_add_22_22_n_114 ,in1[6]);
  xnor csa_tree_add_24_21_groupi_g7104(csa_tree_add_24_21_groupi_n_477 ,csa_tree_add_22_22_n_102 ,in1[4]);
  xnor csa_tree_add_24_21_groupi_g7105(csa_tree_add_24_21_groupi_n_475 ,csa_tree_add_22_22_n_100 ,in1[8]);
  not csa_tree_add_24_21_groupi_g7106(csa_tree_add_24_21_groupi_n_406 ,csa_tree_add_24_21_groupi_n_405);
  not csa_tree_add_24_21_groupi_g7107(csa_tree_add_24_21_groupi_n_404 ,csa_tree_add_24_21_groupi_n_200);
  xnor csa_tree_add_24_21_groupi_g7117(csa_tree_add_24_21_groupi_n_396 ,in1[11] ,in1[10]);
  xnor csa_tree_add_24_21_groupi_g7119(csa_tree_add_24_21_groupi_n_394 ,in1[9] ,in2[0]);
  xnor csa_tree_add_24_21_groupi_g7120(csa_tree_add_24_21_groupi_n_393 ,in1[11] ,in2[0]);
  xnor csa_tree_add_24_21_groupi_g7121(csa_tree_add_24_21_groupi_n_460 ,in1[3] ,in2[7]);
  xnor csa_tree_add_24_21_groupi_g7122(csa_tree_add_24_21_groupi_n_459 ,in1[7] ,in2[17]);
  xnor csa_tree_add_24_21_groupi_g7123(csa_tree_add_24_21_groupi_n_458 ,in1[3] ,in2[9]);
  xnor csa_tree_add_24_21_groupi_g7124(csa_tree_add_24_21_groupi_n_457 ,in1[3] ,in2[10]);
  xnor csa_tree_add_24_21_groupi_g7125(csa_tree_add_24_21_groupi_n_456 ,in1[7] ,in2[14]);
  xnor csa_tree_add_24_21_groupi_g7126(csa_tree_add_24_21_groupi_n_455 ,in1[9] ,in2[9]);
  xnor csa_tree_add_24_21_groupi_g7127(csa_tree_add_24_21_groupi_n_454 ,in1[7] ,in2[8]);
  xnor csa_tree_add_24_21_groupi_g7128(csa_tree_add_24_21_groupi_n_453 ,in1[9] ,in2[10]);
  xnor csa_tree_add_24_21_groupi_g7129(csa_tree_add_24_21_groupi_n_452 ,in1[9] ,in2[2]);
  xnor csa_tree_add_24_21_groupi_g7130(csa_tree_add_24_21_groupi_n_451 ,in1[3] ,in2[4]);
  xnor csa_tree_add_24_21_groupi_g7131(csa_tree_add_24_21_groupi_n_450 ,in1[3] ,in2[3]);
  xnor csa_tree_add_24_21_groupi_g7132(csa_tree_add_24_21_groupi_n_449 ,in1[5] ,in2[9]);
  xnor csa_tree_add_24_21_groupi_g7133(csa_tree_add_24_21_groupi_n_448 ,in1[3] ,in2[15]);
  xnor csa_tree_add_24_21_groupi_g7134(csa_tree_add_24_21_groupi_n_447 ,in1[7] ,in2[2]);
  xnor csa_tree_add_24_21_groupi_g7135(csa_tree_add_24_21_groupi_n_446 ,in1[3] ,in2[12]);
  xnor csa_tree_add_24_21_groupi_g7136(csa_tree_add_24_21_groupi_n_445 ,in1[9] ,in2[4]);
  xnor csa_tree_add_24_21_groupi_g7137(csa_tree_add_24_21_groupi_n_444 ,in1[5] ,in2[1]);
  xnor csa_tree_add_24_21_groupi_g7138(csa_tree_add_24_21_groupi_n_392 ,in3[29] ,in3[28]);
  xnor csa_tree_add_24_21_groupi_g7139(csa_tree_add_24_21_groupi_n_443 ,in1[1] ,in2[8]);
  xnor csa_tree_add_24_21_groupi_g7140(csa_tree_add_24_21_groupi_n_442 ,in1[1] ,in2[16]);
  xnor csa_tree_add_24_21_groupi_g7141(csa_tree_add_24_21_groupi_n_441 ,in1[7] ,in2[3]);
  xnor csa_tree_add_24_21_groupi_g7142(csa_tree_add_24_21_groupi_n_440 ,in1[1] ,in2[1]);
  xnor csa_tree_add_24_21_groupi_g7143(csa_tree_add_24_21_groupi_n_439 ,in1[1] ,in2[2]);
  xnor csa_tree_add_24_21_groupi_g7144(csa_tree_add_24_21_groupi_n_391 ,in3[23] ,in3[22]);
  xnor csa_tree_add_24_21_groupi_g7145(csa_tree_add_24_21_groupi_n_438 ,in1[1] ,in2[13]);
  xnor csa_tree_add_24_21_groupi_g7146(csa_tree_add_24_21_groupi_n_437 ,in1[1] ,in2[17]);
  xnor csa_tree_add_24_21_groupi_g7147(csa_tree_add_24_21_groupi_n_436 ,in1[1] ,in2[10]);
  xnor csa_tree_add_24_21_groupi_g7148(csa_tree_add_24_21_groupi_n_435 ,in1[1] ,in2[4]);
  xnor csa_tree_add_24_21_groupi_g7149(csa_tree_add_24_21_groupi_n_434 ,in1[1] ,in2[12]);
  xnor csa_tree_add_24_21_groupi_g7150(csa_tree_add_24_21_groupi_n_433 ,in1[5] ,in2[13]);
  xnor csa_tree_add_24_21_groupi_g7151(csa_tree_add_24_21_groupi_n_432 ,in1[1] ,in2[14]);
  xnor csa_tree_add_24_21_groupi_g7152(csa_tree_add_24_21_groupi_n_431 ,in1[1] ,in2[11]);
  xnor csa_tree_add_24_21_groupi_g7153(csa_tree_add_24_21_groupi_n_430 ,in1[1] ,in2[3]);
  xnor csa_tree_add_24_21_groupi_g7154(csa_tree_add_24_21_groupi_n_429 ,in1[1] ,in2[9]);
  xnor csa_tree_add_24_21_groupi_g7155(csa_tree_add_24_21_groupi_n_428 ,in1[1] ,in2[6]);
  xnor csa_tree_add_24_21_groupi_g7156(csa_tree_add_24_21_groupi_n_427 ,in1[1] ,in2[5]);
  xnor csa_tree_add_24_21_groupi_g7157(csa_tree_add_24_21_groupi_n_426 ,in1[1] ,in2[7]);
  xnor csa_tree_add_24_21_groupi_g7158(csa_tree_add_24_21_groupi_n_425 ,in1[11] ,in2[11]);
  xnor csa_tree_add_24_21_groupi_g7159(csa_tree_add_24_21_groupi_n_424 ,in1[11] ,in2[6]);
  xnor csa_tree_add_24_21_groupi_g7160(csa_tree_add_24_21_groupi_n_423 ,in1[11] ,in2[13]);
  xnor csa_tree_add_24_21_groupi_g7161(csa_tree_add_24_21_groupi_n_422 ,in1[11] ,in2[17]);
  xnor csa_tree_add_24_21_groupi_g7162(csa_tree_add_24_21_groupi_n_421 ,in1[1] ,in2[15]);
  xnor csa_tree_add_24_21_groupi_g7163(csa_tree_add_24_21_groupi_n_420 ,in1[11] ,in2[12]);
  xnor csa_tree_add_24_21_groupi_g7164(csa_tree_add_24_21_groupi_n_419 ,in1[11] ,in2[4]);
  xnor csa_tree_add_24_21_groupi_g7165(csa_tree_add_24_21_groupi_n_418 ,in1[11] ,in2[2]);
  xnor csa_tree_add_24_21_groupi_g7166(csa_tree_add_24_21_groupi_n_417 ,in1[11] ,in2[3]);
  xnor csa_tree_add_24_21_groupi_g7167(csa_tree_add_24_21_groupi_n_416 ,in1[11] ,in2[15]);
  xnor csa_tree_add_24_21_groupi_g7168(csa_tree_add_24_21_groupi_n_390 ,in3[27] ,in3[26]);
  xnor csa_tree_add_24_21_groupi_g7169(csa_tree_add_24_21_groupi_n_415 ,in1[7] ,in2[10]);
  xnor csa_tree_add_24_21_groupi_g7170(csa_tree_add_24_21_groupi_n_414 ,in1[11] ,in2[1]);
  xnor csa_tree_add_24_21_groupi_g7171(csa_tree_add_24_21_groupi_n_413 ,in1[11] ,in2[8]);
  xnor csa_tree_add_24_21_groupi_g7172(csa_tree_add_24_21_groupi_n_412 ,in1[11] ,in2[14]);
  xnor csa_tree_add_24_21_groupi_g7173(csa_tree_add_24_21_groupi_n_411 ,in1[11] ,in2[5]);
  xnor csa_tree_add_24_21_groupi_g7174(csa_tree_add_24_21_groupi_n_410 ,in1[11] ,in2[10]);
  xnor csa_tree_add_24_21_groupi_g7175(csa_tree_add_24_21_groupi_n_409 ,in1[11] ,in2[7]);
  xnor csa_tree_add_24_21_groupi_g7176(csa_tree_add_24_21_groupi_n_408 ,in1[11] ,in2[9]);
  xnor csa_tree_add_24_21_groupi_g7177(csa_tree_add_24_21_groupi_n_407 ,in1[11] ,in2[16]);
  xnor csa_tree_add_24_21_groupi_g7178(csa_tree_add_24_21_groupi_n_389 ,in3[21] ,in3[20]);
  xnor csa_tree_add_24_21_groupi_g7179(csa_tree_add_24_21_groupi_n_388 ,in3[25] ,in3[24]);
  xnor csa_tree_add_24_21_groupi_g7180(csa_tree_add_24_21_groupi_n_405 ,in3[31] ,in3[30]);
  xnor csa_tree_add_24_21_groupi_g7181(csa_tree_add_24_21_groupi_n_402 ,in1[12] ,in1[11]);
  xnor csa_tree_add_24_21_groupi_g7182(csa_tree_add_24_21_groupi_n_399 ,csa_tree_add_22_22_n_101 ,in1[2]);
  xnor csa_tree_add_24_21_groupi_g7183(csa_tree_add_24_21_groupi_n_397 ,csa_tree_add_22_22_n_103 ,in1[10]);
  not csa_tree_add_24_21_groupi_g7184(csa_tree_add_24_21_groupi_n_386 ,csa_tree_add_24_21_groupi_n_387);
  nor csa_tree_add_24_21_groupi_g7185(csa_tree_add_24_21_groupi_n_385 ,in3[23] ,in3[22]);
  nor csa_tree_add_24_21_groupi_g7186(csa_tree_add_24_21_groupi_n_384 ,in1[2] ,in1[1]);
  and csa_tree_add_24_21_groupi_g7187(csa_tree_add_24_21_groupi_n_383 ,in3[27] ,in3[26]);
  nor csa_tree_add_24_21_groupi_g7188(csa_tree_add_24_21_groupi_n_382 ,in1[8] ,in1[7]);
  nor csa_tree_add_24_21_groupi_g7189(csa_tree_add_24_21_groupi_n_381 ,in1[4] ,in1[3]);
  nor csa_tree_add_24_21_groupi_g7190(csa_tree_add_24_21_groupi_n_380 ,in1[10] ,in1[9]);
  or csa_tree_add_24_21_groupi_g7191(csa_tree_add_24_21_groupi_n_379 ,csa_tree_add_24_21_groupi_n_332 ,csa_tree_add_24_21_groupi_n_330);
  or csa_tree_add_24_21_groupi_g7192(csa_tree_add_24_21_groupi_n_378 ,csa_tree_add_24_21_groupi_n_331 ,csa_tree_add_24_21_groupi_n_329);
  nor csa_tree_add_24_21_groupi_g7193(csa_tree_add_24_21_groupi_n_377 ,in3[29] ,in3[28]);
  nor csa_tree_add_24_21_groupi_g7194(csa_tree_add_24_21_groupi_n_376 ,in3[31] ,in3[30]);
  and csa_tree_add_24_21_groupi_g7195(csa_tree_add_24_21_groupi_n_387 ,in1[0] ,in2[0]);
  or csa_tree_add_24_21_groupi_g7196(csa_tree_add_24_21_groupi_n_374 ,csa_tree_add_24_21_groupi_n_355 ,csa_tree_add_24_21_groupi_n_349);
  or csa_tree_add_24_21_groupi_g7197(csa_tree_add_24_21_groupi_n_373 ,csa_tree_add_24_21_groupi_n_335 ,csa_tree_add_24_21_groupi_n_328);
  or csa_tree_add_24_21_groupi_g7198(csa_tree_add_24_21_groupi_n_372 ,csa_tree_add_22_22_n_96 ,csa_tree_add_22_22_n_114);
  or csa_tree_add_24_21_groupi_g7199(csa_tree_add_24_21_groupi_n_371 ,csa_tree_add_22_22_n_97 ,csa_tree_add_22_22_n_102);
  nor csa_tree_add_24_21_groupi_g7200(csa_tree_add_24_21_groupi_n_370 ,in3[25] ,in3[24]);
  or csa_tree_add_24_21_groupi_g7201(csa_tree_add_24_21_groupi_n_369 ,csa_tree_add_22_22_n_116 ,csa_tree_add_22_22_n_82);
  or csa_tree_add_24_21_groupi_g7202(csa_tree_add_24_21_groupi_n_368 ,in3[27] ,in3[26]);
  nor csa_tree_add_24_21_groupi_g7203(csa_tree_add_24_21_groupi_n_367 ,in1[6] ,in1[5]);
  nor csa_tree_add_24_21_groupi_g7204(csa_tree_add_24_21_groupi_n_366 ,in3[21] ,in3[20]);
  or csa_tree_add_24_21_groupi_g7205(csa_tree_add_24_21_groupi_n_365 ,csa_tree_add_22_22_n_98 ,csa_tree_add_22_22_n_100);
  or csa_tree_add_24_21_groupi_g7206(csa_tree_add_24_21_groupi_n_364 ,csa_tree_add_22_22_n_115 ,csa_tree_add_22_22_n_103);
  and csa_tree_add_24_21_groupi_g7207(csa_tree_add_24_21_groupi_n_375 ,in1[1] ,in1[0]);
  not csa_tree_add_24_21_groupi_g7208(csa_tree_add_24_21_groupi_n_363 ,in3[19]);
  not csa_tree_add_24_21_groupi_g7209(csa_tree_add_24_21_groupi_n_362 ,in3[7]);
  not csa_tree_add_24_21_groupi_g7210(csa_tree_add_24_21_groupi_n_361 ,in3[5]);
  not csa_tree_add_24_21_groupi_g7211(csa_tree_add_24_21_groupi_n_360 ,in3[11]);
  not csa_tree_add_24_21_groupi_g7212(csa_tree_add_24_21_groupi_n_359 ,in3[8]);
  not csa_tree_add_24_21_groupi_g7213(csa_tree_add_24_21_groupi_n_358 ,in3[2]);
  not csa_tree_add_24_21_groupi_g7214(csa_tree_add_24_21_groupi_n_357 ,in3[6]);
  not csa_tree_add_24_21_groupi_g7215(csa_tree_add_24_21_groupi_n_356 ,in3[10]);
  not csa_tree_add_24_21_groupi_g7216(csa_tree_add_24_21_groupi_n_355 ,in3[25]);
  not csa_tree_add_24_21_groupi_g7222(csa_tree_add_24_21_groupi_n_349 ,in3[24]);
  not csa_tree_add_24_21_groupi_g7223(csa_tree_add_24_21_groupi_n_348 ,in3[26]);
  not csa_tree_add_24_21_groupi_g7224(csa_tree_add_24_21_groupi_n_347 ,in2[8]);
  not csa_tree_add_24_21_groupi_g7225(csa_tree_add_24_21_groupi_n_346 ,in2[7]);
  not csa_tree_add_24_21_groupi_g7229(csa_tree_add_24_21_groupi_n_342 ,in3[0]);
  not csa_tree_add_24_21_groupi_g7230(csa_tree_add_24_21_groupi_n_341 ,in3[18]);
  not csa_tree_add_24_21_groupi_g7231(csa_tree_add_24_21_groupi_n_340 ,in3[17]);
  not csa_tree_add_24_21_groupi_g7233(csa_tree_add_24_21_groupi_n_338 ,in3[9]);
  not csa_tree_add_24_21_groupi_g7234(csa_tree_add_24_21_groupi_n_337 ,in3[1]);
  not csa_tree_add_24_21_groupi_g7235(csa_tree_add_24_21_groupi_n_336 ,in3[3]);
  not csa_tree_add_24_21_groupi_g7236(csa_tree_add_24_21_groupi_n_335 ,in3[29]);
  not csa_tree_add_24_21_groupi_g7237(csa_tree_add_24_21_groupi_n_334 ,in3[12]);
  not csa_tree_add_24_21_groupi_g7238(csa_tree_add_24_21_groupi_n_333 ,in3[4]);
  not csa_tree_add_24_21_groupi_g7239(csa_tree_add_24_21_groupi_n_332 ,in3[23]);
  not csa_tree_add_24_21_groupi_g7240(csa_tree_add_24_21_groupi_n_331 ,in3[21]);
  not csa_tree_add_24_21_groupi_g7241(csa_tree_add_24_21_groupi_n_330 ,in3[22]);
  not csa_tree_add_24_21_groupi_g7242(csa_tree_add_24_21_groupi_n_329 ,in3[20]);
  not csa_tree_add_24_21_groupi_g7243(csa_tree_add_24_21_groupi_n_328 ,in3[28]);
  not csa_tree_add_24_21_groupi_g7244(csa_tree_add_24_21_groupi_n_327 ,in2[17]);
  not csa_tree_add_24_21_groupi_g7246(csa_tree_add_24_21_groupi_n_325 ,in2[0]);
  not csa_tree_add_24_21_groupi_drc_bufs7370(csa_tree_add_24_21_groupi_n_293 ,csa_tree_add_24_21_groupi_n_291);
  not csa_tree_add_24_21_groupi_drc_bufs7372(csa_tree_add_24_21_groupi_n_291 ,csa_tree_add_24_21_groupi_n_404);
  not csa_tree_add_24_21_groupi_drc_bufs7386(csa_tree_add_24_21_groupi_n_281 ,csa_tree_add_24_21_groupi_n_279);
  not csa_tree_add_24_21_groupi_drc_bufs7388(csa_tree_add_24_21_groupi_n_279 ,csa_tree_add_24_21_groupi_n_593);
  not csa_tree_add_24_21_groupi_drc_bufs7390(csa_tree_add_24_21_groupi_n_278 ,csa_tree_add_24_21_groupi_n_276);
  not csa_tree_add_24_21_groupi_drc_bufs7391(csa_tree_add_24_21_groupi_n_277 ,csa_tree_add_24_21_groupi_n_276);
  not csa_tree_add_24_21_groupi_drc_bufs7392(csa_tree_add_24_21_groupi_n_276 ,csa_tree_add_24_21_groupi_n_321);
  not csa_tree_add_24_21_groupi_drc_bufs7398(csa_tree_add_24_21_groupi_n_272 ,csa_tree_add_24_21_groupi_n_270);
  not csa_tree_add_24_21_groupi_drc_bufs7400(csa_tree_add_24_21_groupi_n_270 ,csa_tree_add_24_21_groupi_n_314);
  not csa_tree_add_24_21_groupi_drc_bufs7402(csa_tree_add_24_21_groupi_n_269 ,csa_tree_add_24_21_groupi_n_267);
  not csa_tree_add_24_21_groupi_drc_bufs7404(csa_tree_add_24_21_groupi_n_267 ,csa_tree_add_24_21_groupi_n_311);
  not csa_tree_add_24_21_groupi_drc_bufs7406(csa_tree_add_24_21_groupi_n_266 ,csa_tree_add_24_21_groupi_n_264);
  not csa_tree_add_24_21_groupi_drc_bufs7408(csa_tree_add_24_21_groupi_n_264 ,csa_tree_add_24_21_groupi_n_309);
  not csa_tree_add_24_21_groupi_drc_bufs7410(csa_tree_add_24_21_groupi_n_263 ,csa_tree_add_24_21_groupi_n_261);
  not csa_tree_add_24_21_groupi_drc_bufs7412(csa_tree_add_24_21_groupi_n_261 ,csa_tree_add_24_21_groupi_n_318);
  not csa_tree_add_24_21_groupi_drc_bufs7414(csa_tree_add_24_21_groupi_n_260 ,csa_tree_add_24_21_groupi_n_258);
  not csa_tree_add_24_21_groupi_drc_bufs7416(csa_tree_add_24_21_groupi_n_258 ,csa_tree_add_24_21_groupi_n_316);
  not csa_tree_add_24_21_groupi_drc_bufs7419(csa_tree_add_24_21_groupi_n_257 ,csa_tree_add_24_21_groupi_n_320);
  not csa_tree_add_24_21_groupi_drc_bufs7420(csa_tree_add_24_21_groupi_n_320 ,csa_tree_add_24_21_groupi_n_481);
  not csa_tree_add_24_21_groupi_drc_bufs7426(csa_tree_add_24_21_groupi_n_254 ,csa_tree_add_24_21_groupi_n_253);
  not csa_tree_add_24_21_groupi_drc_bufs7428(csa_tree_add_24_21_groupi_n_253 ,csa_tree_add_24_21_groupi_n_281);
  buf csa_tree_add_24_21_groupi_drc_bufs7437(out1[6] ,csa_tree_add_24_21_groupi_n_1912);
  buf csa_tree_add_24_21_groupi_drc_bufs7438(out1[1] ,csa_tree_add_24_21_groupi_n_1332);
  buf csa_tree_add_24_21_groupi_drc_bufs7439(out1[3] ,csa_tree_add_24_21_groupi_n_1710);
  buf csa_tree_add_24_21_groupi_drc_bufs7440(out1[2] ,csa_tree_add_24_21_groupi_n_1535);
  buf csa_tree_add_24_21_groupi_drc_bufs7441(out1[5] ,csa_tree_add_24_21_groupi_n_1841);
  buf csa_tree_add_24_21_groupi_drc_bufs7442(out1[4] ,csa_tree_add_24_21_groupi_n_1762);
  buf csa_tree_add_24_21_groupi_drc_bufs7443(out1[0] ,csa_tree_add_24_21_groupi_n_585);
  buf csa_tree_add_24_21_groupi_drc_bufs7444(out1[31] ,csa_tree_add_24_21_groupi_n_2026);
  buf csa_tree_add_24_21_groupi_drc_bufs7445(out1[29] ,csa_tree_add_24_21_groupi_n_2020);
  buf csa_tree_add_24_21_groupi_drc_bufs7446(out1[14] ,csa_tree_add_24_21_groupi_n_1975);
  buf csa_tree_add_24_21_groupi_drc_bufs7447(out1[17] ,csa_tree_add_24_21_groupi_n_1984);
  buf csa_tree_add_24_21_groupi_drc_bufs7448(out1[22] ,csa_tree_add_24_21_groupi_n_1999);
  buf csa_tree_add_24_21_groupi_drc_bufs7449(out1[18] ,csa_tree_add_24_21_groupi_n_1987);
  buf csa_tree_add_24_21_groupi_drc_bufs7450(out1[26] ,csa_tree_add_24_21_groupi_n_2011);
  buf csa_tree_add_24_21_groupi_drc_bufs7451(out1[7] ,csa_tree_add_24_21_groupi_n_1949);
  buf csa_tree_add_24_21_groupi_drc_bufs7452(out1[27] ,csa_tree_add_24_21_groupi_n_2014);
  buf csa_tree_add_24_21_groupi_drc_bufs7453(out1[21] ,csa_tree_add_24_21_groupi_n_1996);
  buf csa_tree_add_24_21_groupi_drc_bufs7454(out1[16] ,csa_tree_add_24_21_groupi_n_1981);
  buf csa_tree_add_24_21_groupi_drc_bufs7455(out1[19] ,csa_tree_add_24_21_groupi_n_1990);
  buf csa_tree_add_24_21_groupi_drc_bufs7456(out1[25] ,csa_tree_add_24_21_groupi_n_2008);
  buf csa_tree_add_24_21_groupi_drc_bufs7457(out1[24] ,csa_tree_add_24_21_groupi_n_2005);
  buf csa_tree_add_24_21_groupi_drc_bufs7458(out1[28] ,csa_tree_add_24_21_groupi_n_2017);
  buf csa_tree_add_24_21_groupi_drc_bufs7459(out1[30] ,csa_tree_add_24_21_groupi_n_2023);
  buf csa_tree_add_24_21_groupi_drc_bufs7460(out1[15] ,csa_tree_add_24_21_groupi_n_1978);
  buf csa_tree_add_24_21_groupi_drc_bufs7461(out1[12] ,csa_tree_add_24_21_groupi_n_1969);
  buf csa_tree_add_24_21_groupi_drc_bufs7462(out1[10] ,csa_tree_add_24_21_groupi_n_1963);
  buf csa_tree_add_24_21_groupi_drc_bufs7463(out1[11] ,csa_tree_add_24_21_groupi_n_1966);
  buf csa_tree_add_24_21_groupi_drc_bufs7464(out1[13] ,csa_tree_add_24_21_groupi_n_1972);
  buf csa_tree_add_24_21_groupi_drc_bufs7465(out1[23] ,csa_tree_add_24_21_groupi_n_2002);
  buf csa_tree_add_24_21_groupi_drc_bufs7466(out1[8] ,csa_tree_add_24_21_groupi_n_1957);
  buf csa_tree_add_24_21_groupi_drc_bufs7467(out1[20] ,csa_tree_add_24_21_groupi_n_1993);
  buf csa_tree_add_24_21_groupi_drc_bufs7468(out1[9] ,csa_tree_add_24_21_groupi_n_1960);
  not csa_tree_add_24_21_groupi_drc_bufs7499(csa_tree_add_24_21_groupi_n_220 ,csa_tree_add_24_21_groupi_n_218);
  not csa_tree_add_24_21_groupi_drc_bufs7501(csa_tree_add_24_21_groupi_n_218 ,csa_tree_add_24_21_groupi_n_587);
  not csa_tree_add_24_21_groupi_drc_bufs7504(csa_tree_add_24_21_groupi_n_217 ,csa_tree_add_24_21_groupi_n_215);
  not csa_tree_add_24_21_groupi_drc_bufs7506(csa_tree_add_24_21_groupi_n_215 ,csa_tree_add_24_21_groupi_n_586);
  not csa_tree_add_24_21_groupi_drc_bufs7509(csa_tree_add_24_21_groupi_n_214 ,csa_tree_add_24_21_groupi_n_212);
  not csa_tree_add_24_21_groupi_drc_bufs7511(csa_tree_add_24_21_groupi_n_212 ,csa_tree_add_24_21_groupi_n_686);
  not csa_tree_add_24_21_groupi_drc_bufs7514(csa_tree_add_24_21_groupi_n_211 ,csa_tree_add_24_21_groupi_n_209);
  not csa_tree_add_24_21_groupi_drc_bufs7516(csa_tree_add_24_21_groupi_n_209 ,csa_tree_add_24_21_groupi_n_590);
  not csa_tree_add_24_21_groupi_drc_bufs7519(csa_tree_add_24_21_groupi_n_208 ,csa_tree_add_24_21_groupi_n_206);
  not csa_tree_add_24_21_groupi_drc_bufs7521(csa_tree_add_24_21_groupi_n_206 ,csa_tree_add_24_21_groupi_n_589);
  not csa_tree_add_24_21_groupi_drc_bufs7524(csa_tree_add_24_21_groupi_n_205 ,csa_tree_add_24_21_groupi_n_203);
  not csa_tree_add_24_21_groupi_drc_bufs7526(csa_tree_add_24_21_groupi_n_203 ,csa_tree_add_24_21_groupi_n_588);
  not csa_tree_add_24_21_groupi_drc_bufs7539(csa_tree_add_24_21_groupi_n_200 ,csa_tree_add_24_21_groupi_n_198);
  not csa_tree_add_24_21_groupi_drc_bufs7541(csa_tree_add_24_21_groupi_n_198 ,csa_tree_add_24_21_groupi_n_402);
  not csa_tree_add_24_21_groupi_drc_bufs7573(csa_tree_add_24_21_groupi_n_321 ,csa_tree_add_24_21_groupi_n_592);
  not csa_tree_add_24_21_groupi_drc_bufs7577(csa_tree_add_24_21_groupi_n_314 ,csa_tree_add_24_21_groupi_n_475);
  not csa_tree_add_24_21_groupi_drc_bufs7581(csa_tree_add_24_21_groupi_n_311 ,csa_tree_add_24_21_groupi_n_399);
  not csa_tree_add_24_21_groupi_drc_bufs7585(csa_tree_add_24_21_groupi_n_309 ,csa_tree_add_24_21_groupi_n_397);
  not csa_tree_add_24_21_groupi_drc_bufs7589(csa_tree_add_24_21_groupi_n_318 ,csa_tree_add_24_21_groupi_n_479);
  not csa_tree_add_24_21_groupi_drc_bufs7593(csa_tree_add_24_21_groupi_n_316 ,csa_tree_add_24_21_groupi_n_477);
  not csa_tree_add_24_21_groupi_drc_bufs7596(csa_tree_add_24_21_groupi_n_173 ,csa_tree_add_24_21_groupi_n_172);
  not csa_tree_add_24_21_groupi_drc_bufs7597(csa_tree_add_24_21_groupi_n_172 ,csa_tree_add_24_21_groupi_n_325);
  not csa_tree_add_24_21_groupi_drc_bufs7619(csa_tree_add_24_21_groupi_n_166 ,csa_tree_add_24_21_groupi_n_164);
  not csa_tree_add_24_21_groupi_drc_bufs7621(csa_tree_add_24_21_groupi_n_164 ,csa_tree_add_24_21_groupi_n_272);
  not csa_tree_add_24_21_groupi_drc_bufs7627(csa_tree_add_24_21_groupi_n_160 ,csa_tree_add_24_21_groupi_n_158);
  not csa_tree_add_24_21_groupi_drc_bufs7629(csa_tree_add_24_21_groupi_n_158 ,csa_tree_add_24_21_groupi_n_269);
  not csa_tree_add_24_21_groupi_drc_bufs7635(csa_tree_add_24_21_groupi_n_154 ,csa_tree_add_24_21_groupi_n_152);
  not csa_tree_add_24_21_groupi_drc_bufs7637(csa_tree_add_24_21_groupi_n_152 ,csa_tree_add_24_21_groupi_n_266);
  not csa_tree_add_24_21_groupi_drc_bufs7639(csa_tree_add_24_21_groupi_n_151 ,csa_tree_add_24_21_groupi_n_149);
  not csa_tree_add_24_21_groupi_drc_bufs7641(csa_tree_add_24_21_groupi_n_149 ,csa_tree_add_24_21_groupi_n_263);
  not csa_tree_add_24_21_groupi_drc_bufs7643(csa_tree_add_24_21_groupi_n_148 ,csa_tree_add_24_21_groupi_n_146);
  not csa_tree_add_24_21_groupi_drc_bufs7645(csa_tree_add_24_21_groupi_n_146 ,csa_tree_add_24_21_groupi_n_260);
  not csa_tree_add_24_21_groupi_drc_bufs7687(csa_tree_add_24_21_groupi_n_120 ,csa_tree_add_24_21_groupi_n_118);
  not csa_tree_add_24_21_groupi_drc_bufs7688(csa_tree_add_24_21_groupi_n_119 ,csa_tree_add_24_21_groupi_n_118);
  not csa_tree_add_24_21_groupi_drc_bufs7689(csa_tree_add_24_21_groupi_n_118 ,csa_tree_add_24_21_groupi_n_686);
  not csa_tree_add_24_21_groupi_drc_bufs7731(csa_tree_add_24_21_groupi_n_92 ,csa_tree_add_24_21_groupi_n_90);
  not csa_tree_add_24_21_groupi_drc_bufs7732(csa_tree_add_24_21_groupi_n_91 ,csa_tree_add_24_21_groupi_n_90);
  not csa_tree_add_24_21_groupi_drc_bufs7733(csa_tree_add_24_21_groupi_n_90 ,csa_tree_add_24_21_groupi_n_589);
  not csa_tree_add_24_21_groupi_drc_bufs7739(csa_tree_add_24_21_groupi_n_86 ,csa_tree_add_24_21_groupi_n_84);
  not csa_tree_add_24_21_groupi_drc_bufs7740(csa_tree_add_24_21_groupi_n_85 ,csa_tree_add_24_21_groupi_n_84);
  not csa_tree_add_24_21_groupi_drc_bufs7741(csa_tree_add_24_21_groupi_n_84 ,csa_tree_add_24_21_groupi_n_590);
  not csa_tree_add_24_21_groupi_drc_bufs7747(csa_tree_add_24_21_groupi_n_81 ,csa_tree_add_24_21_groupi_n_79);
  not csa_tree_add_24_21_groupi_drc_bufs7748(csa_tree_add_24_21_groupi_n_80 ,csa_tree_add_24_21_groupi_n_79);
  not csa_tree_add_24_21_groupi_drc_bufs7749(csa_tree_add_24_21_groupi_n_79 ,csa_tree_add_24_21_groupi_n_587);
  not csa_tree_add_24_21_groupi_drc_bufs7751(csa_tree_add_24_21_groupi_n_78 ,csa_tree_add_24_21_groupi_n_76);
  not csa_tree_add_24_21_groupi_drc_bufs7752(csa_tree_add_24_21_groupi_n_77 ,csa_tree_add_24_21_groupi_n_76);
  not csa_tree_add_24_21_groupi_drc_bufs7753(csa_tree_add_24_21_groupi_n_76 ,csa_tree_add_24_21_groupi_n_588);
  not csa_tree_add_24_21_groupi_drc_bufs7755(csa_tree_add_24_21_groupi_n_75 ,csa_tree_add_24_21_groupi_n_73);
  not csa_tree_add_24_21_groupi_drc_bufs7756(csa_tree_add_24_21_groupi_n_74 ,csa_tree_add_24_21_groupi_n_73);
  not csa_tree_add_24_21_groupi_drc_bufs7757(csa_tree_add_24_21_groupi_n_73 ,csa_tree_add_24_21_groupi_n_586);
  not csa_tree_add_24_21_groupi_drc_bufs7759(csa_tree_add_24_21_groupi_n_72 ,csa_tree_add_24_21_groupi_n_70);
  not csa_tree_add_24_21_groupi_drc_bufs7761(csa_tree_add_24_21_groupi_n_70 ,csa_tree_add_24_21_groupi_n_208);
  not csa_tree_add_24_21_groupi_drc_bufs7763(csa_tree_add_24_21_groupi_n_69 ,csa_tree_add_24_21_groupi_n_67);
  not csa_tree_add_24_21_groupi_drc_bufs7765(csa_tree_add_24_21_groupi_n_67 ,csa_tree_add_24_21_groupi_n_214);
  not csa_tree_add_24_21_groupi_drc_bufs7767(csa_tree_add_24_21_groupi_n_66 ,csa_tree_add_24_21_groupi_n_64);
  not csa_tree_add_24_21_groupi_drc_bufs7769(csa_tree_add_24_21_groupi_n_64 ,csa_tree_add_24_21_groupi_n_205);
  not csa_tree_add_24_21_groupi_drc_bufs7771(csa_tree_add_24_21_groupi_n_63 ,csa_tree_add_24_21_groupi_n_61);
  not csa_tree_add_24_21_groupi_drc_bufs7773(csa_tree_add_24_21_groupi_n_61 ,csa_tree_add_24_21_groupi_n_217);
  not csa_tree_add_24_21_groupi_drc_bufs7775(csa_tree_add_24_21_groupi_n_60 ,csa_tree_add_24_21_groupi_n_58);
  not csa_tree_add_24_21_groupi_drc_bufs7777(csa_tree_add_24_21_groupi_n_58 ,csa_tree_add_24_21_groupi_n_211);
  not csa_tree_add_24_21_groupi_drc_bufs7779(csa_tree_add_24_21_groupi_n_57 ,csa_tree_add_24_21_groupi_n_55);
  not csa_tree_add_24_21_groupi_drc_bufs7781(csa_tree_add_24_21_groupi_n_55 ,csa_tree_add_24_21_groupi_n_220);
  not csa_tree_add_24_21_groupi_drc_bufs7783(csa_tree_add_24_21_groupi_n_54 ,csa_tree_add_24_21_groupi_n_52);
  not csa_tree_add_24_21_groupi_drc_bufs7785(csa_tree_add_24_21_groupi_n_52 ,csa_tree_add_22_22_n_86);
  not csa_tree_add_24_21_groupi_drc_bufs7799(csa_tree_add_24_21_groupi_n_43 ,csa_tree_add_24_21_groupi_n_42);
  not csa_tree_add_24_21_groupi_drc_bufs7801(csa_tree_add_24_21_groupi_n_42 ,csa_tree_add_24_21_groupi_n_75);
  not csa_tree_add_24_21_groupi_drc_bufs7803(csa_tree_add_24_21_groupi_n_41 ,csa_tree_add_24_21_groupi_n_40);
  not csa_tree_add_24_21_groupi_drc_bufs7805(csa_tree_add_24_21_groupi_n_40 ,csa_tree_add_24_21_groupi_n_78);
  not csa_tree_add_24_21_groupi_drc_bufs7807(csa_tree_add_24_21_groupi_n_39 ,csa_tree_add_24_21_groupi_n_38);
  not csa_tree_add_24_21_groupi_drc_bufs7809(csa_tree_add_24_21_groupi_n_38 ,csa_tree_add_24_21_groupi_n_81);
  not csa_tree_add_24_21_groupi_drc_bufs7815(csa_tree_add_24_21_groupi_n_34 ,csa_tree_add_24_21_groupi_n_33);
  not csa_tree_add_24_21_groupi_drc_bufs7817(csa_tree_add_24_21_groupi_n_33 ,csa_tree_add_24_21_groupi_n_86);
  not csa_tree_add_24_21_groupi_drc_bufs7823(csa_tree_add_24_21_groupi_n_30 ,csa_tree_add_24_21_groupi_n_29);
  not csa_tree_add_24_21_groupi_drc_bufs7825(csa_tree_add_24_21_groupi_n_29 ,csa_tree_add_24_21_groupi_n_92);
  not csa_tree_add_24_21_groupi_drc_bufs7867(csa_tree_add_24_21_groupi_n_3 ,csa_tree_add_24_21_groupi_n_2);
  not csa_tree_add_24_21_groupi_drc_bufs7869(csa_tree_add_24_21_groupi_n_2 ,csa_tree_add_24_21_groupi_n_120);
  xor csa_tree_add_24_21_groupi_g2(csa_tree_add_24_21_groupi_n_1 ,csa_tree_add_24_21_groupi_n_1670 ,csa_tree_add_24_21_groupi_n_1775);
  xor csa_tree_add_24_21_groupi_g7871(csa_tree_add_24_21_groupi_n_0 ,csa_tree_add_24_21_groupi_n_1749 ,csa_tree_add_24_21_groupi_n_1797);
  xnor csa_tree_add_26_22_groupi_g1024(out3[31] ,csa_tree_add_26_22_groupi_n_343 ,csa_tree_add_26_22_groupi_n_179);
  xnor csa_tree_add_26_22_groupi_g1026(out3[30] ,csa_tree_add_26_22_groupi_n_340 ,csa_tree_add_26_22_groupi_n_124);
  and csa_tree_add_26_22_groupi_g1027(csa_tree_add_26_22_groupi_n_341 ,csa_tree_add_26_22_groupi_n_141 ,csa_tree_add_26_22_groupi_n_340);
  xnor csa_tree_add_26_22_groupi_g1029(out3[29] ,csa_tree_add_26_22_groupi_n_337 ,csa_tree_add_26_22_groupi_n_130);
  and csa_tree_add_26_22_groupi_g1030(csa_tree_add_26_22_groupi_n_338 ,csa_tree_add_26_22_groupi_n_167 ,csa_tree_add_26_22_groupi_n_337);
  xnor csa_tree_add_26_22_groupi_g1032(out3[28] ,csa_tree_add_26_22_groupi_n_334 ,csa_tree_add_26_22_groupi_n_83);
  and csa_tree_add_26_22_groupi_g1033(csa_tree_add_26_22_groupi_n_335 ,csa_tree_add_26_22_groupi_n_163 ,csa_tree_add_26_22_groupi_n_334);
  xnor csa_tree_add_26_22_groupi_g1035(out3[27] ,csa_tree_add_26_22_groupi_n_331 ,csa_tree_add_26_22_groupi_n_99);
  and csa_tree_add_26_22_groupi_g1036(csa_tree_add_26_22_groupi_n_332 ,csa_tree_add_26_22_groupi_n_132 ,csa_tree_add_26_22_groupi_n_331);
  xnor csa_tree_add_26_22_groupi_g1038(out3[26] ,csa_tree_add_26_22_groupi_n_328 ,csa_tree_add_26_22_groupi_n_120);
  and csa_tree_add_26_22_groupi_g1039(csa_tree_add_26_22_groupi_n_329 ,csa_tree_add_26_22_groupi_n_164 ,csa_tree_add_26_22_groupi_n_328);
  xnor csa_tree_add_26_22_groupi_g1041(out3[25] ,csa_tree_add_26_22_groupi_n_325 ,csa_tree_add_26_22_groupi_n_128);
  and csa_tree_add_26_22_groupi_g1042(csa_tree_add_26_22_groupi_n_326 ,csa_tree_add_26_22_groupi_n_161 ,csa_tree_add_26_22_groupi_n_325);
  xnor csa_tree_add_26_22_groupi_g1044(out3[24] ,csa_tree_add_26_22_groupi_n_322 ,csa_tree_add_26_22_groupi_n_87);
  and csa_tree_add_26_22_groupi_g1045(csa_tree_add_26_22_groupi_n_323 ,csa_tree_add_26_22_groupi_n_156 ,csa_tree_add_26_22_groupi_n_322);
  xnor csa_tree_add_26_22_groupi_g1047(out3[23] ,csa_tree_add_26_22_groupi_n_319 ,csa_tree_add_26_22_groupi_n_91);
  and csa_tree_add_26_22_groupi_g1048(csa_tree_add_26_22_groupi_n_320 ,csa_tree_add_26_22_groupi_n_139 ,csa_tree_add_26_22_groupi_n_319);
  xnor csa_tree_add_26_22_groupi_g1050(out3[22] ,csa_tree_add_26_22_groupi_n_316 ,csa_tree_add_26_22_groupi_n_101);
  and csa_tree_add_26_22_groupi_g1051(csa_tree_add_26_22_groupi_n_317 ,csa_tree_add_26_22_groupi_n_133 ,csa_tree_add_26_22_groupi_n_316);
  xnor csa_tree_add_26_22_groupi_g1053(out3[21] ,csa_tree_add_26_22_groupi_n_313 ,csa_tree_add_26_22_groupi_n_122);
  and csa_tree_add_26_22_groupi_g1054(csa_tree_add_26_22_groupi_n_314 ,csa_tree_add_26_22_groupi_n_137 ,csa_tree_add_26_22_groupi_n_313);
  xnor csa_tree_add_26_22_groupi_g1056(out3[20] ,csa_tree_add_26_22_groupi_n_310 ,csa_tree_add_26_22_groupi_n_93);
  and csa_tree_add_26_22_groupi_g1057(csa_tree_add_26_22_groupi_n_311 ,csa_tree_add_26_22_groupi_n_143 ,csa_tree_add_26_22_groupi_n_310);
  xnor csa_tree_add_26_22_groupi_g1059(out3[19] ,csa_tree_add_26_22_groupi_n_307 ,csa_tree_add_26_22_groupi_n_126);
  and csa_tree_add_26_22_groupi_g1060(csa_tree_add_26_22_groupi_n_308 ,csa_tree_add_26_22_groupi_n_166 ,csa_tree_add_26_22_groupi_n_307);
  or csa_tree_add_26_22_groupi_g1061(csa_tree_add_26_22_groupi_n_307 ,csa_tree_add_26_22_groupi_n_157 ,csa_tree_add_26_22_groupi_n_305);
  xnor csa_tree_add_26_22_groupi_g1062(out3[18] ,csa_tree_add_26_22_groupi_n_304 ,csa_tree_add_26_22_groupi_n_178);
  and csa_tree_add_26_22_groupi_g1063(csa_tree_add_26_22_groupi_n_305 ,csa_tree_add_26_22_groupi_n_154 ,csa_tree_add_26_22_groupi_n_304);
  or csa_tree_add_26_22_groupi_g1064(csa_tree_add_26_22_groupi_n_304 ,csa_tree_add_26_22_groupi_n_160 ,csa_tree_add_26_22_groupi_n_302);
  xnor csa_tree_add_26_22_groupi_g1065(out3[17] ,csa_tree_add_26_22_groupi_n_301 ,csa_tree_add_26_22_groupi_n_177);
  and csa_tree_add_26_22_groupi_g1066(csa_tree_add_26_22_groupi_n_302 ,csa_tree_add_26_22_groupi_n_155 ,csa_tree_add_26_22_groupi_n_301);
  or csa_tree_add_26_22_groupi_g1067(csa_tree_add_26_22_groupi_n_301 ,csa_tree_add_26_22_groupi_n_199 ,csa_tree_add_26_22_groupi_n_299);
  xor csa_tree_add_26_22_groupi_g1068(out3[16] ,csa_tree_add_26_22_groupi_n_298 ,csa_tree_add_26_22_groupi_n_212);
  and csa_tree_add_26_22_groupi_g1069(csa_tree_add_26_22_groupi_n_299 ,csa_tree_add_26_22_groupi_n_198 ,csa_tree_add_26_22_groupi_n_298);
  or csa_tree_add_26_22_groupi_g1070(csa_tree_add_26_22_groupi_n_298 ,csa_tree_add_26_22_groupi_n_233 ,csa_tree_add_26_22_groupi_n_296);
  xnor csa_tree_add_26_22_groupi_g1071(out3[15] ,csa_tree_add_26_22_groupi_n_295 ,csa_tree_add_26_22_groupi_n_242);
  and csa_tree_add_26_22_groupi_g1072(csa_tree_add_26_22_groupi_n_296 ,csa_tree_add_26_22_groupi_n_228 ,csa_tree_add_26_22_groupi_n_295);
  or csa_tree_add_26_22_groupi_g1073(csa_tree_add_26_22_groupi_n_295 ,csa_tree_add_26_22_groupi_n_218 ,csa_tree_add_26_22_groupi_n_293);
  xnor csa_tree_add_26_22_groupi_g1074(out3[14] ,csa_tree_add_26_22_groupi_n_292 ,csa_tree_add_26_22_groupi_n_254);
  and csa_tree_add_26_22_groupi_g1075(csa_tree_add_26_22_groupi_n_293 ,csa_tree_add_26_22_groupi_n_221 ,csa_tree_add_26_22_groupi_n_292);
  or csa_tree_add_26_22_groupi_g1076(csa_tree_add_26_22_groupi_n_292 ,csa_tree_add_26_22_groupi_n_220 ,csa_tree_add_26_22_groupi_n_290);
  xnor csa_tree_add_26_22_groupi_g1077(out3[13] ,csa_tree_add_26_22_groupi_n_289 ,csa_tree_add_26_22_groupi_n_253);
  and csa_tree_add_26_22_groupi_g1078(csa_tree_add_26_22_groupi_n_290 ,csa_tree_add_26_22_groupi_n_219 ,csa_tree_add_26_22_groupi_n_289);
  or csa_tree_add_26_22_groupi_g1079(csa_tree_add_26_22_groupi_n_289 ,csa_tree_add_26_22_groupi_n_225 ,csa_tree_add_26_22_groupi_n_287);
  xnor csa_tree_add_26_22_groupi_g1080(out3[12] ,csa_tree_add_26_22_groupi_n_286 ,csa_tree_add_26_22_groupi_n_252);
  and csa_tree_add_26_22_groupi_g1081(csa_tree_add_26_22_groupi_n_287 ,csa_tree_add_26_22_groupi_n_217 ,csa_tree_add_26_22_groupi_n_286);
  or csa_tree_add_26_22_groupi_g1082(csa_tree_add_26_22_groupi_n_286 ,csa_tree_add_26_22_groupi_n_216 ,csa_tree_add_26_22_groupi_n_284);
  xnor csa_tree_add_26_22_groupi_g1083(out3[11] ,csa_tree_add_26_22_groupi_n_283 ,csa_tree_add_26_22_groupi_n_251);
  and csa_tree_add_26_22_groupi_g1084(csa_tree_add_26_22_groupi_n_284 ,csa_tree_add_26_22_groupi_n_213 ,csa_tree_add_26_22_groupi_n_283);
  or csa_tree_add_26_22_groupi_g1085(csa_tree_add_26_22_groupi_n_283 ,csa_tree_add_26_22_groupi_n_222 ,csa_tree_add_26_22_groupi_n_281);
  xnor csa_tree_add_26_22_groupi_g1086(out3[10] ,csa_tree_add_26_22_groupi_n_280 ,csa_tree_add_26_22_groupi_n_250);
  and csa_tree_add_26_22_groupi_g1087(csa_tree_add_26_22_groupi_n_281 ,csa_tree_add_26_22_groupi_n_214 ,csa_tree_add_26_22_groupi_n_280);
  or csa_tree_add_26_22_groupi_g1088(csa_tree_add_26_22_groupi_n_280 ,csa_tree_add_26_22_groupi_n_215 ,csa_tree_add_26_22_groupi_n_278);
  xnor csa_tree_add_26_22_groupi_g1089(out3[9] ,csa_tree_add_26_22_groupi_n_277 ,csa_tree_add_26_22_groupi_n_245);
  and csa_tree_add_26_22_groupi_g1090(csa_tree_add_26_22_groupi_n_278 ,csa_tree_add_26_22_groupi_n_239 ,csa_tree_add_26_22_groupi_n_277);
  or csa_tree_add_26_22_groupi_g1091(csa_tree_add_26_22_groupi_n_277 ,csa_tree_add_26_22_groupi_n_238 ,csa_tree_add_26_22_groupi_n_275);
  xnor csa_tree_add_26_22_groupi_g1092(out3[8] ,csa_tree_add_26_22_groupi_n_274 ,csa_tree_add_26_22_groupi_n_248);
  and csa_tree_add_26_22_groupi_g1093(csa_tree_add_26_22_groupi_n_275 ,csa_tree_add_26_22_groupi_n_237 ,csa_tree_add_26_22_groupi_n_274);
  or csa_tree_add_26_22_groupi_g1094(csa_tree_add_26_22_groupi_n_274 ,csa_tree_add_26_22_groupi_n_236 ,csa_tree_add_26_22_groupi_n_272);
  xnor csa_tree_add_26_22_groupi_g1095(out3[7] ,csa_tree_add_26_22_groupi_n_271 ,csa_tree_add_26_22_groupi_n_247);
  and csa_tree_add_26_22_groupi_g1096(csa_tree_add_26_22_groupi_n_272 ,csa_tree_add_26_22_groupi_n_235 ,csa_tree_add_26_22_groupi_n_271);
  or csa_tree_add_26_22_groupi_g1097(csa_tree_add_26_22_groupi_n_271 ,csa_tree_add_26_22_groupi_n_241 ,csa_tree_add_26_22_groupi_n_269);
  xnor csa_tree_add_26_22_groupi_g1098(out3[6] ,csa_tree_add_26_22_groupi_n_268 ,csa_tree_add_26_22_groupi_n_246);
  and csa_tree_add_26_22_groupi_g1099(csa_tree_add_26_22_groupi_n_269 ,csa_tree_add_26_22_groupi_n_232 ,csa_tree_add_26_22_groupi_n_268);
  or csa_tree_add_26_22_groupi_g1100(csa_tree_add_26_22_groupi_n_268 ,csa_tree_add_26_22_groupi_n_231 ,csa_tree_add_26_22_groupi_n_266);
  xnor csa_tree_add_26_22_groupi_g1101(out3[5] ,csa_tree_add_26_22_groupi_n_265 ,csa_tree_add_26_22_groupi_n_243);
  and csa_tree_add_26_22_groupi_g1102(csa_tree_add_26_22_groupi_n_266 ,csa_tree_add_26_22_groupi_n_230 ,csa_tree_add_26_22_groupi_n_265);
  or csa_tree_add_26_22_groupi_g1103(csa_tree_add_26_22_groupi_n_265 ,csa_tree_add_26_22_groupi_n_229 ,csa_tree_add_26_22_groupi_n_263);
  xnor csa_tree_add_26_22_groupi_g1104(out3[4] ,csa_tree_add_26_22_groupi_n_262 ,csa_tree_add_26_22_groupi_n_244);
  and csa_tree_add_26_22_groupi_g1105(csa_tree_add_26_22_groupi_n_263 ,csa_tree_add_26_22_groupi_n_227 ,csa_tree_add_26_22_groupi_n_262);
  or csa_tree_add_26_22_groupi_g1106(csa_tree_add_26_22_groupi_n_262 ,csa_tree_add_26_22_groupi_n_224 ,csa_tree_add_26_22_groupi_n_260);
  xnor csa_tree_add_26_22_groupi_g1107(out3[3] ,csa_tree_add_26_22_groupi_n_258 ,csa_tree_add_26_22_groupi_n_255);
  and csa_tree_add_26_22_groupi_g1108(csa_tree_add_26_22_groupi_n_260 ,csa_tree_add_26_22_groupi_n_223 ,csa_tree_add_26_22_groupi_n_258);
  xor csa_tree_add_26_22_groupi_g1109(out3[2] ,csa_tree_add_26_22_groupi_n_226 ,csa_tree_add_26_22_groupi_n_256);
  or csa_tree_add_26_22_groupi_g1110(csa_tree_add_26_22_groupi_n_258 ,csa_tree_add_26_22_groupi_n_234 ,csa_tree_add_26_22_groupi_n_257);
  and csa_tree_add_26_22_groupi_g1111(csa_tree_add_26_22_groupi_n_257 ,csa_tree_add_26_22_groupi_n_240 ,csa_tree_add_26_22_groupi_n_226);
  xnor csa_tree_add_26_22_groupi_g1112(csa_tree_add_26_22_groupi_n_256 ,csa_tree_add_26_22_groupi_n_194 ,n_36);
  xnor csa_tree_add_26_22_groupi_g1113(csa_tree_add_26_22_groupi_n_255 ,csa_tree_add_26_22_groupi_n_148 ,csa_tree_add_26_22_groupi_n_206);
  xnor csa_tree_add_26_22_groupi_g1114(csa_tree_add_26_22_groupi_n_254 ,csa_tree_add_26_22_groupi_n_147 ,csa_tree_add_26_22_groupi_n_211);
  xnor csa_tree_add_26_22_groupi_g1115(csa_tree_add_26_22_groupi_n_253 ,csa_tree_add_26_22_groupi_n_150 ,csa_tree_add_26_22_groupi_n_204);
  xnor csa_tree_add_26_22_groupi_g1116(csa_tree_add_26_22_groupi_n_252 ,csa_tree_add_26_22_groupi_n_152 ,csa_tree_add_26_22_groupi_n_203);
  xnor csa_tree_add_26_22_groupi_g1117(csa_tree_add_26_22_groupi_n_251 ,csa_tree_add_26_22_groupi_n_149 ,csa_tree_add_26_22_groupi_n_202);
  xnor csa_tree_add_26_22_groupi_g1118(csa_tree_add_26_22_groupi_n_250 ,csa_tree_add_26_22_groupi_n_171 ,csa_tree_add_26_22_groupi_n_201);
  xor csa_tree_add_26_22_groupi_g1119(out3[1] ,csa_tree_add_26_22_groupi_n_176 ,csa_tree_add_26_22_groupi_n_195);
  xnor csa_tree_add_26_22_groupi_g1120(csa_tree_add_26_22_groupi_n_248 ,csa_tree_add_26_22_groupi_n_151 ,csa_tree_add_26_22_groupi_n_200);
  xnor csa_tree_add_26_22_groupi_g1121(csa_tree_add_26_22_groupi_n_247 ,csa_tree_add_26_22_groupi_n_174 ,csa_tree_add_26_22_groupi_n_205);
  xnor csa_tree_add_26_22_groupi_g1122(csa_tree_add_26_22_groupi_n_246 ,csa_tree_add_26_22_groupi_n_170 ,csa_tree_add_26_22_groupi_n_210);
  xnor csa_tree_add_26_22_groupi_g1123(csa_tree_add_26_22_groupi_n_245 ,csa_tree_add_26_22_groupi_n_175 ,csa_tree_add_26_22_groupi_n_192);
  xnor csa_tree_add_26_22_groupi_g1124(csa_tree_add_26_22_groupi_n_244 ,csa_tree_add_26_22_groupi_n_145 ,csa_tree_add_26_22_groupi_n_207);
  xnor csa_tree_add_26_22_groupi_g1125(csa_tree_add_26_22_groupi_n_243 ,csa_tree_add_26_22_groupi_n_153 ,csa_tree_add_26_22_groupi_n_209);
  xnor csa_tree_add_26_22_groupi_g1126(csa_tree_add_26_22_groupi_n_242 ,csa_tree_add_26_22_groupi_n_146 ,csa_tree_add_26_22_groupi_n_208);
  and csa_tree_add_26_22_groupi_g1127(csa_tree_add_26_22_groupi_n_241 ,csa_tree_add_26_22_groupi_n_170 ,csa_tree_add_26_22_groupi_n_210);
  or csa_tree_add_26_22_groupi_g1128(csa_tree_add_26_22_groupi_n_240 ,n_36 ,csa_tree_add_26_22_groupi_n_193);
  or csa_tree_add_26_22_groupi_g1129(csa_tree_add_26_22_groupi_n_239 ,csa_tree_add_26_22_groupi_n_175 ,csa_tree_add_26_22_groupi_n_192);
  and csa_tree_add_26_22_groupi_g1130(csa_tree_add_26_22_groupi_n_238 ,csa_tree_add_26_22_groupi_n_151 ,csa_tree_add_26_22_groupi_n_200);
  or csa_tree_add_26_22_groupi_g1131(csa_tree_add_26_22_groupi_n_237 ,csa_tree_add_26_22_groupi_n_151 ,csa_tree_add_26_22_groupi_n_200);
  and csa_tree_add_26_22_groupi_g1132(csa_tree_add_26_22_groupi_n_236 ,csa_tree_add_26_22_groupi_n_174 ,csa_tree_add_26_22_groupi_n_205);
  or csa_tree_add_26_22_groupi_g1133(csa_tree_add_26_22_groupi_n_235 ,csa_tree_add_26_22_groupi_n_174 ,csa_tree_add_26_22_groupi_n_205);
  nor csa_tree_add_26_22_groupi_g1134(csa_tree_add_26_22_groupi_n_234 ,csa_tree_add_26_22_groupi_n_0 ,csa_tree_add_26_22_groupi_n_194);
  and csa_tree_add_26_22_groupi_g1135(csa_tree_add_26_22_groupi_n_233 ,csa_tree_add_26_22_groupi_n_146 ,csa_tree_add_26_22_groupi_n_208);
  or csa_tree_add_26_22_groupi_g1136(csa_tree_add_26_22_groupi_n_232 ,csa_tree_add_26_22_groupi_n_170 ,csa_tree_add_26_22_groupi_n_210);
  and csa_tree_add_26_22_groupi_g1137(csa_tree_add_26_22_groupi_n_231 ,csa_tree_add_26_22_groupi_n_153 ,csa_tree_add_26_22_groupi_n_209);
  or csa_tree_add_26_22_groupi_g1138(csa_tree_add_26_22_groupi_n_230 ,csa_tree_add_26_22_groupi_n_153 ,csa_tree_add_26_22_groupi_n_209);
  and csa_tree_add_26_22_groupi_g1139(csa_tree_add_26_22_groupi_n_229 ,csa_tree_add_26_22_groupi_n_145 ,csa_tree_add_26_22_groupi_n_207);
  or csa_tree_add_26_22_groupi_g1140(csa_tree_add_26_22_groupi_n_228 ,csa_tree_add_26_22_groupi_n_146 ,csa_tree_add_26_22_groupi_n_208);
  or csa_tree_add_26_22_groupi_g1141(csa_tree_add_26_22_groupi_n_227 ,csa_tree_add_26_22_groupi_n_145 ,csa_tree_add_26_22_groupi_n_207);
  and csa_tree_add_26_22_groupi_g1142(csa_tree_add_26_22_groupi_n_225 ,csa_tree_add_26_22_groupi_n_152 ,csa_tree_add_26_22_groupi_n_203);
  and csa_tree_add_26_22_groupi_g1143(csa_tree_add_26_22_groupi_n_224 ,csa_tree_add_26_22_groupi_n_148 ,csa_tree_add_26_22_groupi_n_206);
  or csa_tree_add_26_22_groupi_g1144(csa_tree_add_26_22_groupi_n_223 ,csa_tree_add_26_22_groupi_n_148 ,csa_tree_add_26_22_groupi_n_206);
  and csa_tree_add_26_22_groupi_g1145(csa_tree_add_26_22_groupi_n_222 ,csa_tree_add_26_22_groupi_n_171 ,csa_tree_add_26_22_groupi_n_201);
  or csa_tree_add_26_22_groupi_g1146(csa_tree_add_26_22_groupi_n_221 ,csa_tree_add_26_22_groupi_n_147 ,csa_tree_add_26_22_groupi_n_211);
  and csa_tree_add_26_22_groupi_g1147(csa_tree_add_26_22_groupi_n_220 ,csa_tree_add_26_22_groupi_n_150 ,csa_tree_add_26_22_groupi_n_204);
  or csa_tree_add_26_22_groupi_g1148(csa_tree_add_26_22_groupi_n_219 ,csa_tree_add_26_22_groupi_n_150 ,csa_tree_add_26_22_groupi_n_204);
  and csa_tree_add_26_22_groupi_g1149(csa_tree_add_26_22_groupi_n_218 ,csa_tree_add_26_22_groupi_n_147 ,csa_tree_add_26_22_groupi_n_211);
  or csa_tree_add_26_22_groupi_g1150(csa_tree_add_26_22_groupi_n_217 ,csa_tree_add_26_22_groupi_n_152 ,csa_tree_add_26_22_groupi_n_203);
  and csa_tree_add_26_22_groupi_g1151(csa_tree_add_26_22_groupi_n_216 ,csa_tree_add_26_22_groupi_n_149 ,csa_tree_add_26_22_groupi_n_202);
  and csa_tree_add_26_22_groupi_g1152(csa_tree_add_26_22_groupi_n_215 ,csa_tree_add_26_22_groupi_n_175 ,csa_tree_add_26_22_groupi_n_192);
  or csa_tree_add_26_22_groupi_g1153(csa_tree_add_26_22_groupi_n_214 ,csa_tree_add_26_22_groupi_n_171 ,csa_tree_add_26_22_groupi_n_201);
  or csa_tree_add_26_22_groupi_g1154(csa_tree_add_26_22_groupi_n_213 ,csa_tree_add_26_22_groupi_n_149 ,csa_tree_add_26_22_groupi_n_202);
  xnor csa_tree_add_26_22_groupi_g1155(csa_tree_add_26_22_groupi_n_212 ,csa_tree_add_26_22_groupi_n_85 ,csa_tree_add_26_22_groupi_n_173);
  or csa_tree_add_26_22_groupi_g1156(csa_tree_add_26_22_groupi_n_226 ,csa_tree_add_26_22_groupi_n_158 ,csa_tree_add_26_22_groupi_n_197);
  nor csa_tree_add_26_22_groupi_g1157(csa_tree_add_26_22_groupi_n_199 ,csa_tree_add_26_22_groupi_n_85 ,csa_tree_add_26_22_groupi_n_172);
  or csa_tree_add_26_22_groupi_g1158(csa_tree_add_26_22_groupi_n_198 ,csa_tree_add_26_22_groupi_n_84 ,csa_tree_add_26_22_groupi_n_173);
  and csa_tree_add_26_22_groupi_g1159(csa_tree_add_26_22_groupi_n_197 ,csa_tree_add_26_22_groupi_n_176 ,csa_tree_add_26_22_groupi_n_168);
  xnor csa_tree_add_26_22_groupi_g1160(out3[0] ,csa_tree_add_26_22_groupi_n_80 ,in11[0]);
  xnor csa_tree_add_26_22_groupi_g1161(csa_tree_add_26_22_groupi_n_195 ,csa_tree_add_26_22_groupi_n_97 ,n_35);
  xnor csa_tree_add_26_22_groupi_g1162(csa_tree_add_26_22_groupi_n_211 ,csa_tree_add_26_22_groupi_n_68 ,n_48);
  xnor csa_tree_add_26_22_groupi_g1163(csa_tree_add_26_22_groupi_n_210 ,csa_tree_add_26_22_groupi_n_75 ,n_40);
  xnor csa_tree_add_26_22_groupi_g1164(csa_tree_add_26_22_groupi_n_209 ,csa_tree_add_26_22_groupi_n_74 ,n_39);
  xnor csa_tree_add_26_22_groupi_g1165(csa_tree_add_26_22_groupi_n_208 ,csa_tree_add_26_22_groupi_n_72 ,n_49);
  xnor csa_tree_add_26_22_groupi_g1166(csa_tree_add_26_22_groupi_n_207 ,csa_tree_add_26_22_groupi_n_78 ,n_38);
  xnor csa_tree_add_26_22_groupi_g1167(csa_tree_add_26_22_groupi_n_206 ,csa_tree_add_26_22_groupi_n_70 ,n_37);
  xnor csa_tree_add_26_22_groupi_g1168(csa_tree_add_26_22_groupi_n_205 ,csa_tree_add_26_22_groupi_n_77 ,n_41);
  xnor csa_tree_add_26_22_groupi_g1169(csa_tree_add_26_22_groupi_n_204 ,csa_tree_add_26_22_groupi_n_73 ,n_47);
  xnor csa_tree_add_26_22_groupi_g1170(csa_tree_add_26_22_groupi_n_203 ,csa_tree_add_26_22_groupi_n_81 ,n_46);
  xnor csa_tree_add_26_22_groupi_g1171(csa_tree_add_26_22_groupi_n_202 ,csa_tree_add_26_22_groupi_n_103 ,n_45);
  xnor csa_tree_add_26_22_groupi_g1172(csa_tree_add_26_22_groupi_n_201 ,csa_tree_add_26_22_groupi_n_71 ,n_44);
  xnor csa_tree_add_26_22_groupi_g1173(csa_tree_add_26_22_groupi_n_200 ,csa_tree_add_26_22_groupi_n_76 ,n_42);
  not csa_tree_add_26_22_groupi_g1174(csa_tree_add_26_22_groupi_n_193 ,csa_tree_add_26_22_groupi_n_194);
  xnor csa_tree_add_26_22_groupi_g1188(csa_tree_add_26_22_groupi_n_178 ,csa_tree_add_26_22_groupi_n_30 ,csa_tree_add_26_22_groupi_n_89);
  xnor csa_tree_add_26_22_groupi_g1189(csa_tree_add_26_22_groupi_n_177 ,csa_tree_add_26_22_groupi_n_32 ,csa_tree_add_26_22_groupi_n_95);
  xnor csa_tree_add_26_22_groupi_g1190(csa_tree_add_26_22_groupi_n_194 ,csa_tree_add_26_22_groupi_n_37 ,csa_tree_add_26_22_groupi_n_69);
  xnor csa_tree_add_26_22_groupi_g1191(csa_tree_add_26_22_groupi_n_192 ,csa_tree_add_26_22_groupi_n_102 ,n_43);
  not csa_tree_add_26_22_groupi_g1192(csa_tree_add_26_22_groupi_n_172 ,csa_tree_add_26_22_groupi_n_173);
  or csa_tree_add_26_22_groupi_g1194(csa_tree_add_26_22_groupi_n_168 ,n_35 ,csa_tree_add_26_22_groupi_n_96);
  nor csa_tree_add_26_22_groupi_g1202(csa_tree_add_26_22_groupi_n_160 ,csa_tree_add_26_22_groupi_n_32 ,csa_tree_add_26_22_groupi_n_95);
  nor csa_tree_add_26_22_groupi_g1204(csa_tree_add_26_22_groupi_n_158 ,csa_tree_add_26_22_groupi_n_1 ,csa_tree_add_26_22_groupi_n_97);
  nor csa_tree_add_26_22_groupi_g1205(csa_tree_add_26_22_groupi_n_157 ,csa_tree_add_26_22_groupi_n_30 ,csa_tree_add_26_22_groupi_n_89);
  or csa_tree_add_26_22_groupi_g1207(csa_tree_add_26_22_groupi_n_155 ,csa_tree_add_26_22_groupi_n_31 ,csa_tree_add_26_22_groupi_n_94);
  or csa_tree_add_26_22_groupi_g1208(csa_tree_add_26_22_groupi_n_154 ,csa_tree_add_26_22_groupi_n_29 ,csa_tree_add_26_22_groupi_n_88);
  or csa_tree_add_26_22_groupi_g1209(csa_tree_add_26_22_groupi_n_176 ,csa_tree_add_26_22_groupi_n_12 ,csa_tree_add_26_22_groupi_n_110);
  or csa_tree_add_26_22_groupi_g1210(csa_tree_add_26_22_groupi_n_175 ,csa_tree_add_26_22_groupi_n_8 ,csa_tree_add_26_22_groupi_n_107);
  or csa_tree_add_26_22_groupi_g1211(csa_tree_add_26_22_groupi_n_174 ,csa_tree_add_26_22_groupi_n_42 ,csa_tree_add_26_22_groupi_n_117);
  or csa_tree_add_26_22_groupi_g1212(csa_tree_add_26_22_groupi_n_173 ,csa_tree_add_26_22_groupi_n_41 ,csa_tree_add_26_22_groupi_n_116);
  or csa_tree_add_26_22_groupi_g1213(csa_tree_add_26_22_groupi_n_171 ,csa_tree_add_26_22_groupi_n_15 ,csa_tree_add_26_22_groupi_n_104);
  or csa_tree_add_26_22_groupi_g1214(csa_tree_add_26_22_groupi_n_170 ,csa_tree_add_26_22_groupi_n_44 ,csa_tree_add_26_22_groupi_n_115);
  or csa_tree_add_26_22_groupi_g1229(csa_tree_add_26_22_groupi_n_153 ,csa_tree_add_26_22_groupi_n_50 ,csa_tree_add_26_22_groupi_n_113);
  or csa_tree_add_26_22_groupi_g1230(csa_tree_add_26_22_groupi_n_152 ,csa_tree_add_26_22_groupi_n_52 ,csa_tree_add_26_22_groupi_n_108);
  or csa_tree_add_26_22_groupi_g1231(csa_tree_add_26_22_groupi_n_151 ,csa_tree_add_26_22_groupi_n_10 ,csa_tree_add_26_22_groupi_n_118);
  or csa_tree_add_26_22_groupi_g1232(csa_tree_add_26_22_groupi_n_150 ,csa_tree_add_26_22_groupi_n_13 ,csa_tree_add_26_22_groupi_n_109);
  or csa_tree_add_26_22_groupi_g1233(csa_tree_add_26_22_groupi_n_149 ,csa_tree_add_26_22_groupi_n_53 ,csa_tree_add_26_22_groupi_n_106);
  or csa_tree_add_26_22_groupi_g1234(csa_tree_add_26_22_groupi_n_148 ,csa_tree_add_26_22_groupi_n_18 ,csa_tree_add_26_22_groupi_n_105);
  or csa_tree_add_26_22_groupi_g1235(csa_tree_add_26_22_groupi_n_147 ,csa_tree_add_26_22_groupi_n_17 ,csa_tree_add_26_22_groupi_n_111);
  or csa_tree_add_26_22_groupi_g1236(csa_tree_add_26_22_groupi_n_146 ,csa_tree_add_26_22_groupi_n_39 ,csa_tree_add_26_22_groupi_n_114);
  or csa_tree_add_26_22_groupi_g1237(csa_tree_add_26_22_groupi_n_145 ,csa_tree_add_26_22_groupi_n_14 ,csa_tree_add_26_22_groupi_n_112);
  and csa_tree_add_26_22_groupi_g1244(csa_tree_add_26_22_groupi_n_118 ,in11[7] ,csa_tree_add_26_22_groupi_n_48);
  and csa_tree_add_26_22_groupi_g1245(csa_tree_add_26_22_groupi_n_117 ,in11[6] ,csa_tree_add_26_22_groupi_n_49);
  and csa_tree_add_26_22_groupi_g1246(csa_tree_add_26_22_groupi_n_116 ,n_17 ,csa_tree_add_26_22_groupi_n_19);
  and csa_tree_add_26_22_groupi_g1247(csa_tree_add_26_22_groupi_n_115 ,n_7 ,csa_tree_add_26_22_groupi_n_46);
  and csa_tree_add_26_22_groupi_g1248(csa_tree_add_26_22_groupi_n_114 ,n_48 ,csa_tree_add_26_22_groupi_n_21);
  and csa_tree_add_26_22_groupi_g1249(csa_tree_add_26_22_groupi_n_113 ,in11[4] ,csa_tree_add_26_22_groupi_n_9);
  and csa_tree_add_26_22_groupi_g1250(csa_tree_add_26_22_groupi_n_112 ,n_37 ,csa_tree_add_26_22_groupi_n_20);
  and csa_tree_add_26_22_groupi_g1251(csa_tree_add_26_22_groupi_n_111 ,n_15 ,csa_tree_add_26_22_groupi_n_22);
  and csa_tree_add_26_22_groupi_g1252(csa_tree_add_26_22_groupi_n_110 ,in11[0] ,csa_tree_add_26_22_groupi_n_40);
  and csa_tree_add_26_22_groupi_g1253(csa_tree_add_26_22_groupi_n_109 ,n_14 ,csa_tree_add_26_22_groupi_n_47);
  and csa_tree_add_26_22_groupi_g1254(csa_tree_add_26_22_groupi_n_108 ,n_45 ,csa_tree_add_26_22_groupi_n_51);
  and csa_tree_add_26_22_groupi_g1255(csa_tree_add_26_22_groupi_n_107 ,n_42 ,csa_tree_add_26_22_groupi_n_43);
  and csa_tree_add_26_22_groupi_g1256(csa_tree_add_26_22_groupi_n_106 ,n_44 ,csa_tree_add_26_22_groupi_n_45);
  nor csa_tree_add_26_22_groupi_g1257(csa_tree_add_26_22_groupi_n_105 ,csa_tree_add_26_22_groupi_n_37 ,csa_tree_add_26_22_groupi_n_16);
  and csa_tree_add_26_22_groupi_g1258(csa_tree_add_26_22_groupi_n_104 ,n_43 ,csa_tree_add_26_22_groupi_n_11);
  xnor csa_tree_add_26_22_groupi_g1259(csa_tree_add_26_22_groupi_n_103 ,n_13 ,in11[11]);
  xnor csa_tree_add_26_22_groupi_g1260(csa_tree_add_26_22_groupi_n_102 ,n_11 ,in11[9]);
  not csa_tree_add_26_22_groupi_g1269(csa_tree_add_26_22_groupi_n_96 ,csa_tree_add_26_22_groupi_n_97);
  not csa_tree_add_26_22_groupi_g1270(csa_tree_add_26_22_groupi_n_94 ,csa_tree_add_26_22_groupi_n_95);
  not csa_tree_add_26_22_groupi_g1273(csa_tree_add_26_22_groupi_n_88 ,csa_tree_add_26_22_groupi_n_89);
  not csa_tree_add_26_22_groupi_g1275(csa_tree_add_26_22_groupi_n_84 ,csa_tree_add_26_22_groupi_n_85);
  xnor csa_tree_add_26_22_groupi_g1277(csa_tree_add_26_22_groupi_n_81 ,n_14 ,in11[12]);
  xnor csa_tree_add_26_22_groupi_g1278(csa_tree_add_26_22_groupi_n_80 ,n_34 ,n_2);
  xnor csa_tree_add_26_22_groupi_g1280(csa_tree_add_26_22_groupi_n_78 ,n_6 ,in11[4]);
  xnor csa_tree_add_26_22_groupi_g1281(csa_tree_add_26_22_groupi_n_77 ,n_9 ,in11[7]);
  xnor csa_tree_add_26_22_groupi_g1282(csa_tree_add_26_22_groupi_n_76 ,n_10 ,in11[8]);
  xnor csa_tree_add_26_22_groupi_g1283(csa_tree_add_26_22_groupi_n_75 ,n_8 ,in11[6]);
  xnor csa_tree_add_26_22_groupi_g1284(csa_tree_add_26_22_groupi_n_74 ,n_7 ,in11[5]);
  xnor csa_tree_add_26_22_groupi_g1285(csa_tree_add_26_22_groupi_n_73 ,n_15 ,in11[13]);
  xnor csa_tree_add_26_22_groupi_g1286(csa_tree_add_26_22_groupi_n_72 ,n_17 ,in11[15]);
  xnor csa_tree_add_26_22_groupi_g1287(csa_tree_add_26_22_groupi_n_71 ,n_12 ,in11[10]);
  xnor csa_tree_add_26_22_groupi_g1288(csa_tree_add_26_22_groupi_n_70 ,n_5 ,in11[3]);
  xnor csa_tree_add_26_22_groupi_g1289(csa_tree_add_26_22_groupi_n_69 ,n_4 ,in11[2]);
  xnor csa_tree_add_26_22_groupi_g1290(csa_tree_add_26_22_groupi_n_68 ,n_16 ,in11[14]);
  xnor csa_tree_add_26_22_groupi_g1293(csa_tree_add_26_22_groupi_n_97 ,n_3 ,in11[1]);
  xnor csa_tree_add_26_22_groupi_g1294(csa_tree_add_26_22_groupi_n_95 ,n_51 ,n_19);
  xnor csa_tree_add_26_22_groupi_g1299(csa_tree_add_26_22_groupi_n_85 ,n_50 ,n_18);
  and csa_tree_add_26_22_groupi_g1308(csa_tree_add_26_22_groupi_n_53 ,in11[10] ,n_12);
  and csa_tree_add_26_22_groupi_g1309(csa_tree_add_26_22_groupi_n_52 ,in11[11] ,n_13);
  or csa_tree_add_26_22_groupi_g1310(csa_tree_add_26_22_groupi_n_51 ,in11[11] ,n_13);
  and csa_tree_add_26_22_groupi_g1311(csa_tree_add_26_22_groupi_n_50 ,n_38 ,n_6);
  or csa_tree_add_26_22_groupi_g1312(csa_tree_add_26_22_groupi_n_49 ,n_40 ,n_8);
  or csa_tree_add_26_22_groupi_g1313(csa_tree_add_26_22_groupi_n_48 ,n_41 ,n_9);
  or csa_tree_add_26_22_groupi_g1314(csa_tree_add_26_22_groupi_n_47 ,in11[12] ,n_46);
  or csa_tree_add_26_22_groupi_g1315(csa_tree_add_26_22_groupi_n_46 ,in11[5] ,n_39);
  or csa_tree_add_26_22_groupi_g1316(csa_tree_add_26_22_groupi_n_45 ,in11[10] ,n_12);
  and csa_tree_add_26_22_groupi_g1317(csa_tree_add_26_22_groupi_n_44 ,in11[5] ,n_39);
  or csa_tree_add_26_22_groupi_g1318(csa_tree_add_26_22_groupi_n_43 ,in11[8] ,n_10);
  and csa_tree_add_26_22_groupi_g1319(csa_tree_add_26_22_groupi_n_42 ,n_40 ,n_8);
  and csa_tree_add_26_22_groupi_g1320(csa_tree_add_26_22_groupi_n_41 ,in11[15] ,n_49);
  or csa_tree_add_26_22_groupi_g1321(csa_tree_add_26_22_groupi_n_40 ,n_34 ,n_2);
  and csa_tree_add_26_22_groupi_g1322(csa_tree_add_26_22_groupi_n_39 ,in11[14] ,n_16);
  not csa_tree_add_26_22_groupi_g1333(csa_tree_add_26_22_groupi_n_31 ,csa_tree_add_26_22_groupi_n_32);
  not csa_tree_add_26_22_groupi_g1334(csa_tree_add_26_22_groupi_n_29 ,csa_tree_add_26_22_groupi_n_30);
  or csa_tree_add_26_22_groupi_g1338(csa_tree_add_26_22_groupi_n_22 ,in11[13] ,n_47);
  or csa_tree_add_26_22_groupi_g1339(csa_tree_add_26_22_groupi_n_21 ,in11[14] ,n_16);
  or csa_tree_add_26_22_groupi_g1340(csa_tree_add_26_22_groupi_n_20 ,in11[3] ,n_5);
  or csa_tree_add_26_22_groupi_g1341(csa_tree_add_26_22_groupi_n_19 ,in11[15] ,n_49);
  and csa_tree_add_26_22_groupi_g1342(csa_tree_add_26_22_groupi_n_18 ,in11[2] ,n_4);
  and csa_tree_add_26_22_groupi_g1343(csa_tree_add_26_22_groupi_n_17 ,in11[13] ,n_47);
  nor csa_tree_add_26_22_groupi_g1344(csa_tree_add_26_22_groupi_n_16 ,in11[2] ,n_4);
  and csa_tree_add_26_22_groupi_g1345(csa_tree_add_26_22_groupi_n_15 ,in11[9] ,n_11);
  and csa_tree_add_26_22_groupi_g1346(csa_tree_add_26_22_groupi_n_14 ,in11[3] ,n_5);
  and csa_tree_add_26_22_groupi_g1347(csa_tree_add_26_22_groupi_n_13 ,in11[12] ,n_46);
  and csa_tree_add_26_22_groupi_g1348(csa_tree_add_26_22_groupi_n_12 ,n_34 ,n_2);
  or csa_tree_add_26_22_groupi_g1349(csa_tree_add_26_22_groupi_n_11 ,in11[9] ,n_11);
  and csa_tree_add_26_22_groupi_g1350(csa_tree_add_26_22_groupi_n_10 ,n_41 ,n_9);
  or csa_tree_add_26_22_groupi_g1351(csa_tree_add_26_22_groupi_n_9 ,n_38 ,n_6);
  and csa_tree_add_26_22_groupi_g1352(csa_tree_add_26_22_groupi_n_8 ,in11[8] ,n_10);
  or csa_tree_add_26_22_groupi_g1353(csa_tree_add_26_22_groupi_n_37 ,csa_tree_add_26_22_groupi_n_3 ,csa_tree_add_26_22_groupi_n_7);
  or csa_tree_add_26_22_groupi_g1356(csa_tree_add_26_22_groupi_n_32 ,csa_tree_add_26_22_groupi_n_4 ,csa_tree_add_26_22_groupi_n_6);
  or csa_tree_add_26_22_groupi_g1357(csa_tree_add_26_22_groupi_n_30 ,csa_tree_add_26_22_groupi_n_2 ,csa_tree_add_26_22_groupi_n_5);
  not csa_tree_add_26_22_groupi_g1361(csa_tree_add_26_22_groupi_n_7 ,n_3);
  not csa_tree_add_26_22_groupi_g1362(csa_tree_add_26_22_groupi_n_6 ,n_18);
  not csa_tree_add_26_22_groupi_g1363(csa_tree_add_26_22_groupi_n_5 ,n_19);
  not csa_tree_add_26_22_groupi_g1364(csa_tree_add_26_22_groupi_n_4 ,n_50);
  not csa_tree_add_26_22_groupi_g1365(csa_tree_add_26_22_groupi_n_3 ,in11[1]);
  not csa_tree_add_26_22_groupi_g1366(csa_tree_add_26_22_groupi_n_2 ,n_51);
  not csa_tree_add_26_22_groupi_g1367(csa_tree_add_26_22_groupi_n_1 ,n_35);
  not csa_tree_add_26_22_groupi_g1368(csa_tree_add_26_22_groupi_n_0 ,n_36);
  not g7872(csa_tree_add_24_21_groupi_n_468 ,in1[1]);
  buf g7873(csa_tree_add_24_21_groupi_n_395 ,in2[0]);
  not g7874(csa_tree_add_26_22_groupi_n_89 ,n_52);
  not g7875(csa_tree_add_26_22_groupi_n_126 ,n_53);
  not g7877(csa_tree_add_26_22_groupi_n_93 ,n_54);
  not g7878(csa_tree_add_26_22_groupi_n_166 ,csa_tree_add_26_22_groupi_n_126);
  not g7880(csa_tree_add_26_22_groupi_n_122 ,n_55);
  not g7881(csa_tree_add_26_22_groupi_n_143 ,csa_tree_add_26_22_groupi_n_93);
  not g7883(csa_tree_add_26_22_groupi_n_101 ,n_56);
  not g7884(csa_tree_add_26_22_groupi_n_137 ,csa_tree_add_26_22_groupi_n_122);
  buf g7885(csa_tree_add_26_22_groupi_n_310 ,csa_tree_add_26_22_groupi_n_308);
  not g7887(csa_tree_add_26_22_groupi_n_91 ,n_57);
  not g7888(csa_tree_add_26_22_groupi_n_133 ,csa_tree_add_26_22_groupi_n_101);
  buf g7889(csa_tree_add_26_22_groupi_n_313 ,csa_tree_add_26_22_groupi_n_311);
  not g7891(csa_tree_add_26_22_groupi_n_87 ,n_58);
  not g7892(csa_tree_add_26_22_groupi_n_139 ,csa_tree_add_26_22_groupi_n_91);
  buf g7893(csa_tree_add_26_22_groupi_n_316 ,csa_tree_add_26_22_groupi_n_314);
  not g7895(csa_tree_add_26_22_groupi_n_128 ,n_59);
  not g7896(csa_tree_add_26_22_groupi_n_156 ,csa_tree_add_26_22_groupi_n_87);
  buf g7897(csa_tree_add_26_22_groupi_n_319 ,csa_tree_add_26_22_groupi_n_317);
  not g7899(csa_tree_add_26_22_groupi_n_120 ,n_60);
  not g7900(csa_tree_add_26_22_groupi_n_161 ,csa_tree_add_26_22_groupi_n_128);
  buf g7901(csa_tree_add_26_22_groupi_n_322 ,csa_tree_add_26_22_groupi_n_320);
  not g7903(csa_tree_add_26_22_groupi_n_99 ,n_61);
  not g7904(csa_tree_add_26_22_groupi_n_164 ,csa_tree_add_26_22_groupi_n_120);
  buf g7905(csa_tree_add_26_22_groupi_n_325 ,csa_tree_add_26_22_groupi_n_323);
  not g7907(csa_tree_add_26_22_groupi_n_83 ,n_62);
  not g7908(csa_tree_add_26_22_groupi_n_132 ,csa_tree_add_26_22_groupi_n_99);
  buf g7909(csa_tree_add_26_22_groupi_n_328 ,csa_tree_add_26_22_groupi_n_326);
  not g7911(csa_tree_add_26_22_groupi_n_130 ,n_63);
  not g7912(csa_tree_add_26_22_groupi_n_163 ,csa_tree_add_26_22_groupi_n_83);
  buf g7913(csa_tree_add_26_22_groupi_n_331 ,csa_tree_add_26_22_groupi_n_329);
  not g7915(csa_tree_add_26_22_groupi_n_124 ,n_64);
  not g7916(csa_tree_add_26_22_groupi_n_167 ,csa_tree_add_26_22_groupi_n_130);
  buf g7917(csa_tree_add_26_22_groupi_n_334 ,csa_tree_add_26_22_groupi_n_332);
  not g7920(csa_tree_add_26_22_groupi_n_141 ,csa_tree_add_26_22_groupi_n_124);
  buf g7921(csa_tree_add_26_22_groupi_n_337 ,csa_tree_add_26_22_groupi_n_335);
  not g7922(csa_tree_add_26_22_groupi_n_179 ,n_65);
  buf g7923(csa_tree_add_26_22_groupi_n_340 ,csa_tree_add_26_22_groupi_n_338);
  buf g7924(csa_tree_add_26_22_groupi_n_343 ,csa_tree_add_26_22_groupi_n_341);

endmodule

module top(in1, in2, in3, in4, in5, out1);

  input [31:0] in1, in2, in3;

  input [5:0] in4, in5;

  output [63:0] out1;
  wire [31:0] in1, in2, in3;
  wire [5:0] in4, in5;
  wire [63:0] out1;
  wire csa_tree_add_8_49_groupi_n_0, csa_tree_add_8_49_groupi_n_1, csa_tree_add_8_49_groupi_n_2, csa_tree_add_8_49_groupi_n_3, csa_tree_add_8_49_groupi_n_4, csa_tree_add_8_49_groupi_n_5, csa_tree_add_8_49_groupi_n_6, csa_tree_add_8_49_groupi_n_7;
  wire csa_tree_add_8_49_groupi_n_8, csa_tree_add_8_49_groupi_n_9, csa_tree_add_8_49_groupi_n_10, csa_tree_add_8_49_groupi_n_11, csa_tree_add_8_49_groupi_n_12, csa_tree_add_8_49_groupi_n_13, csa_tree_add_8_49_groupi_n_14, csa_tree_add_8_49_groupi_n_15;
  wire csa_tree_add_8_49_groupi_n_16, csa_tree_add_8_49_groupi_n_17, csa_tree_add_8_49_groupi_n_18, csa_tree_add_8_49_groupi_n_19, csa_tree_add_8_49_groupi_n_20, csa_tree_add_8_49_groupi_n_21, csa_tree_add_8_49_groupi_n_22, csa_tree_add_8_49_groupi_n_23;
  wire csa_tree_add_8_49_groupi_n_24, csa_tree_add_8_49_groupi_n_25, csa_tree_add_8_49_groupi_n_26, csa_tree_add_8_49_groupi_n_27, csa_tree_add_8_49_groupi_n_28, csa_tree_add_8_49_groupi_n_29, csa_tree_add_8_49_groupi_n_30, csa_tree_add_8_49_groupi_n_31;
  wire csa_tree_add_8_49_groupi_n_32, csa_tree_add_8_49_groupi_n_33, csa_tree_add_8_49_groupi_n_34, csa_tree_add_8_49_groupi_n_35, csa_tree_add_8_49_groupi_n_36, csa_tree_add_8_49_groupi_n_37, csa_tree_add_8_49_groupi_n_38, csa_tree_add_8_49_groupi_n_39;
  wire csa_tree_add_8_49_groupi_n_40, csa_tree_add_8_49_groupi_n_41, csa_tree_add_8_49_groupi_n_42, csa_tree_add_8_49_groupi_n_43, csa_tree_add_8_49_groupi_n_44, csa_tree_add_8_49_groupi_n_45, csa_tree_add_8_49_groupi_n_46, csa_tree_add_8_49_groupi_n_47;
  wire csa_tree_add_8_49_groupi_n_48, csa_tree_add_8_49_groupi_n_49, csa_tree_add_8_49_groupi_n_50, csa_tree_add_8_49_groupi_n_51, csa_tree_add_8_49_groupi_n_52, csa_tree_add_8_49_groupi_n_53, csa_tree_add_8_49_groupi_n_54, csa_tree_add_8_49_groupi_n_55;
  wire csa_tree_add_8_49_groupi_n_56, csa_tree_add_8_49_groupi_n_57, csa_tree_add_8_49_groupi_n_58, csa_tree_add_8_49_groupi_n_59, csa_tree_add_8_49_groupi_n_60, csa_tree_add_8_49_groupi_n_61, csa_tree_add_8_49_groupi_n_62, csa_tree_add_8_49_groupi_n_63;
  wire csa_tree_add_8_49_groupi_n_64, csa_tree_add_8_49_groupi_n_65, csa_tree_add_8_49_groupi_n_66, csa_tree_add_8_49_groupi_n_67, csa_tree_add_8_49_groupi_n_68, csa_tree_add_8_49_groupi_n_69, csa_tree_add_8_49_groupi_n_70, csa_tree_add_8_49_groupi_n_71;
  wire csa_tree_add_8_49_groupi_n_72, csa_tree_add_8_49_groupi_n_73, csa_tree_add_8_49_groupi_n_74, csa_tree_add_8_49_groupi_n_75, csa_tree_add_8_49_groupi_n_76, csa_tree_add_8_49_groupi_n_77, csa_tree_add_8_49_groupi_n_78, csa_tree_add_8_49_groupi_n_79;
  wire csa_tree_add_8_49_groupi_n_80, csa_tree_add_8_49_groupi_n_81, csa_tree_add_8_49_groupi_n_82, csa_tree_add_8_49_groupi_n_83, csa_tree_add_8_49_groupi_n_84, csa_tree_add_8_49_groupi_n_85, csa_tree_add_8_49_groupi_n_86, csa_tree_add_8_49_groupi_n_87;
  wire csa_tree_add_8_49_groupi_n_88, csa_tree_add_8_49_groupi_n_89, csa_tree_add_8_49_groupi_n_90, csa_tree_add_8_49_groupi_n_91, csa_tree_add_8_49_groupi_n_92, csa_tree_add_8_49_groupi_n_93, csa_tree_add_8_49_groupi_n_94, csa_tree_add_8_49_groupi_n_95;
  wire csa_tree_add_8_49_groupi_n_96, csa_tree_add_8_49_groupi_n_97, csa_tree_add_8_49_groupi_n_98, csa_tree_add_8_49_groupi_n_99, csa_tree_add_8_49_groupi_n_100, csa_tree_add_8_49_groupi_n_101, csa_tree_add_8_49_groupi_n_102, csa_tree_add_8_49_groupi_n_103;
  wire csa_tree_add_8_49_groupi_n_104, csa_tree_add_8_49_groupi_n_105, csa_tree_add_8_49_groupi_n_106, csa_tree_add_8_49_groupi_n_107, csa_tree_add_8_49_groupi_n_108, csa_tree_add_8_49_groupi_n_109, csa_tree_add_8_49_groupi_n_110, csa_tree_add_8_49_groupi_n_111;
  wire csa_tree_add_8_49_groupi_n_112, csa_tree_add_8_49_groupi_n_113, csa_tree_add_8_49_groupi_n_114, csa_tree_add_8_49_groupi_n_115, csa_tree_add_8_49_groupi_n_116, csa_tree_add_8_49_groupi_n_117, csa_tree_add_8_49_groupi_n_118, csa_tree_add_8_49_groupi_n_119;
  wire csa_tree_add_8_49_groupi_n_120, csa_tree_add_8_49_groupi_n_121, csa_tree_add_8_49_groupi_n_122, csa_tree_add_8_49_groupi_n_123, csa_tree_add_8_49_groupi_n_124, csa_tree_add_8_49_groupi_n_125, csa_tree_add_8_49_groupi_n_126, csa_tree_add_8_49_groupi_n_127;
  wire csa_tree_add_8_49_groupi_n_128, csa_tree_add_8_49_groupi_n_129, csa_tree_add_8_49_groupi_n_130, csa_tree_add_8_49_groupi_n_131, csa_tree_add_8_49_groupi_n_132, csa_tree_add_8_49_groupi_n_133, csa_tree_add_8_49_groupi_n_134, csa_tree_add_8_49_groupi_n_135;
  wire csa_tree_add_8_49_groupi_n_136, csa_tree_add_8_49_groupi_n_137, csa_tree_add_8_49_groupi_n_138, csa_tree_add_8_49_groupi_n_139, csa_tree_add_8_49_groupi_n_140, csa_tree_add_8_49_groupi_n_141, csa_tree_add_8_49_groupi_n_142, csa_tree_add_8_49_groupi_n_143;
  wire csa_tree_add_8_49_groupi_n_144, csa_tree_add_8_49_groupi_n_145, csa_tree_add_8_49_groupi_n_146, csa_tree_add_8_49_groupi_n_147, csa_tree_add_8_49_groupi_n_148, csa_tree_add_8_49_groupi_n_149, csa_tree_add_8_49_groupi_n_150, csa_tree_add_8_49_groupi_n_151;
  wire csa_tree_add_8_49_groupi_n_152, csa_tree_add_8_49_groupi_n_153, csa_tree_add_8_49_groupi_n_154, csa_tree_add_8_49_groupi_n_155, csa_tree_add_8_49_groupi_n_156, csa_tree_add_8_49_groupi_n_157, csa_tree_add_8_49_groupi_n_158, csa_tree_add_8_49_groupi_n_159;
  wire csa_tree_add_8_49_groupi_n_160, csa_tree_add_8_49_groupi_n_161, csa_tree_add_8_49_groupi_n_162, csa_tree_add_8_49_groupi_n_163, csa_tree_add_8_49_groupi_n_164, csa_tree_add_8_49_groupi_n_165, csa_tree_add_8_49_groupi_n_166, csa_tree_add_8_49_groupi_n_167;
  wire csa_tree_add_8_49_groupi_n_168, csa_tree_add_8_49_groupi_n_169, csa_tree_add_8_49_groupi_n_170, csa_tree_add_8_49_groupi_n_171, csa_tree_add_8_49_groupi_n_172, csa_tree_add_8_49_groupi_n_173, csa_tree_add_8_49_groupi_n_174, csa_tree_add_8_49_groupi_n_175;
  wire csa_tree_add_8_49_groupi_n_176, csa_tree_add_8_49_groupi_n_177, csa_tree_add_8_49_groupi_n_178, csa_tree_add_8_49_groupi_n_179, csa_tree_add_8_49_groupi_n_180, csa_tree_add_8_49_groupi_n_181, csa_tree_add_8_49_groupi_n_182, csa_tree_add_8_49_groupi_n_183;
  wire csa_tree_add_8_49_groupi_n_184, csa_tree_add_8_49_groupi_n_185, csa_tree_add_8_49_groupi_n_186, csa_tree_add_8_49_groupi_n_187, csa_tree_add_8_49_groupi_n_188, csa_tree_add_8_49_groupi_n_189, csa_tree_add_8_49_groupi_n_190, csa_tree_add_8_49_groupi_n_191;
  wire csa_tree_add_8_49_groupi_n_192, csa_tree_add_8_49_groupi_n_193, csa_tree_add_8_49_groupi_n_194, csa_tree_add_8_49_groupi_n_195, csa_tree_add_8_49_groupi_n_196, csa_tree_add_8_49_groupi_n_197, csa_tree_add_8_49_groupi_n_198, csa_tree_add_8_49_groupi_n_199;
  wire csa_tree_add_8_49_groupi_n_200, csa_tree_add_8_49_groupi_n_201, csa_tree_add_8_49_groupi_n_202, csa_tree_add_8_49_groupi_n_203, csa_tree_add_8_49_groupi_n_204, csa_tree_add_8_49_groupi_n_205, csa_tree_add_8_49_groupi_n_206, csa_tree_add_8_49_groupi_n_207;
  wire csa_tree_add_8_49_groupi_n_208, csa_tree_add_8_49_groupi_n_209, csa_tree_add_8_49_groupi_n_210, csa_tree_add_8_49_groupi_n_211, csa_tree_add_8_49_groupi_n_212, csa_tree_add_8_49_groupi_n_213, csa_tree_add_8_49_groupi_n_214, csa_tree_add_8_49_groupi_n_215;
  wire csa_tree_add_8_49_groupi_n_216, csa_tree_add_8_49_groupi_n_217, csa_tree_add_8_49_groupi_n_218, csa_tree_add_8_49_groupi_n_219, csa_tree_add_8_49_groupi_n_220, csa_tree_add_8_49_groupi_n_221, csa_tree_add_8_49_groupi_n_222, csa_tree_add_8_49_groupi_n_223;
  wire csa_tree_add_8_49_groupi_n_224, csa_tree_add_8_49_groupi_n_225, csa_tree_add_8_49_groupi_n_226, csa_tree_add_8_49_groupi_n_227, csa_tree_add_8_49_groupi_n_228, csa_tree_add_8_49_groupi_n_229, csa_tree_add_8_49_groupi_n_230, csa_tree_add_8_49_groupi_n_231;
  wire csa_tree_add_8_49_groupi_n_232, csa_tree_add_8_49_groupi_n_233, csa_tree_add_8_49_groupi_n_234, csa_tree_add_8_49_groupi_n_235, csa_tree_add_8_49_groupi_n_236, csa_tree_add_8_49_groupi_n_237, csa_tree_add_8_49_groupi_n_238, csa_tree_add_8_49_groupi_n_239;
  wire csa_tree_add_8_49_groupi_n_240, csa_tree_add_8_49_groupi_n_241, csa_tree_add_8_49_groupi_n_242, csa_tree_add_8_49_groupi_n_243, csa_tree_add_8_49_groupi_n_244, csa_tree_add_8_49_groupi_n_245, csa_tree_add_8_49_groupi_n_246, csa_tree_add_8_49_groupi_n_247;
  wire csa_tree_add_8_49_groupi_n_248, csa_tree_add_8_49_groupi_n_249, csa_tree_add_8_49_groupi_n_250, csa_tree_add_8_49_groupi_n_251, csa_tree_add_8_49_groupi_n_252, csa_tree_add_8_49_groupi_n_253, csa_tree_add_8_49_groupi_n_254, csa_tree_add_8_49_groupi_n_255;
  wire csa_tree_add_8_49_groupi_n_256, csa_tree_add_8_49_groupi_n_257, csa_tree_add_8_49_groupi_n_258, csa_tree_add_8_49_groupi_n_259, csa_tree_add_8_49_groupi_n_260, csa_tree_add_8_49_groupi_n_261, csa_tree_add_8_49_groupi_n_262, csa_tree_add_8_49_groupi_n_263;
  wire csa_tree_add_8_49_groupi_n_264, csa_tree_add_8_49_groupi_n_265, csa_tree_add_8_49_groupi_n_266, csa_tree_add_8_49_groupi_n_267, csa_tree_add_8_49_groupi_n_268, csa_tree_add_8_49_groupi_n_269, csa_tree_add_8_49_groupi_n_270, csa_tree_add_8_49_groupi_n_271;
  wire csa_tree_add_8_49_groupi_n_272, csa_tree_add_8_49_groupi_n_273, csa_tree_add_8_49_groupi_n_274, csa_tree_add_8_49_groupi_n_275, csa_tree_add_8_49_groupi_n_276, csa_tree_add_8_49_groupi_n_277, csa_tree_add_8_49_groupi_n_278, csa_tree_add_8_49_groupi_n_279;
  wire csa_tree_add_8_49_groupi_n_280, csa_tree_add_8_49_groupi_n_281, csa_tree_add_8_49_groupi_n_282, csa_tree_add_8_49_groupi_n_283, csa_tree_add_8_49_groupi_n_284, csa_tree_add_8_49_groupi_n_285, csa_tree_add_8_49_groupi_n_286, csa_tree_add_8_49_groupi_n_287;
  wire csa_tree_add_8_49_groupi_n_288, csa_tree_add_8_49_groupi_n_289, csa_tree_add_8_49_groupi_n_290, csa_tree_add_8_49_groupi_n_291, csa_tree_add_8_49_groupi_n_292, csa_tree_add_8_49_groupi_n_293, csa_tree_add_8_49_groupi_n_294, csa_tree_add_8_49_groupi_n_295;
  wire csa_tree_add_8_49_groupi_n_296, csa_tree_add_8_49_groupi_n_297, csa_tree_add_8_49_groupi_n_298, csa_tree_add_8_49_groupi_n_299, csa_tree_add_8_49_groupi_n_300, csa_tree_add_8_49_groupi_n_301, csa_tree_add_8_49_groupi_n_302, csa_tree_add_8_49_groupi_n_303;
  wire csa_tree_add_8_49_groupi_n_304, csa_tree_add_8_49_groupi_n_305, csa_tree_add_8_49_groupi_n_306, csa_tree_add_8_49_groupi_n_307, csa_tree_add_8_49_groupi_n_308, csa_tree_add_8_49_groupi_n_309, csa_tree_add_8_49_groupi_n_310, csa_tree_add_8_49_groupi_n_311;
  wire csa_tree_add_8_49_groupi_n_312, csa_tree_add_8_49_groupi_n_313, csa_tree_add_8_49_groupi_n_314, csa_tree_add_8_49_groupi_n_315, csa_tree_add_8_49_groupi_n_316, csa_tree_add_8_49_groupi_n_317, csa_tree_add_8_49_groupi_n_318, csa_tree_add_8_49_groupi_n_319;
  wire csa_tree_add_8_49_groupi_n_320, csa_tree_add_8_49_groupi_n_321, csa_tree_add_8_49_groupi_n_322, csa_tree_add_8_49_groupi_n_323, csa_tree_add_8_49_groupi_n_324, csa_tree_add_8_49_groupi_n_325, csa_tree_add_8_49_groupi_n_326, csa_tree_add_8_49_groupi_n_327;
  wire csa_tree_add_8_49_groupi_n_328, csa_tree_add_8_49_groupi_n_329, csa_tree_add_8_49_groupi_n_330, csa_tree_add_8_49_groupi_n_331, csa_tree_add_8_49_groupi_n_332, csa_tree_add_8_49_groupi_n_333, csa_tree_add_8_49_groupi_n_334, csa_tree_add_8_49_groupi_n_335;
  wire csa_tree_add_8_49_groupi_n_336, csa_tree_add_8_49_groupi_n_337, csa_tree_add_8_49_groupi_n_338, csa_tree_add_8_49_groupi_n_339, csa_tree_add_8_49_groupi_n_340, csa_tree_add_8_49_groupi_n_341, csa_tree_add_8_49_groupi_n_342, csa_tree_add_8_49_groupi_n_343;
  wire csa_tree_add_8_49_groupi_n_344, csa_tree_add_8_49_groupi_n_345, csa_tree_add_8_49_groupi_n_346, csa_tree_add_8_49_groupi_n_347, csa_tree_add_8_49_groupi_n_348, csa_tree_add_8_49_groupi_n_349, csa_tree_add_8_49_groupi_n_350, csa_tree_add_8_49_groupi_n_351;
  wire csa_tree_add_8_49_groupi_n_352, csa_tree_add_8_49_groupi_n_353, csa_tree_add_8_49_groupi_n_354, csa_tree_add_8_49_groupi_n_355, csa_tree_add_8_49_groupi_n_356, csa_tree_add_8_49_groupi_n_357, csa_tree_add_8_49_groupi_n_358, csa_tree_add_8_49_groupi_n_359;
  wire csa_tree_add_8_49_groupi_n_360, csa_tree_add_8_49_groupi_n_361, csa_tree_add_8_49_groupi_n_362, csa_tree_add_8_49_groupi_n_363, csa_tree_add_8_49_groupi_n_364, csa_tree_add_8_49_groupi_n_365, csa_tree_add_8_49_groupi_n_366, csa_tree_add_8_49_groupi_n_367;
  wire csa_tree_add_8_49_groupi_n_368, csa_tree_add_8_49_groupi_n_369, csa_tree_add_8_49_groupi_n_370, csa_tree_add_8_49_groupi_n_371, csa_tree_add_8_49_groupi_n_372, csa_tree_add_8_49_groupi_n_373, csa_tree_add_8_49_groupi_n_374, csa_tree_add_8_49_groupi_n_375;
  wire csa_tree_add_8_49_groupi_n_376, csa_tree_add_8_49_groupi_n_377, csa_tree_add_8_49_groupi_n_378, csa_tree_add_8_49_groupi_n_379, csa_tree_add_8_49_groupi_n_380, csa_tree_add_8_49_groupi_n_381, csa_tree_add_8_49_groupi_n_382, csa_tree_add_8_49_groupi_n_383;
  wire csa_tree_add_8_49_groupi_n_384, csa_tree_add_8_49_groupi_n_385, csa_tree_add_8_49_groupi_n_386, csa_tree_add_8_49_groupi_n_387, csa_tree_add_8_49_groupi_n_388, csa_tree_add_8_49_groupi_n_389, csa_tree_add_8_49_groupi_n_390, csa_tree_add_8_49_groupi_n_391;
  wire csa_tree_add_8_49_groupi_n_392, csa_tree_add_8_49_groupi_n_393, csa_tree_add_8_49_groupi_n_394, csa_tree_add_8_49_groupi_n_395, csa_tree_add_8_49_groupi_n_396, csa_tree_add_8_49_groupi_n_397, csa_tree_add_8_49_groupi_n_398, csa_tree_add_8_49_groupi_n_399;
  wire csa_tree_add_8_49_groupi_n_400, csa_tree_add_8_49_groupi_n_401, csa_tree_add_8_49_groupi_n_402, csa_tree_add_8_49_groupi_n_403, csa_tree_add_8_49_groupi_n_404, csa_tree_add_8_49_groupi_n_405, csa_tree_add_8_49_groupi_n_406, csa_tree_add_8_49_groupi_n_407;
  wire csa_tree_add_8_49_groupi_n_408, csa_tree_add_8_49_groupi_n_409, csa_tree_add_8_49_groupi_n_410, csa_tree_add_8_49_groupi_n_411, csa_tree_add_8_49_groupi_n_412, csa_tree_add_8_49_groupi_n_413, csa_tree_add_8_49_groupi_n_414, csa_tree_add_8_49_groupi_n_415;
  wire csa_tree_add_8_49_groupi_n_416, csa_tree_add_8_49_groupi_n_417, csa_tree_add_8_49_groupi_n_418, csa_tree_add_8_49_groupi_n_419, csa_tree_add_8_49_groupi_n_420, csa_tree_add_8_49_groupi_n_421, csa_tree_add_8_49_groupi_n_422, csa_tree_add_8_49_groupi_n_423;
  wire csa_tree_add_8_49_groupi_n_424, csa_tree_add_8_49_groupi_n_425, csa_tree_add_8_49_groupi_n_426, csa_tree_add_8_49_groupi_n_427, csa_tree_add_8_49_groupi_n_428, csa_tree_add_8_49_groupi_n_429, csa_tree_add_8_49_groupi_n_430, csa_tree_add_8_49_groupi_n_431;
  wire csa_tree_add_8_49_groupi_n_432, csa_tree_add_8_49_groupi_n_433, csa_tree_add_8_49_groupi_n_434, csa_tree_add_8_49_groupi_n_435, csa_tree_add_8_49_groupi_n_436, csa_tree_add_8_49_groupi_n_437, csa_tree_add_8_49_groupi_n_438, csa_tree_add_8_49_groupi_n_439;
  wire csa_tree_add_8_49_groupi_n_440, csa_tree_add_8_49_groupi_n_441, csa_tree_add_8_49_groupi_n_442, csa_tree_add_8_49_groupi_n_443, csa_tree_add_8_49_groupi_n_444, csa_tree_add_8_49_groupi_n_445, csa_tree_add_8_49_groupi_n_446, csa_tree_add_8_49_groupi_n_447;
  wire csa_tree_add_8_49_groupi_n_449, csa_tree_add_8_49_groupi_n_450, csa_tree_add_8_49_groupi_n_451, csa_tree_add_8_49_groupi_n_452, csa_tree_add_8_49_groupi_n_453, csa_tree_add_8_49_groupi_n_454, csa_tree_add_8_49_groupi_n_455, csa_tree_add_8_49_groupi_n_456;
  wire csa_tree_add_8_49_groupi_n_457, csa_tree_add_8_49_groupi_n_458, csa_tree_add_8_49_groupi_n_459, csa_tree_add_8_49_groupi_n_460, csa_tree_add_8_49_groupi_n_461, csa_tree_add_8_49_groupi_n_462, csa_tree_add_8_49_groupi_n_463, csa_tree_add_8_49_groupi_n_464;
  wire csa_tree_add_8_49_groupi_n_465, csa_tree_add_8_49_groupi_n_466, csa_tree_add_8_49_groupi_n_467, csa_tree_add_8_49_groupi_n_468, csa_tree_add_8_49_groupi_n_469, csa_tree_add_8_49_groupi_n_470, csa_tree_add_8_49_groupi_n_471, csa_tree_add_8_49_groupi_n_472;
  wire csa_tree_add_8_49_groupi_n_473, csa_tree_add_8_49_groupi_n_474, csa_tree_add_8_49_groupi_n_475, csa_tree_add_8_49_groupi_n_476, csa_tree_add_8_49_groupi_n_477, csa_tree_add_8_49_groupi_n_478, csa_tree_add_8_49_groupi_n_479, csa_tree_add_8_49_groupi_n_480;
  wire csa_tree_add_8_49_groupi_n_481, csa_tree_add_8_49_groupi_n_482, csa_tree_add_8_49_groupi_n_483, csa_tree_add_8_49_groupi_n_484, csa_tree_add_8_49_groupi_n_485, csa_tree_add_8_49_groupi_n_486, csa_tree_add_8_49_groupi_n_487, csa_tree_add_8_49_groupi_n_488;
  wire csa_tree_add_8_49_groupi_n_489, csa_tree_add_8_49_groupi_n_490, csa_tree_add_8_49_groupi_n_491, csa_tree_add_8_49_groupi_n_492, csa_tree_add_8_49_groupi_n_493, csa_tree_add_8_49_groupi_n_494, csa_tree_add_8_49_groupi_n_495, csa_tree_add_8_49_groupi_n_496;
  wire csa_tree_add_8_49_groupi_n_497, csa_tree_add_8_49_groupi_n_498, csa_tree_add_8_49_groupi_n_499, csa_tree_add_8_49_groupi_n_500, csa_tree_add_8_49_groupi_n_501, csa_tree_add_8_49_groupi_n_502, csa_tree_add_8_49_groupi_n_503, csa_tree_add_8_49_groupi_n_504;
  wire csa_tree_add_8_49_groupi_n_505, csa_tree_add_8_49_groupi_n_506, csa_tree_add_8_49_groupi_n_507, csa_tree_add_8_49_groupi_n_508, csa_tree_add_8_49_groupi_n_509, csa_tree_add_8_49_groupi_n_510, csa_tree_add_8_49_groupi_n_511, csa_tree_add_8_49_groupi_n_512;
  wire csa_tree_add_8_49_groupi_n_513, csa_tree_add_8_49_groupi_n_514, csa_tree_add_8_49_groupi_n_515, csa_tree_add_8_49_groupi_n_516, csa_tree_add_8_49_groupi_n_517, csa_tree_add_8_49_groupi_n_518, csa_tree_add_8_49_groupi_n_519, csa_tree_add_8_49_groupi_n_520;
  wire csa_tree_add_8_49_groupi_n_521, csa_tree_add_8_49_groupi_n_522, csa_tree_add_8_49_groupi_n_523, csa_tree_add_8_49_groupi_n_524, csa_tree_add_8_49_groupi_n_525, csa_tree_add_8_49_groupi_n_526, csa_tree_add_8_49_groupi_n_527, csa_tree_add_8_49_groupi_n_528;
  wire csa_tree_add_8_49_groupi_n_529, csa_tree_add_8_49_groupi_n_530, csa_tree_add_8_49_groupi_n_531, csa_tree_add_8_49_groupi_n_532, csa_tree_add_8_49_groupi_n_533, csa_tree_add_8_49_groupi_n_534, csa_tree_add_8_49_groupi_n_535, csa_tree_add_8_49_groupi_n_536;
  wire csa_tree_add_8_49_groupi_n_537, csa_tree_add_8_49_groupi_n_538, csa_tree_add_8_49_groupi_n_539, csa_tree_add_8_49_groupi_n_540, csa_tree_add_8_49_groupi_n_541, csa_tree_add_8_49_groupi_n_542, csa_tree_add_8_49_groupi_n_543, csa_tree_add_8_49_groupi_n_544;
  wire csa_tree_add_8_49_groupi_n_545, csa_tree_add_8_49_groupi_n_546, csa_tree_add_8_49_groupi_n_547, csa_tree_add_8_49_groupi_n_548, csa_tree_add_8_49_groupi_n_549, csa_tree_add_8_49_groupi_n_550, csa_tree_add_8_49_groupi_n_551, csa_tree_add_8_49_groupi_n_552;
  wire csa_tree_add_8_49_groupi_n_553, csa_tree_add_8_49_groupi_n_554, csa_tree_add_8_49_groupi_n_556, csa_tree_add_8_49_groupi_n_557, csa_tree_add_8_49_groupi_n_558, csa_tree_add_8_49_groupi_n_559, csa_tree_add_8_49_groupi_n_560, csa_tree_add_8_49_groupi_n_561;
  wire csa_tree_add_8_49_groupi_n_562, csa_tree_add_8_49_groupi_n_563, csa_tree_add_8_49_groupi_n_564, csa_tree_add_8_49_groupi_n_565, csa_tree_add_8_49_groupi_n_566, csa_tree_add_8_49_groupi_n_567, csa_tree_add_8_49_groupi_n_568, csa_tree_add_8_49_groupi_n_569;
  wire csa_tree_add_8_49_groupi_n_570, csa_tree_add_8_49_groupi_n_571, csa_tree_add_8_49_groupi_n_572, csa_tree_add_8_49_groupi_n_574, csa_tree_add_8_49_groupi_n_576, csa_tree_add_8_49_groupi_n_577, csa_tree_add_8_49_groupi_n_579, csa_tree_add_8_49_groupi_n_580;
  wire csa_tree_add_8_49_groupi_n_582, csa_tree_add_8_49_groupi_n_583, csa_tree_add_8_49_groupi_n_585, csa_tree_add_8_49_groupi_n_586, csa_tree_add_8_49_groupi_n_588, csa_tree_add_8_49_groupi_n_589, csa_tree_add_8_49_groupi_n_591, csa_tree_add_8_49_groupi_n_592;
  wire csa_tree_add_8_49_groupi_n_594, csa_tree_add_8_49_groupi_n_595, csa_tree_add_8_49_groupi_n_597, csa_tree_add_8_49_groupi_n_598, csa_tree_add_8_49_groupi_n_600, csa_tree_add_8_49_groupi_n_601, csa_tree_add_8_49_groupi_n_603, csa_tree_add_8_49_groupi_n_604;
  wire csa_tree_add_8_49_groupi_n_606, csa_tree_add_8_49_groupi_n_607, csa_tree_add_8_49_groupi_n_609, csa_tree_add_8_49_groupi_n_610, csa_tree_add_8_49_groupi_n_612, csa_tree_add_8_49_groupi_n_613, csa_tree_add_8_49_groupi_n_615, csa_tree_add_8_49_groupi_n_616;
  wire csa_tree_add_8_49_groupi_n_618, csa_tree_add_8_49_groupi_n_619, csa_tree_add_8_49_groupi_n_621, csa_tree_add_8_49_groupi_n_622, csa_tree_add_8_49_groupi_n_624, csa_tree_add_8_49_groupi_n_625, csa_tree_add_8_49_groupi_n_627, csa_tree_add_8_49_groupi_n_628;
  wire csa_tree_add_8_49_groupi_n_630, csa_tree_add_8_49_groupi_n_631, csa_tree_add_8_49_groupi_n_633, csa_tree_add_8_49_groupi_n_634, csa_tree_add_8_49_groupi_n_636, csa_tree_add_8_49_groupi_n_637, csa_tree_add_8_49_groupi_n_639, csa_tree_add_8_49_groupi_n_640;
  wire csa_tree_add_8_49_groupi_n_642, csa_tree_add_8_49_groupi_n_643, csa_tree_add_8_49_groupi_n_645, csa_tree_add_8_49_groupi_n_646, csa_tree_add_8_49_groupi_n_648, csa_tree_add_8_49_groupi_n_649, csa_tree_add_8_49_groupi_n_651, csa_tree_add_8_49_groupi_n_652;
  wire csa_tree_add_8_49_groupi_n_654, csa_tree_add_8_49_groupi_n_655, csa_tree_add_8_49_groupi_n_657, csa_tree_add_8_49_groupi_n_658, csa_tree_add_8_49_groupi_n_660, csa_tree_add_8_49_groupi_n_661, csa_tree_add_8_49_groupi_n_663, csa_tree_add_8_49_groupi_n_664;
  wire csa_tree_add_8_49_groupi_n_666, csa_tree_add_8_49_groupi_n_667, csa_tree_add_8_49_groupi_n_669, csa_tree_add_8_49_groupi_n_670, csa_tree_add_8_49_groupi_n_672, csa_tree_add_8_49_groupi_n_673, csa_tree_add_8_49_groupi_n_675, csa_tree_add_8_49_groupi_n_676;
  wire csa_tree_add_8_49_groupi_n_678, csa_tree_add_8_49_groupi_n_679, csa_tree_add_8_49_groupi_n_681, csa_tree_add_8_49_groupi_n_682, csa_tree_add_8_49_groupi_n_684, csa_tree_add_8_49_groupi_n_685, csa_tree_add_8_49_groupi_n_687, csa_tree_add_8_49_groupi_n_688;
  wire csa_tree_add_8_49_groupi_n_690, csa_tree_add_8_49_groupi_n_691, csa_tree_add_8_49_groupi_n_693, csa_tree_add_8_49_groupi_n_694, csa_tree_add_8_49_groupi_n_696, csa_tree_add_8_49_groupi_n_697, csa_tree_add_8_49_groupi_n_699, csa_tree_add_8_49_groupi_n_700;
  wire csa_tree_add_8_49_groupi_n_702, csa_tree_add_8_49_groupi_n_703, csa_tree_add_8_49_groupi_n_705, csa_tree_add_8_49_groupi_n_706, csa_tree_add_8_49_groupi_n_708, csa_tree_add_8_49_groupi_n_709, csa_tree_add_8_49_groupi_n_711, csa_tree_add_8_49_groupi_n_712;
  wire csa_tree_add_8_49_groupi_n_714, csa_tree_add_8_49_groupi_n_715, csa_tree_add_8_49_groupi_n_717, csa_tree_add_8_49_groupi_n_718, csa_tree_add_8_49_groupi_n_720, csa_tree_add_8_49_groupi_n_721, csa_tree_add_8_49_groupi_n_723, csa_tree_add_8_49_groupi_n_724;
  wire csa_tree_add_8_49_groupi_n_726, csa_tree_add_8_49_groupi_n_727, csa_tree_add_8_49_groupi_n_729, csa_tree_add_8_49_groupi_n_730, csa_tree_add_8_49_groupi_n_732, csa_tree_add_8_49_groupi_n_733, csa_tree_add_8_49_groupi_n_735, csa_tree_add_8_49_groupi_n_736;
  wire csa_tree_add_8_49_groupi_n_738, csa_tree_add_8_49_groupi_n_739, csa_tree_add_8_49_groupi_n_741, csa_tree_add_8_49_groupi_n_742, csa_tree_add_8_49_groupi_n_744, csa_tree_add_8_49_groupi_n_745, csa_tree_add_8_49_groupi_n_747, csa_tree_add_8_49_groupi_n_748;
  wire csa_tree_add_8_49_groupi_n_750, csa_tree_add_8_49_groupi_n_751, csa_tree_add_8_49_groupi_n_753, n_0, n_1, n_2, n_3, n_4;
  wire n_5, n_6, n_7, n_8, n_9, n_10, n_9, n_10;
  wire n_17, n_18, n_17, n_18, n_17, n_18, n_17, n_18;
  wire n_17, n_18, n_27, n_28, n_17, n_18, n_27, n_28;
  wire n_29, n_30, n_17, n_18, n_146, n_148, n_148, n_36;
  wire n_37, n_146, n_148, n_213, n_41, n_42, n_132, n_134;
  wire n_132, n_134, n_134, n_143, n_265, n_50, n_51, n_52;
  wire n_132, n_134, n_143, n_265, n_265, n_143, n_265, n_60;
  wire n_61, n_132, n_134, n_134, n_132, n_134, n_134, n_132;
  wire n_134, n_70, n_71, n_117, n_119, n_119, n_117, n_119;
  wire n_119, n_108, n_110, n_110, n_123, n_125, n_125, n_123;
  wire n_125, n_125, n_108, n_110, n_110, n_117, n_119, n_119;
  wire n_108, n_110, n_110, n_117, n_119, n_119, n_108, n_110;
  wire n_110, n_108, n_110, n_110, n_108, n_110, n_110, n_108;
  wire n_110, n_110, n_123, n_125, n_125, n_117, n_119, n_119;
  wire n_117, n_119, n_119, n_123, n_125, n_125, n_123, n_125;
  wire n_125, n_123, n_125, n_125, n_176, n_178, n_178, n_132;
  wire n_134, n_134, n_132, n_134, n_134, n_143, n_265, n_265;
  wire n_141, n_143, n_143, n_144, n_259, n_146, n_148, n_148;
  wire n_123, n_125, n_125, n_123, n_125, n_125, n_176, n_178;
  wire n_178, n_108, n_110, n_110, n_117, n_119, n_119, n_176;
  wire n_178, n_178, n_117, n_119, n_119, n_176, n_178, n_178;
  wire n_176, n_178, n_178, n_176, n_178, n_178, n_176, n_178;
  wire n_178, n_176, n_178, n_178, n_146, n_148, n_187, n_188;
  wire n_189, n_214, n_216, n_216, n_195, n_197, n_195, n_197;
  wire n_197, n_197, n_199, n_235, n_237, n_237, n_204, n_204;
  wire n_206, n_206, n_208, n_208, n_210, n_210, n_213, n_212;
  wire n_213, n_214, n_216, n_216, n_217, n_218, n_219, n_235;
  wire n_237, n_237, n_235, n_237, n_237, n_235, n_237, n_237;
  wire n_235, n_237, n_237, n_213, n_342, n_342, n_235, n_237;
  wire n_237, n_343, n_195, n_195, n_235, n_237, n_245, n_245;
  wire n_245, n_245, n_249, n_249, n_249, n_249, n_253, n_253;
  wire n_253, n_253, n_257, n_257, n_257, n_257, n_259, n_141;
  wire n_265, n_262, n_265, n_141, n_265, n_266, n_265, n_342;
  wire n_212, n_342, n_271, n_272, n_273, n_274, n_275, n_276;
  wire n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284;
  wire n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292;
  wire n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300;
  wire n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308;
  wire n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316;
  wire n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324;
  wire n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332;
  wire n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_342;
  wire n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348;
  wire n_349, n_350, n_351, n_352, n_353, n_354, n_355, n_356;
  wire n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364;
  wire n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372;
  wire n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380;
  wire n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388;
  wire n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396;
  wire n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404;
  wire n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412;
  wire n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420;
  wire n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444;
  wire n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460;
  wire n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476;
  wire n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484;
  wire n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492;
  wire n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500;
  wire n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508;
  wire n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516;
  wire n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524;
  wire n_525, n_526, n_527, n_528, n_529, n_530, n_531, n_532;
  wire n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540;
  wire n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548;
  wire n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556;
  wire n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564;
  wire n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572;
  wire n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580;
  wire n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_588;
  wire n_589, n_590, n_591, n_592, n_593, n_594, n_595, n_596;
  wire n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604;
  wire n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612;
  wire n_613, n_614, n_615, n_616, n_617, n_618, n_619, n_620;
  wire n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628;
  wire n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636;
  wire n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644;
  wire n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652;
  wire n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660;
  wire n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668;
  wire n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676;
  wire n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684;
  wire n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692;
  wire n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700;
  wire n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708;
  wire n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716;
  wire n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724;
  wire n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732;
  wire n_733, n_734, n_735, n_736, n_737, n_738, n_739, n_740;
  wire n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748;
  wire n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756;
  wire n_757, n_758, n_759, n_760, n_761, n_762, n_763, n_764;
  wire n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772;
  wire n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780;
  wire n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788;
  wire n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796;
  wire n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804;
  wire n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812;
  wire n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820;
  wire n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828;
  wire n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836;
  wire n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844;
  wire n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852;
  wire n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860;
  wire n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868;
  wire n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876;
  wire n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884;
  wire n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892;
  wire n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900;
  wire n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908;
  wire n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_930, n_929, n_930;
  wire n_937, n_938, n_937, n_938, n_937, n_938, n_937, n_938;
  wire n_937, n_938, n_947, n_948, n_937, n_938, n_947, n_948;
  wire n_949, n_950, n_937, n_938, n_1066, n_1068, n_1068, n_956;
  wire n_957, n_1066, n_1068, n_1133, n_961, n_962, n_1052, n_1054;
  wire n_1052, n_1054, n_1054, n_1063, n_1185, n_970, n_971, n_972;
  wire n_1052, n_1054, n_1063, n_1185, n_1185, n_1063, n_1185, n_980;
  wire n_981, n_1052, n_1054, n_1054, n_1052, n_1054, n_1054, n_1052;
  wire n_1054, n_990, n_991, n_1037, n_1039, n_1039, n_1037, n_1039;
  wire n_1039, n_1028, n_1030, n_1030, n_1043, n_1045, n_1045, n_1043;
  wire n_1045, n_1045, n_1028, n_1030, n_1030, n_1037, n_1039, n_1039;
  wire n_1028, n_1030, n_1030, n_1037, n_1039, n_1039, n_1028, n_1030;
  wire n_1030, n_1028, n_1030, n_1030, n_1028, n_1030, n_1030, n_1028;
  wire n_1030, n_1030, n_1043, n_1045, n_1045, n_1037, n_1039, n_1039;
  wire n_1037, n_1039, n_1039, n_1043, n_1045, n_1045, n_1043, n_1045;
  wire n_1045, n_1043, n_1045, n_1045, n_1096, n_1098, n_1098, n_1052;
  wire n_1054, n_1054, n_1052, n_1054, n_1054, n_1063, n_1185, n_1185;
  wire n_1061, n_1063, n_1063, n_1064, n_1179, n_1066, n_1068, n_1068;
  wire n_1043, n_1045, n_1045, n_1043, n_1045, n_1045, n_1096, n_1098;
  wire n_1098, n_1028, n_1030, n_1030, n_1037, n_1039, n_1039, n_1096;
  wire n_1098, n_1098, n_1037, n_1039, n_1039, n_1096, n_1098, n_1098;
  wire n_1096, n_1098, n_1098, n_1096, n_1098, n_1098, n_1096, n_1098;
  wire n_1098, n_1096, n_1098, n_1098, n_1066, n_1068, n_1107, n_1108;
  wire n_1109, n_1134, n_1136, n_1136, n_1115, n_1117, n_1115, n_1117;
  wire n_1117, n_1117, n_1119, n_1152, n_1154, n_1154, n_1124, n_1124;
  wire n_1126, n_1126, n_1128, n_1128, n_1130, n_1130, n_1133, n_1132;
  wire n_1133, n_1134, n_1136, n_1136, n_1137, n_1138, n_1139, n_1152;
  wire n_1154, n_1154, n_1152, n_1154, n_1154, n_1152, n_1154, n_1154;
  wire n_1133, n_1262, n_1262, n_1152, n_1154, n_1154, n_1152, n_1154;
  wire n_1154, n_1263, n_1115, n_1115, n_1152, n_1154, n_1165, n_1165;
  wire n_1165, n_1165, n_1169, n_1169, n_1169, n_1169, n_1173, n_1173;
  wire n_1173, n_1173, n_1177, n_1177, n_1177, n_1177, n_1179, n_1061;
  wire n_1185, n_1182, n_1185, n_1061, n_1185, n_1186, n_1185, n_1262;
  wire n_1132, n_1262, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196;
  wire n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204;
  wire n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212;
  wire n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220;
  wire n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228;
  wire n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236;
  wire n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244;
  wire n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252;
  wire n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1262;
  wire n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268;
  wire n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276;
  wire n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284;
  wire n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292;
  wire n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300;
  wire n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308;
  wire n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316;
  wire n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324;
  wire n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332;
  wire n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340;
  wire n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348;
  wire n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356;
  wire n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364;
  wire n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372;
  wire n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380;
  wire n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388;
  wire n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396;
  wire n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404;
  wire n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412;
  wire n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420;
  wire n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428;
  wire n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436;
  wire n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444;
  wire n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452;
  wire n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460;
  wire n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468;
  wire n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476;
  wire n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484;
  wire n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492;
  wire n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500;
  wire n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508;
  wire n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516;
  wire n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524;
  wire n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532;
  wire n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540;
  wire n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548;
  wire n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556;
  wire n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564;
  wire n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572;
  wire n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580;
  wire n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588;
  wire n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596;
  wire n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604;
  wire n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612;
  wire n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620;
  wire n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628;
  wire n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636;
  wire n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644;
  wire n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652;
  wire n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660;
  wire n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668;
  wire n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676;
  wire n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684;
  wire n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692;
  wire n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700;
  wire n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708;
  wire n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716;
  wire n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724;
  wire n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732;
  wire n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740;
  wire n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748;
  wire n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756;
  wire n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764;
  wire n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772;
  wire n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780;
  wire n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788;
  wire n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796;
  wire n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804;
  wire n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812;
  wire n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820;
  wire n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828;
  wire n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836;
  wire n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844;
  wire n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852;
  wire n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860;
  wire n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868;
  wire n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876;
  wire n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884;
  wire n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892;
  wire n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900;
  wire n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908;
  wire n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916;
  wire n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924;
  wire n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932;
  wire n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940;
  or g5390__2398(n_1874 ,n_1521 ,n_1805);
  or g5391__5107(n_1873 ,n_1583 ,n_1810);
  or g5392__6260(n_1861 ,n_1749 ,n_1811);
  or g5393__4319(n_1872 ,n_1561 ,n_1809);
  or g5394__8428(n_1871 ,n_1666 ,n_1808);
  or g5395__5526(n_1870 ,n_1642 ,n_1807);
  or g5396__6783(n_1875 ,n_1443 ,n_1812);
  or g5397__3680(n_1864 ,n_1719 ,n_1804);
  or g5398__1617(n_1868 ,n_1663 ,n_927);
  or g5399__2802(n_1866 ,n_1707 ,n_925);
  or g5400__1705(n_1865 ,n_1693 ,n_1803);
  or g5401__5122(n_1869 ,n_1634 ,n_1806);
  or g5402__8246(n_1863 ,n_1702 ,n_924);
  or g5403__7098(n_1862 ,n_1697 ,n_926);
  or g5404__6131(n_1867 ,n_1694 ,n_928);
  and g5405__1881(n_1876 ,in5[5] ,n_1800);
  and g5406__5115(n_1812 ,in5[5] ,n_1793);
  and g5407__7482(n_1811 ,in5[5] ,n_1794);
  or g5408__4733(n_1859 ,n_1768 ,n_1791);
  or g5409__6161(n_1857 ,n_1766 ,n_1789);
  or g5410__9315(n_1856 ,n_923 ,n_1788);
  or g5411__9945(n_1854 ,n_1764 ,n_1790);
  and g5412__2883(n_1810 ,in5[5] ,n_1795);
  or g5413__2346(n_1852 ,n_1729 ,n_1772);
  or g5414__1666(n_1851 ,n_1692 ,n_1786);
  or g5415__7410(n_1850 ,n_1725 ,n_1785);
  or g5416__6417(n_1849 ,n_1723 ,n_1784);
  or g5417__5477(n_1847 ,n_1718 ,n_1783);
  or g5418__2398(n_1846 ,n_1745 ,n_1782);
  and g5419__5107(n_1844 ,n_1185 ,n_1800);
  and g5420__6260(n_1843 ,n_971 ,n_1793);
  and g5421__4319(n_1842 ,n_1054 ,n_1799);
  and g5422__8428(n_1841 ,n_981 ,n_1795);
  and g5423__5526(n_1840 ,n_1054 ,n_1796);
  and g5424__6783(n_1839 ,n_1185 ,n_1797);
  and g5425__3680(n_1838 ,n_1054 ,n_1802);
  and g5426__1617(n_1837 ,n_962 ,n_1801);
  and g5427__2802(n_1809 ,in5[5] ,n_1796);
  and g5428__1705(n_1832 ,n_1054 ,n_1798);
  and g5429__5122(n_1829 ,n_1185 ,n_1794);
  and g5430__8246(n_1808 ,in5[5] ,n_1797);
  and g5431__7098(n_1807 ,in5[5] ,n_1802);
  and g5432__6131(n_1806 ,in5[5] ,n_1801);
  and g5434__1881(n_1805 ,in5[5] ,n_1799);
  and g5435__5115(n_1804 ,in5[5] ,n_1798);
  or g5437__7482(n_1860 ,n_1747 ,n_1769);
  or g5438__4733(n_1845 ,n_1751 ,n_1781);
  and g5439__6161(n_1831 ,n_1054 ,n_1773);
  and g5440__9315(n_1834 ,n_1185 ,n_1774);
  or g5441__9945(n_1848 ,n_922 ,n_1771);
  nor g5445__2883(n_1803 ,n_1054 ,n_1779);
  or g5446__2346(n_1853 ,n_1770 ,n_1792);
  or g5447__1666(n_1858 ,n_1767 ,n_1780);
  or g5448__7410(n_1855 ,n_1765 ,n_1787);
  and g5449__6417(n_1836 ,n_1054 ,n_1776);
  and g5450__5477(n_1833 ,n_991 ,n_1778);
  and g5451__2398(n_1830 ,n_1054 ,n_1775);
  and g5452__5107(n_1835 ,n_1185 ,n_1777);
  or g5453__6260(n_1792 ,n_1635 ,n_1730);
  or g5454__4319(n_1791 ,n_1444 ,n_1743);
  or g5455__8428(n_1790 ,n_1643 ,n_1731);
  or g5456__5526(n_1789 ,n_1575 ,n_1740);
  or g5457__6783(n_1788 ,n_1562 ,n_1737);
  or g5458__3680(n_1787 ,n_1664 ,n_1734);
  or g5459__1617(n_1786 ,n_1726 ,n_1727);
  or g5460__2802(n_1785 ,n_921 ,n_1724);
  or g5461__1705(n_1784 ,n_1733 ,n_1696);
  or g5462__5122(n_1783 ,n_1636 ,n_1744);
  or g5463__8246(n_1782 ,n_1619 ,n_1700);
  or g5464__7098(n_1781 ,n_920 ,n_1695);
  or g5465__6131(n_1780 ,n_1520 ,n_1742);
  or g5466__1881(n_1802 ,n_1712 ,n_1711);
  or g5467__5115(n_1801 ,n_1698 ,n_1710);
  or g5468__7482(n_1800 ,n_1739 ,n_1738);
  or g5469__4733(n_1799 ,n_1705 ,n_1746);
  or g5470__6161(n_1798 ,n_1571 ,n_1703);
  or g5471__9315(n_1797 ,n_1714 ,n_1713);
  or g5472__9945(n_1796 ,n_1699 ,n_1715);
  or g5473__2883(n_1795 ,n_1732 ,n_1736);
  or g5474__2346(n_1794 ,n_1509 ,n_1748);
  or g5475__1666(n_1793 ,n_1735 ,n_1716);
  not g5476(n_1779 ,n_1778);
  or g5482__7410(n_1772 ,n_1665 ,n_1728);
  or g5483__6417(n_1771 ,n_1640 ,n_1741);
  and g5484__5477(n_1824 ,n_1054 ,n_1720);
  and g5485__2398(n_1821 ,n_962 ,n_1721);
  and g5486__5107(n_1828 ,n_1054 ,n_1753);
  and g5487__6260(n_1827 ,n_1185 ,n_1755);
  and g5488__4319(n_1826 ,n_1054 ,n_1757);
  and g5489__8428(n_1825 ,n_1185 ,n_1759);
  and g5490__5526(n_1823 ,n_1054 ,n_1761);
  and g5491__6783(n_1822 ,n_971 ,n_1763);
  nor g5492__3680(n_1770 ,n_1185 ,n_1722);
  nor g5493__1617(n_1769 ,n_1054 ,n_1752);
  nor g5494__2802(n_1768 ,n_1054 ,n_1754);
  nor g5495__1705(n_1767 ,n_1054 ,n_1756);
  nor g5496__5122(n_1766 ,n_1185 ,n_1758);
  nor g5497__8246(n_1765 ,n_1054 ,n_1760);
  nor g5498__7098(n_1764 ,n_972 ,n_1762);
  or g5500__6131(n_1778 ,n_1639 ,n_1704);
  or g5501__1881(n_1777 ,n_1638 ,n_1708);
  or g5502__5115(n_1776 ,n_1637 ,n_1709);
  or g5503__7482(n_1775 ,n_1518 ,n_1750);
  or g5504__4733(n_1774 ,n_1641 ,n_1706);
  or g5505__6161(n_1773 ,n_1564 ,n_1701);
  not g5506(n_1763 ,n_1762);
  not g5507(n_1761 ,n_1760);
  not g5508(n_1759 ,n_1758);
  not g5509(n_1757 ,n_1756);
  not g5510(n_1755 ,n_1754);
  not g5511(n_1753 ,n_1752);
  nor g5512__9315(n_1751 ,n_1154 ,n_1691);
  nor g5513__9945(n_1750 ,in5[4] ,n_1677);
  nor g5514__2883(n_1749 ,n_1154 ,n_1668);
  nor g5515__2346(n_1748 ,in5[4] ,n_1691);
  nor g5516__1666(n_1747 ,n_1154 ,n_1687);
  nor g5517__7410(n_1746 ,in5[4] ,n_1683);
  nor g5518__6417(n_1745 ,n_1154 ,n_1677);
  and g5519__5477(n_1744 ,n_1117 ,n_1656);
  nor g5520__2398(n_1743 ,n_1154 ,n_1676);
  nor g5521__5107(n_1742 ,n_1154 ,n_1683);
  nor g5522__6260(n_1741 ,n_1262 ,n_1655);
  nor g5523__4319(n_1740 ,n_1262 ,n_1679);
  and g5524__8428(n_1739 ,in5[4] ,n_1672);
  nor g5525__5526(n_1738 ,in5[4] ,n_1687);
  nor g5526__6783(n_1737 ,n_1154 ,n_1678);
  nor g5527__3680(n_1736 ,in5[4] ,n_1679);
  and g5528__1617(n_1735 ,in5[4] ,n_1688);
  nor g5529__2802(n_1734 ,n_1154 ,n_1674);
  and g5530__1705(n_1733 ,in5[5] ,n_1690);
  and g5531__5122(n_1732 ,in5[4] ,n_1685);
  nor g5532__8246(n_1731 ,n_1262 ,n_1670);
  nor g5533__7098(n_1730 ,n_1154 ,n_1669);
  and g5534__6131(n_1729 ,in5[5] ,n_1684);
  nor g5535__1881(n_1728 ,n_1154 ,n_1667);
  nor g5536__5115(n_1727 ,n_1154 ,n_1662);
  and g5537__7482(n_1726 ,in5[5] ,n_1682);
  and g5538__4733(n_1725 ,n_1117 ,n_1647);
  nor g5539__6161(n_1724 ,n_1154 ,n_1648);
  nor g5540__9315(n_1723 ,n_1154 ,n_1653);
  or g5541__9945(n_1762 ,in5[4] ,n_1671);
  or g5542__2883(n_1760 ,in5[4] ,n_1675);
  or g5543__2346(n_1758 ,in5[4] ,n_1686);
  or g5544__1666(n_1756 ,in5[4] ,n_1651);
  or g5545__7410(n_1754 ,in5[4] ,n_1689);
  or g5546__6417(n_1752 ,in5[4] ,n_1673);
  not g5547(n_1722 ,n_1721);
  nor g5549__5477(n_1719 ,n_1154 ,n_1654);
  nor g5550__2398(n_1718 ,n_1154 ,n_1661);
  and g5551__5107(n_1819 ,n_1185 ,n_1682);
  and g5552__6260(n_1717 ,n_1054 ,n_1690);
  nor g5553__4319(n_1716 ,in5[4] ,n_1676);
  nor g5554__8428(n_1715 ,in5[4] ,n_1678);
  nor g5555__5526(n_1714 ,n_1136 ,n_1675);
  nor g5556__6783(n_1713 ,in5[4] ,n_1674);
  nor g5557__3680(n_1712 ,n_1068 ,n_1671);
  nor g5558__1617(n_1711 ,in5[4] ,n_1670);
  nor g5559__2802(n_1710 ,in5[4] ,n_1669);
  nor g5560__1705(n_1709 ,in5[4] ,n_1667);
  nor g5561__5122(n_1708 ,in5[4] ,n_1662);
  and g5562__8246(n_1707 ,n_1133 ,n_1647);
  nor g5563__7098(n_1706 ,in5[4] ,n_1648);
  nor g5564__6131(n_1705 ,n_1068 ,n_1651);
  nor g5565__1881(n_1704 ,in5[4] ,n_1653);
  nor g5566__5115(n_1703 ,in5[4] ,n_1655);
  and g5567__7482(n_1702 ,n_1133 ,n_1656);
  and g5568__4733(n_1820 ,n_1185 ,n_1684);
  nor g5569__6161(n_1701 ,in5[4] ,n_1661);
  and g5570__9315(n_1700 ,n_1117 ,n_1680);
  nor g5572__9945(n_1699 ,n_1109 ,n_1660);
  nor g5573__2883(n_1698 ,n_1068 ,n_1658);
  nor g5574__2346(n_1697 ,n_1154 ,n_1681);
  and g5575__1666(n_1696 ,n_1117 ,n_1649);
  and g5576__7410(n_1818 ,n_1054 ,n_1652);
  nor g5577__6417(n_1695 ,n_1115 ,n_1668);
  nor g5578__5477(n_1694 ,n_1154 ,n_1645);
  nor g5579__2398(n_1693 ,n_1154 ,n_1650);
  and g5580__5107(n_1692 ,n_1117 ,n_1646);
  and g5582__6260(n_1721 ,n_1068 ,n_1657);
  and g5583__4319(n_1720 ,n_1068 ,n_1659);
  not g5584(n_1689 ,n_1688);
  not g5585(n_1686 ,n_1685);
  not g5586(n_1681 ,n_1680);
  not g5587(n_1673 ,n_1672);
  nor g5588__8428(n_1666 ,n_1154 ,n_1632);
  nor g5589__5526(n_1665 ,n_1115 ,n_1633);
  nor g5590__6783(n_1664 ,n_1119 ,n_1632);
  nor g5591__3680(n_1663 ,n_1154 ,n_1633);
  and g5592__1617(n_1691 ,n_1625 ,n_1623);
  and g5593__2802(n_1690 ,n_1068 ,n_1589);
  or g5594__1705(n_1688 ,n_1626 ,n_1616);
  and g5595__5122(n_1687 ,n_1622 ,n_1606);
  or g5596__8246(n_1685 ,n_1621 ,n_1620);
  and g5597__7098(n_1684 ,n_1068 ,n_1590);
  and g5598__6131(n_1683 ,n_1629 ,n_1627);
  and g5599__1881(n_1682 ,n_1068 ,n_1588);
  or g5600__5115(n_1680 ,n_1569 ,n_1614);
  and g5601__7482(n_1679 ,n_1617 ,n_1624);
  and g5602__4733(n_1678 ,n_1631 ,n_1613);
  and g5603__6161(n_1677 ,n_1630 ,n_1618);
  and g5604__9315(n_1676 ,n_1607 ,n_1602);
  and g5605__9945(n_1675 ,n_1516 ,n_1610);
  and g5606__2883(n_1674 ,n_1609 ,n_1608);
  or g5607__2346(n_1672 ,n_1576 ,n_1611);
  and g5608__1666(n_1671 ,n_1468 ,n_1605);
  and g5609__7410(n_1670 ,n_1603 ,n_1604);
  and g5610__6417(n_1669 ,n_1600 ,n_1599);
  and g5611__5477(n_1668 ,n_1560 ,n_1628);
  and g5612__2398(n_1667 ,n_1586 ,n_1585);
  not g5613(n_1660 ,n_1659);
  not g5614(n_1658 ,n_1657);
  not g5617(n_1650 ,n_1649);
  not g5618(n_1646 ,n_1645);
  and g5619__5107(n_1644 ,n_981 ,n_1597);
  nor g5620__6260(n_1643 ,n_1139 ,n_1598);
  nor g5621__4319(n_1642 ,n_1154 ,n_1598);
  nor g5622__8428(n_1641 ,n_1136 ,n_1594);
  and g5623__5526(n_1815 ,n_1054 ,n_1591);
  nor g5624__6783(n_1640 ,n_1054 ,n_1596);
  and g5625__3680(n_1639 ,in5[4] ,n_1589);
  and g5626__1617(n_1638 ,in5[4] ,n_1588);
  and g5627__2802(n_1637 ,in5[4] ,n_1590);
  nor g5628__1705(n_1636 ,n_991 ,n_1592);
  nor g5629__5122(n_1635 ,n_1115 ,n_1593);
  nor g5630__8246(n_1634 ,n_1262 ,n_1593);
  and g5631__7098(n_1662 ,n_1582 ,n_1581);
  and g5632__6131(n_1661 ,n_1612 ,n_1565);
  or g5633__1881(n_1659 ,n_1517 ,n_1615);
  or g5634__5115(n_1657 ,n_1403 ,n_1601);
  or g5635__7482(n_1656 ,n_1566 ,n_1567);
  and g5636__4733(n_1655 ,n_1570 ,n_1568);
  and g5637__6161(n_1654 ,n_1514 ,n_1572);
  and g5638__9315(n_1653 ,n_1574 ,n_1573);
  and g5639__9945(n_1652 ,n_957 ,n_1595);
  and g5640__2883(n_1651 ,n_1563 ,n_1587);
  or g5641__2346(n_1649 ,n_1515 ,n_1577);
  and g5642__1666(n_1648 ,n_1579 ,n_1578);
  or g5643__7410(n_1647 ,n_1445 ,n_1580);
  and g5644__6417(n_1645 ,n_1402 ,n_1584);
  or g5645__5477(n_1631 ,n_938 ,n_1559);
  or g5646__2398(n_1630 ,n_1098 ,n_1540);
  or g5647__5107(n_1629 ,n_938 ,n_1558);
  or g5648__6260(n_1628 ,n_938 ,n_1528);
  or g5649__4319(n_1627 ,in5[3] ,n_1556);
  and g5650__8428(n_1626 ,in5[3] ,n_1557);
  or g5651__5526(n_1625 ,n_1098 ,n_1531);
  or g5652__6783(n_1624 ,in5[3] ,n_1552);
  or g5653__3680(n_1623 ,in5[3] ,n_1530);
  or g5654__1617(n_1622 ,n_1098 ,n_1554);
  and g5655__2802(n_1621 ,in5[3] ,n_1536);
  nor g5656__1705(n_1620 ,in5[3] ,n_1539);
  and g5657__5122(n_1619 ,in5[5] ,n_1527);
  or g5658__8246(n_1618 ,in5[3] ,n_1538);
  or g5659__7098(n_1617 ,n_1098 ,n_1553);
  nor g5660__6131(n_1616 ,in5[3] ,n_1551);
  and g5661__1881(n_1814 ,n_1054 ,n_1527);
  nor g5662__5115(n_1615 ,in5[3] ,n_1549);
  and g5663__7482(n_1614 ,in5[3] ,n_1522);
  or g5664__4733(n_1613 ,in5[3] ,n_1547);
  or g5665__6161(n_1612 ,n_1098 ,n_1545);
  nor g5666__9315(n_1611 ,in5[3] ,n_1555);
  or g5667__9945(n_1610 ,in5[3] ,n_1545);
  or g5668__2883(n_1609 ,n_1098 ,n_1544);
  or g5669__2346(n_1608 ,in5[3] ,n_1542);
  or g5670__1666(n_1607 ,n_1098 ,n_1543);
  or g5671__7410(n_1606 ,in5[3] ,n_1534);
  or g5672__6417(n_1605 ,in5[3] ,n_1540);
  or g5673__5477(n_1604 ,in5[3] ,n_1523);
  or g5674__2398(n_1603 ,n_1098 ,n_1538);
  or g5675__5107(n_1602 ,in5[3] ,n_1532);
  nor g5676__6260(n_1601 ,in5[3] ,n_1531);
  or g5677__4319(n_1600 ,n_1098 ,n_1530);
  or g5678__8428(n_1599 ,in5[3] ,n_1528);
  or g5679__5526(n_1633 ,n_938 ,n_1534);
  or g5680__6783(n_1632 ,n_1098 ,n_1546);
  not g5681(n_1597 ,n_1596);
  not g5682(n_1595 ,n_1594);
  not g5683(n_1592 ,n_1591);
  or g5684__3680(n_1587 ,in5[3] ,n_1537);
  or g5685__1617(n_1586 ,n_1098 ,n_1555);
  or g5686__2802(n_1585 ,in5[3] ,n_1554);
  or g5687__1705(n_1584 ,n_1098 ,n_1532);
  nor g5688__5122(n_1583 ,n_1154 ,n_1526);
  or g5689__8246(n_1582 ,n_938 ,n_1551);
  or g5690__7098(n_1581 ,in5[3] ,n_1543);
  nor g5691__6131(n_1580 ,n_1098 ,n_1556);
  or g5692__1881(n_1579 ,n_1098 ,n_1537);
  or g5693__5115(n_1578 ,in5[3] ,n_1558);
  nor g5694__7482(n_1577 ,n_1098 ,n_1552);
  and g5695__4733(n_1576 ,in5[3] ,n_1548);
  nor g5696__6161(n_1575 ,n_1119 ,n_1526);
  or g5697__9315(n_1574 ,n_1098 ,n_1539);
  or g5698__9945(n_1573 ,in5[3] ,n_1553);
  or g5699__2883(n_1572 ,n_938 ,n_1547);
  nor g5700__2346(n_1571 ,n_1068 ,n_1533);
  or g5701__1666(n_1570 ,n_1098 ,n_1549);
  nor g5702__7410(n_1569 ,in5[3] ,n_1541);
  or g5703__6417(n_1568 ,in5[3] ,n_1559);
  nor g5704__5477(n_1567 ,n_1098 ,n_1542);
  nor g5705__2398(n_1566 ,in5[3] ,n_1546);
  or g5706__5107(n_1565 ,in5[3] ,n_1544);
  nor g5707__6260(n_1564 ,n_1108 ,n_1524);
  or g5708__4319(n_1563 ,n_938 ,n_1529);
  nor g5709__8428(n_1562 ,n_1138 ,n_1550);
  nor g5710__5526(n_1561 ,n_1154 ,n_1550);
  or g5711__6783(n_1560 ,in5[3] ,n_1535);
  or g5712__3680(n_1598 ,n_1098 ,n_1541);
  or g5713__1617(n_1596 ,in5[4] ,n_1533);
  or g5714__2802(n_1594 ,in5[3] ,n_1529);
  or g5715__1705(n_1593 ,n_938 ,n_1535);
  and g5716__5122(n_1591 ,n_1068 ,n_1525);
  and g5717__8246(n_1590 ,n_1098 ,n_1548);
  and g5718__7098(n_1589 ,n_1098 ,n_1536);
  and g5719__6131(n_1588 ,n_938 ,n_1557);
  and g5720__1881(n_1559 ,n_1485 ,n_1484);
  and g5721__5115(n_1558 ,n_1501 ,n_1507);
  or g5722__7482(n_1557 ,n_1446 ,n_1500);
  and g5723__4733(n_1556 ,n_1506 ,n_1504);
  and g5724__6161(n_1555 ,n_1487 ,n_1452);
  and g5725__9315(n_1554 ,n_1505 ,n_1479);
  and g5726__9945(n_1553 ,n_1497 ,n_1496);
  and g5727__2883(n_1552 ,n_1495 ,n_1493);
  and g5728__2346(n_1551 ,n_1492 ,n_1483);
  or g5729__1666(n_1550 ,n_1098 ,n_1512);
  and g5730__7410(n_1549 ,n_1486 ,n_1488);
  or g5731__6417(n_1548 ,n_1490 ,n_1458);
  and g5732__5477(n_1547 ,n_1482 ,n_1481);
  and g5733__2398(n_1546 ,n_1348 ,n_1480);
  and g5734__5107(n_1545 ,n_1489 ,n_1491);
  and g5735__6260(n_1544 ,n_1511 ,n_1450);
  and g5736__4319(n_1543 ,n_1470 ,n_1465);
  and g5737__8428(n_1542 ,n_1447 ,n_1471);
  and g5738__5526(n_1541 ,n_1405 ,n_1469);
  and g5739__6783(n_1540 ,n_1466 ,n_1467);
  and g5740__3680(n_1539 ,n_1494 ,n_1499);
  and g5741__1617(n_1538 ,n_1464 ,n_1459);
  not g5742(n_1525 ,n_1524);
  not g5743(n_1523 ,n_1522);
  nor g5745__2802(n_1521 ,n_1154 ,n_1477);
  nor g5746__1705(n_1520 ,n_1138 ,n_1477);
  and g5747__5122(n_1519 ,n_1054 ,n_1475);
  nor g5748__8246(n_1518 ,n_1068 ,n_1473);
  nor g5749__7098(n_1517 ,n_1098 ,n_1513);
  or g5750__6131(n_1516 ,n_1098 ,n_1478);
  nor g5751__1881(n_1515 ,in5[3] ,n_1476);
  or g5752__5115(n_1514 ,in5[3] ,n_1512);
  and g5753__7482(n_1537 ,n_1449 ,n_1448);
  or g5754__4733(n_1536 ,n_1343 ,n_1503);
  and g5755__6161(n_1535 ,n_1472 ,n_1460);
  and g5756__9315(n_1534 ,n_1457 ,n_1463);
  or g5757__9945(n_1533 ,in5[3] ,n_1513);
  and g5758__2883(n_1532 ,n_1456 ,n_1454);
  and g5759__2346(n_1531 ,n_1502 ,n_1498);
  and g5760__1666(n_1530 ,n_1508 ,n_1455);
  and g5761__7410(n_1529 ,n_1404 ,n_1451);
  and g5762__6417(n_1528 ,n_1453 ,n_1510);
  and g5763__5477(n_1527 ,n_1108 ,n_1474);
  or g5764__2398(n_1526 ,n_938 ,n_1476);
  or g5765__5107(n_1524 ,in5[3] ,n_1478);
  or g5766__6260(n_1522 ,n_1462 ,n_1461);
  or g5767__4319(n_1511 ,n_1045 ,n_1427);
  or g5768__8428(n_1510 ,in5[2] ,n_1441);
  nor g5769__5526(n_1509 ,n_1136 ,n_1411);
  or g5770__6783(n_1508 ,n_930 ,n_1434);
  or g5771__3680(n_1507 ,in5[2] ,n_1440);
  or g5772__1617(n_1506 ,n_1045 ,n_1439);
  or g5773__2802(n_1505 ,n_1045 ,n_1436);
  or g5774__1705(n_1504 ,in5[2] ,n_1430);
  nor g5775__5122(n_1503 ,in5[2] ,n_1435);
  or g5776__8246(n_1502 ,n_1045 ,n_1435);
  or g5777__7098(n_1501 ,n_1045 ,n_1437);
  nor g5778__6131(n_1500 ,in5[2] ,n_1417);
  or g5779__1881(n_1499 ,in5[2] ,n_1434);
  or g5780__5115(n_1498 ,in5[2] ,n_1428);
  or g5781__7482(n_1497 ,n_1045 ,n_1431);
  or g5782__4733(n_1496 ,in5[2] ,n_1442);
  or g5783__6161(n_1495 ,n_1045 ,n_1441);
  or g5784__9315(n_1494 ,n_1045 ,n_1428);
  or g5785__9945(n_1493 ,in5[2] ,n_1406);
  or g5786__2883(n_1492 ,n_1045 ,n_1407);
  or g5787__2346(n_1491 ,in5[2] ,n_1407);
  and g5788__1666(n_1490 ,in5[2] ,n_1422);
  or g5789__7410(n_1489 ,n_1045 ,n_1417);
  or g5790__6417(n_1488 ,in5[2] ,n_1426);
  or g5791__5477(n_1487 ,n_1045 ,n_1426);
  or g5792__2398(n_1486 ,n_1045 ,n_1419);
  or g5793__5107(n_1485 ,n_1045 ,n_1416);
  or g5794__6260(n_1484 ,in5[2] ,n_1436);
  or g5795__4319(n_1483 ,in5[2] ,n_1427);
  or g5796__8428(n_1482 ,n_1045 ,n_1424);
  or g5797__5526(n_1481 ,in5[2] ,n_1438);
  or g5798__6783(n_1480 ,n_1045 ,n_1420);
  or g5799__3680(n_1479 ,in5[2] ,n_1424);
  or g5800__1617(n_1513 ,in5[2] ,n_1423);
  or g5801__2802(n_1512 ,n_930 ,n_1415);
  not g5803(n_1474 ,n_1473);
  or g5804__1705(n_1472 ,in5[2] ,n_1429);
  or g5805__5122(n_1471 ,in5[2] ,n_1409);
  or g5806__8246(n_1470 ,n_930 ,n_1414);
  or g5807__7098(n_1469 ,n_1045 ,n_1430);
  or g5808__6131(n_1468 ,n_938 ,n_1412);
  or g5809__1881(n_1467 ,in5[2] ,n_1418);
  or g5810__5115(n_1466 ,n_1045 ,n_1432);
  or g5811__7482(n_1465 ,in5[2] ,n_1421);
  or g5812__4733(n_1464 ,n_1045 ,n_1433);
  or g5813__6161(n_1463 ,in5[2] ,n_1415);
  nor g5814__9315(n_1462 ,n_1045 ,n_1440);
  nor g5815__9945(n_1461 ,in5[2] ,n_1439);
  or g5816__2883(n_1460 ,n_1045 ,n_1406);
  or g5817__2346(n_1459 ,in5[2] ,n_1437);
  nor g5818__1666(n_1458 ,in5[2] ,n_1419);
  or g5819__7410(n_1457 ,n_1045 ,n_1438);
  or g5820__6417(n_1456 ,n_1045 ,n_1409);
  or g5821__5477(n_1455 ,in5[2] ,n_1431);
  or g5822__2398(n_1454 ,in5[2] ,n_1420);
  or g5823__5107(n_1453 ,n_1045 ,n_1442);
  or g5824__6260(n_1452 ,in5[2] ,n_1416);
  or g5825__4319(n_1451 ,in5[2] ,n_1432);
  or g5826__8428(n_1450 ,in5[2] ,n_1414);
  or g5827__5526(n_1449 ,n_1045 ,n_1418);
  or g5828__6783(n_1448 ,in5[2] ,n_1433);
  or g5829__3680(n_1447 ,n_1045 ,n_1421);
  nor g5830__1617(n_1446 ,n_1045 ,n_1408);
  nor g5831__2802(n_1445 ,in5[3] ,n_1425);
  nor g5832__1705(n_1444 ,n_1139 ,n_1413);
  nor g5833__5122(n_1443 ,n_1154 ,n_1413);
  or g5834__8246(n_1478 ,in5[2] ,n_1408);
  or g5835__7098(n_1477 ,n_938 ,n_1425);
  or g5836__6131(n_1476 ,n_1045 ,n_1429);
  and g5837__1881(n_1475 ,n_957 ,n_1410);
  or g5838__5115(n_1473 ,in5[3] ,n_1412);
  and g5839__7482(n_1442 ,n_1392 ,n_1380);
  and g5840__4733(n_1441 ,n_1397 ,n_1335);
  and g5841__6161(n_1440 ,n_1389 ,n_1357);
  and g5842__9315(n_1439 ,n_1393 ,n_1352);
  and g5843__9945(n_1438 ,n_1340 ,n_1345);
  and g5844__2883(n_1437 ,n_1384 ,n_1377);
  and g5845__2346(n_1436 ,n_1341 ,n_1349);
  and g5846__1666(n_1435 ,n_1383 ,n_1398);
  and g5847__7410(n_1434 ,n_1374 ,n_1353);
  and g5848__6417(n_1433 ,n_1371 ,n_1368);
  and g5849__5477(n_1432 ,n_1338 ,n_1369);
  and g5850__2398(n_1431 ,n_1378 ,n_1396);
  and g5851__5107(n_1430 ,n_1346 ,n_1388);
  and g5852__6260(n_1429 ,n_1316 ,n_1375);
  and g5853__4319(n_1428 ,n_1390 ,n_1354);
  and g5854__8428(n_1427 ,n_1381 ,n_1362);
  and g5855__5526(n_1426 ,n_1364 ,n_1355);
  or g5856__6783(n_1425 ,n_930 ,n_1399);
  and g5857__3680(n_1424 ,n_1382 ,n_1360);
  not g5858(n_1423 ,n_1422);
  not g5859(n_1411 ,n_1410);
  or g5860__1617(n_1405 ,in5[2] ,n_1399);
  or g5861__2802(n_1404 ,n_1045 ,n_1366);
  nor g5862__1705(n_1403 ,n_1098 ,n_1400);
  or g5863__5122(n_1402 ,in5[3] ,n_1367);
  or g5864__8246(n_1422 ,n_1347 ,n_1351);
  and g5865__7098(n_1421 ,n_1356 ,n_1337);
  and g5866__6131(n_1420 ,n_1365 ,n_1344);
  and g5867__1881(n_1419 ,n_1342 ,n_1395);
  and g5868__5115(n_1418 ,n_1359 ,n_1387);
  and g5869__7482(n_1417 ,n_1373 ,n_1379);
  and g5870__4733(n_1416 ,n_1385 ,n_1386);
  and g5871__6161(n_1415 ,n_1391 ,n_1336);
  and g5872__9315(n_1414 ,n_1361 ,n_1358);
  or g5873__9945(n_1413 ,n_938 ,n_1367);
  or g5874__2883(n_1412 ,in5[2] ,n_1366);
  and g5875__2346(n_1410 ,n_938 ,n_1401);
  and g5876__1666(n_1409 ,n_1394 ,n_1350);
  and g5877__7410(n_1408 ,n_1317 ,n_1363);
  and g5878__6417(n_1407 ,n_1372 ,n_1370);
  and g5879__5477(n_1406 ,n_1376 ,n_1339);
  not g5880(n_1401 ,n_1400);
  or g5881__2398(n_1398 ,in5[1] ,n_1322);
  or g5882__5107(n_1397 ,n_1030 ,n_1313);
  or g5883__6260(n_1396 ,in5[1] ,n_1298);
  or g5884__4319(n_1395 ,in5[1] ,n_1324);
  or g5885__8428(n_1394 ,n_1030 ,n_1325);
  or g5886__5526(n_1393 ,n_1030 ,n_1305);
  or g5887__6783(n_1392 ,n_1030 ,n_1320);
  or g5888__3680(n_1391 ,n_1030 ,n_1327);
  or g5889__1617(n_1390 ,n_1030 ,n_1303);
  or g5890__2802(n_1389 ,n_1030 ,n_1308);
  or g5891__1705(n_1388 ,in5[1] ,n_1327);
  or g5892__5122(n_1387 ,in5[1] ,n_1312);
  or g5893__8246(n_1386 ,in5[1] ,n_1326);
  or g5894__7098(n_1385 ,n_1030 ,n_1330);
  or g5895__6131(n_1384 ,n_1030 ,n_1326);
  or g5896__1881(n_1383 ,n_1030 ,n_1309);
  or g5897__5115(n_1382 ,n_1030 ,n_1323);
  or g5898__7482(n_1381 ,n_1030 ,n_1334);
  or g5899__4733(n_1380 ,in5[1] ,n_1300);
  or g5900__6161(n_1379 ,in5[1] ,n_1303);
  or g5901__9315(n_1378 ,n_1030 ,n_1314);
  or g5902__9945(n_1377 ,in5[1] ,n_1321);
  or g5903__2883(n_1376 ,n_1030 ,n_1306);
  or g5904__2346(n_1375 ,n_1030 ,n_1301);
  or g5905__1666(n_1374 ,n_1030 ,n_1319);
  or g5906__7410(n_1373 ,n_950 ,n_1322);
  or g5907__6417(n_1372 ,n_1030 ,n_1307);
  or g5908__5477(n_1371 ,n_1030 ,n_1318);
  or g5909__2398(n_1370 ,in5[1] ,n_1319);
  or g5910__5107(n_1369 ,in5[1] ,n_1310);
  or g5911__6260(n_1368 ,in5[1] ,n_1330);
  or g5912__4319(n_1400 ,in5[2] ,n_1331);
  or g5913__8428(n_1399 ,n_1030 ,n_1299);
  or g5914__5526(n_1365 ,n_1030 ,n_1302);
  or g5915__6783(n_1364 ,n_1030 ,n_1312);
  or g5916__3680(n_1363 ,in5[1] ,n_1309);
  or g5917__1617(n_1362 ,in5[1] ,n_1314);
  or g5918__2802(n_1361 ,n_1030 ,n_1298);
  or g5919__1705(n_1360 ,in5[1] ,n_1305);
  or g5920__5122(n_1359 ,n_1030 ,n_1324);
  or g5921__8246(n_1358 ,in5[1] ,n_1320);
  or g5922__7098(n_1357 ,in5[1] ,n_1323);
  or g5923__6131(n_1356 ,n_1030 ,n_1300);
  or g5924__1881(n_1355 ,in5[1] ,n_1318);
  or g5925__5115(n_1354 ,in5[1] ,n_1307);
  or g5926__7482(n_1353 ,in5[1] ,n_1334);
  or g5927__4733(n_1352 ,in5[1] ,n_1315);
  and g5928__6161(n_1351 ,n_1030 ,n_1332);
  or g5929__9315(n_1350 ,in5[1] ,n_1306);
  or g5930__9945(n_1349 ,in5[1] ,n_1308);
  or g5931__2883(n_1348 ,in5[2] ,n_1311);
  and g5932__2346(n_1347 ,in5[1] ,n_1328);
  or g5933__1666(n_1346 ,n_1030 ,n_1304);
  or g5934__7410(n_1345 ,in5[1] ,n_1304);
  or g5935__6417(n_1344 ,in5[1] ,n_1301);
  nor g5936__5477(n_1343 ,n_1045 ,n_1331);
  or g5937__2398(n_1342 ,n_1030 ,n_1310);
  or g5938__5107(n_1341 ,n_1030 ,n_1321);
  or g5939__6260(n_1340 ,n_1030 ,n_1315);
  or g5940__4319(n_1339 ,in5[1] ,n_1302);
  or g5941__8428(n_1338 ,n_1030 ,n_1333);
  or g5942__5526(n_1337 ,in5[1] ,n_1313);
  or g5943__6783(n_1336 ,in5[1] ,n_1299);
  or g5944__3680(n_1335 ,in5[1] ,n_1325);
  or g5945__1617(n_1367 ,n_1045 ,n_1311);
  or g5946__2802(n_1366 ,in5[1] ,n_1329);
  not g5947(n_1333 ,n_1332);
  not g5948(n_1329 ,n_1328);
  or g5949__1705(n_1317 ,n_1030 ,n_1297);
  or g5950__5122(n_1316 ,in5[1] ,n_1264);
  and g5951__8246(n_1334 ,n_1255 ,n_1294);
  or g5952__7098(n_1332 ,n_1244 ,n_1277);
  or g5953__6131(n_1331 ,in5[1] ,n_1297);
  and g5954__1881(n_1330 ,n_1257 ,n_1286);
  or g5955__5115(n_1328 ,n_1259 ,n_1287);
  and g5956__7482(n_1327 ,n_1239 ,n_1269);
  and g5957__4733(n_1326 ,n_1243 ,n_1291);
  and g5958__6161(n_1325 ,n_1241 ,n_1267);
  and g5959__9315(n_1324 ,n_1242 ,n_1274);
  and g5960__9945(n_1323 ,n_1230 ,n_1265);
  and g5961__2883(n_1322 ,n_1233 ,n_1288);
  and g5962__2346(n_1321 ,n_1238 ,n_1278);
  and g5963__1666(n_1320 ,n_1231 ,n_1268);
  and g5964__7410(n_1319 ,n_1252 ,n_1284);
  and g5965__6417(n_1318 ,n_1250 ,n_1282);
  and g5966__5477(n_1315 ,n_1232 ,n_1293);
  and g5967__2398(n_1314 ,n_1254 ,n_1295);
  and g5968__5107(n_1313 ,n_1256 ,n_1271);
  and g5969__6260(n_1312 ,n_1246 ,n_1289);
  or g5970__4319(n_1311 ,n_950 ,n_1264);
  and g5971__8428(n_1310 ,n_1253 ,n_1292);
  and g5972__5526(n_1309 ,n_1240 ,n_1290);
  and g5973__6783(n_1308 ,n_1247 ,n_1296);
  and g5974__3680(n_1307 ,n_1249 ,n_1281);
  and g5975__1617(n_1306 ,n_1235 ,n_1270);
  and g5976__2802(n_1305 ,n_1237 ,n_1276);
  and g5977__1705(n_1304 ,n_1280 ,n_1273);
  and g5978__5122(n_1303 ,n_1248 ,n_1279);
  and g5979__8246(n_1302 ,n_1251 ,n_1266);
  and g5980__7098(n_1301 ,n_1236 ,n_1272);
  and g5981__6131(n_1300 ,n_1245 ,n_1283);
  and g5982__1881(n_1299 ,n_1258 ,n_1285);
  and g5983__5115(n_1298 ,n_1234 ,n_1275);
  or g5984__7482(n_1296 ,n_1200 ,in5[0]);
  or g5985__4733(n_1295 ,n_1229 ,in5[0]);
  or g5986__6161(n_1294 ,n_1210 ,in5[0]);
  or g5987__9315(n_1293 ,n_1222 ,in5[0]);
  or g5988__9945(n_1292 ,n_1214 ,in5[0]);
  or g5989__2883(n_1291 ,n_1199 ,in5[0]);
  or g5990__2346(n_1290 ,n_1225 ,in5[0]);
  or g5991__1666(n_1289 ,n_1221 ,in5[0]);
  or g5992__7410(n_1288 ,n_1205 ,in5[0]);
  and g5993__6417(n_1287 ,in2[1] ,n_1039);
  or g5994__5477(n_1286 ,n_1203 ,in5[0]);
  or g5995__2398(n_1285 ,n_1213 ,in5[0]);
  or g5996__5107(n_1284 ,n_1208 ,in5[0]);
  or g5997__6260(n_1283 ,n_1204 ,in5[0]);
  or g5998__4319(n_1282 ,n_1207 ,in5[0]);
  or g5999__8428(n_1281 ,n_1206 ,in5[0]);
  or g6000__5526(n_1280 ,n_1227 ,n_1039);
  or g6001__6783(n_1279 ,n_1226 ,in5[0]);
  or g6002__3680(n_1278 ,n_1202 ,in5[0]);
  and g6003__1617(n_1277 ,in2[3] ,n_1039);
  or g6004__2802(n_1276 ,n_1215 ,in5[0]);
  or g6005__1705(n_1275 ,n_1223 ,in5[0]);
  or g6006__5122(n_1274 ,n_1228 ,in5[0]);
  or g6007__8246(n_1273 ,n_1201 ,in5[0]);
  or g6008__7098(n_1272 ,n_1224 ,in5[0]);
  or g6009__6131(n_1271 ,n_1217 ,in5[0]);
  or g6010__1881(n_1270 ,n_1227 ,in5[0]);
  or g6011__5115(n_1269 ,n_1197 ,in5[0]);
  or g6012__7482(n_1268 ,n_1219 ,in5[0]);
  or g6013__4733(n_1267 ,n_1218 ,in5[0]);
  or g6014__6161(n_1266 ,n_1216 ,in5[0]);
  or g6015__9315(n_1265 ,n_1220 ,in5[0]);
  or g6016__9945(n_1297 ,n_1209 ,in5[0]);
  not g6017(n_1263 ,n_1191);
  not g6022(n_1262 ,n_1133);
  nor g6028__2883(n_1259 ,n_1039 ,n_1209);
  or g6029__2346(n_1258 ,n_1224 ,n_1039);
  or g6030__1666(n_1257 ,n_1210 ,n_1039);
  or g6031__7410(n_1256 ,n_1220 ,n_1039);
  or g6032__6417(n_1255 ,n_1207 ,n_1039);
  or g6033__5477(n_1254 ,n_1203 ,n_1039);
  or g6034__2398(n_1253 ,n_1205 ,n_1039);
  or g6035__5107(n_1252 ,n_1221 ,n_1039);
  or g6036__6260(n_1251 ,n_1201 ,n_1039);
  or g6037__4319(n_1250 ,n_1208 ,n_1039);
  or g6038__8428(n_1249 ,n_1228 ,n_1039);
  or g6039__5526(n_1248 ,n_1214 ,n_1039);
  or g6040__6783(n_1247 ,n_1219 ,n_1039);
  or g6041__3680(n_1246 ,n_1206 ,n_948);
  or g6042__1617(n_1245 ,n_1200 ,n_948);
  nor g6043__2802(n_1244 ,n_1039 ,n_1225);
  or g6044__1705(n_1243 ,n_1229 ,n_1039);
  or g6045__5122(n_1242 ,n_1226 ,n_1039);
  or g6046__8246(n_1241 ,n_1215 ,n_1039);
  or g6047__7098(n_1240 ,n_1198 ,n_1039);
  or g6048__6131(n_1239 ,n_1216 ,n_1039);
  or g6049__1881(n_1238 ,n_1223 ,n_1039);
  or g6050__5115(n_1237 ,n_1217 ,n_1039);
  or g6051__7482(n_1236 ,n_1197 ,n_1039);
  or g6052__4733(n_1235 ,n_1222 ,n_1039);
  or g6053__6161(n_1234 ,n_1199 ,n_1039);
  or g6054__9315(n_1233 ,n_1196 ,n_1039);
  or g6055__9945(n_1232 ,n_1218 ,n_948);
  or g6056__2883(n_1231 ,n_1202 ,n_948);
  or g6057__2346(n_1230 ,n_1204 ,n_1039);
  or g6058__1666(n_1264 ,n_1213 ,n_1039);
  or g6059__7410(n_1191 ,in5[5] ,in5[4]);
  and g6060__6417(n_1261 ,in5[4] ,n_1054);
  not g6061(n_1229 ,in2[14]);
  not g6062(n_1228 ,in2[7]);
  not g6063(n_1227 ,in2[26]);
  not g6064(n_1226 ,in2[6]);
  not g6065(n_1225 ,in2[2]);
  not g6066(n_1224 ,in2[30]);
  not g6067(n_1223 ,in2[16]);
  not g6068(n_1222 ,in2[25]);
  not g6069(n_1221 ,in2[9]);
  not g6070(n_1220 ,in2[21]);
  not g6071(n_1219 ,in2[18]);
  not g6072(n_1218 ,in2[24]);
  not g6073(n_1217 ,in2[22]);
  not g6074(n_1216 ,in2[28]);
  not g6075(n_1215 ,in2[23]);
  not g6076(n_1214 ,in2[5]);
  not g6077(n_1213 ,in2[31]);
  not g6078(n_1212 ,in5[1]);
  not g6079(n_1211 ,in5[2]);
  not g6080(n_1210 ,in2[12]);
  not g6081(n_1209 ,in2[0]);
  not g6082(n_1208 ,in2[10]);
  not g6083(n_1207 ,in2[11]);
  not g6084(n_1206 ,in2[8]);
  not g6085(n_1205 ,in2[4]);
  not g6086(n_1204 ,in2[20]);
  not g6087(n_1203 ,in2[13]);
  not g6088(n_1202 ,in2[17]);
  not g6089(n_1201 ,in2[27]);
  not g6090(n_1200 ,in2[19]);
  not g6091(n_1199 ,in2[15]);
  not g6092(n_1198 ,in2[1]);
  not g6093(n_1197 ,in2[29]);
  not g6094(n_1196 ,in2[3]);
  not g6095(n_1195 ,in5[4]);
  not g6096(n_1194 ,in5[0]);
  not g6097(n_1193 ,in5[5]);
  not g6098(n_1192 ,in5[3]);
  not drc_bufs6099(n_1186 ,n_1064);
  not drc_bufs6100(n_1185 ,n_1063);
  not drc_bufs6103(n_1182 ,n_1064);
  not drc_bufs6106(n_1179 ,n_1193);
  not drc_bufs6113(n_1177 ,n_1124);
  not drc_bufs6121(n_1173 ,n_1130);
  not drc_bufs6129(n_1169 ,n_1126);
  not drc_bufs6137(n_1165 ,n_1128);
  not drc_bufs6172(n_1154 ,n_1152);
  not drc_bufs6174(n_1152 ,n_1262);
  not drc_bufs6192(n_1139 ,n_1137);
  not drc_bufs6193(n_1138 ,n_1137);
  not drc_bufs6194(n_1137 ,n_1191);
  buf drc_bufs6214(n_1817 ,n_1717);
  buf drc_bufs6215(n_1813 ,n_1519);
  buf drc_bufs6216(n_1816 ,n_1644);
  not drc_bufs6242(n_1136 ,n_1134);
  not drc_bufs6244(n_1134 ,n_1195);
  not drc_bufs6344(n_1133 ,n_1132);
  not drc_bufs6350(n_1132 ,n_1261);
  not drc_bufs6352(n_1130 ,n_1211);
  not drc_bufs6356(n_1128 ,n_1212);
  not drc_bufs6360(n_1126 ,n_1194);
  not drc_bufs6364(n_1124 ,n_1192);
  not drc_bufs6372(n_1119 ,n_1117);
  not drc_bufs6376(n_1117 ,n_1115);
  not drc_bufs6378(n_1115 ,n_1263);
  not drc_bufs6388(n_1109 ,n_1107);
  not drc_bufs6389(n_1108 ,n_1107);
  not drc_bufs6390(n_1107 ,n_1195);
  not drc_bufs6404(n_1098 ,n_1096);
  not drc_bufs6406(n_1096 ,n_1177);
  not drc_bufs6444(n_1068 ,n_1066);
  not drc_bufs6446(n_1066 ,n_1136);
  not drc_bufs6449(n_1064 ,n_1193);
  not drc_bufs6452(n_1063 ,n_1061);
  not drc_bufs6454(n_1061 ,n_1179);
  not drc_bufs6464(n_1054 ,n_1052);
  not drc_bufs6466(n_1052 ,n_1185);
  not drc_bufs6476(n_1045 ,n_1043);
  not drc_bufs6478(n_1043 ,n_1173);
  not drc_bufs6484(n_1039 ,n_1037);
  not drc_bufs6486(n_1037 ,n_1169);
  not drc_bufs6496(n_1030 ,n_1028);
  not drc_bufs6498(n_1028 ,n_1165);
  not drc_bufs6548(n_991 ,n_990);
  not drc_bufs6550(n_990 ,n_1186);
  not drc_bufs6565(n_981 ,n_980);
  not drc_bufs6566(n_980 ,n_1186);
  not drc_bufs6580(n_972 ,n_970);
  not drc_bufs6581(n_971 ,n_970);
  not drc_bufs6582(n_970 ,n_1182);
  not drc_bufs6597(n_962 ,n_961);
  not drc_bufs6598(n_961 ,n_1182);
  not drc_bufs6609(n_957 ,n_956);
  not drc_bufs6610(n_956 ,n_1109);
  not drc_bufs6620(n_950 ,n_949);
  not drc_bufs6622(n_949 ,n_1030);
  not drc_bufs6624(n_948 ,n_947);
  not drc_bufs6626(n_947 ,n_1039);
  not drc_bufs6644(n_938 ,n_937);
  not drc_bufs6646(n_937 ,n_1098);
  not drc_bufs6660(n_930 ,n_929);
  not drc_bufs6662(n_929 ,n_1045);
  and g2__5477(n_928 ,n_961 ,n_1777);
  and g6664__2398(n_927 ,n_1052 ,n_1776);
  and g6665__5107(n_926 ,n_1063 ,n_1775);
  and g6666__6260(n_925 ,n_990 ,n_1774);
  and g6667__4319(n_924 ,n_1052 ,n_1773);
  and g6668__8428(n_923 ,n_1052 ,n_1720);
  nor g6669__5526(n_922 ,n_1115 ,n_1654);
  and g6670__6783(n_921 ,n_1063 ,n_1652);
  and g6671__3680(n_920 ,n_980 ,n_1475);
  or g6672__1617(n_1938 ,n_600 ,n_902);
  or g6673__2802(n_1937 ,n_662 ,n_917);
  or g6674__1705(n_1925 ,n_832 ,n_918);
  or g6675__5122(n_1936 ,n_640 ,n_908);
  or g6676__8246(n_1935 ,n_746 ,n_905);
  or g6677__7098(n_1934 ,n_723 ,n_904);
  or g6678__6131(n_1939 ,n_523 ,n_919);
  or g6679__1881(n_1928 ,n_802 ,n_901);
  or g6680__5115(n_1932 ,n_743 ,n_7);
  or g6681__7482(n_1930 ,n_789 ,n_5);
  or g6682__4733(n_1929 ,n_773 ,n_898);
  or g6683__6161(n_1933 ,n_714 ,n_903);
  or g6684__9315(n_1927 ,n_784 ,n_4);
  or g6685__9945(n_1926 ,n_778 ,n_6);
  or g6686__2883(n_1931 ,n_774 ,n_8);
  and g6687__2346(n_1940 ,in4[5] ,n_891);
  and g6688__1666(n_919 ,in4[5] ,n_884);
  and g6689__7410(n_918 ,in4[5] ,n_885);
  or g6690__6417(n_1923 ,n_851 ,n_882);
  or g6691__5477(n_1921 ,n_849 ,n_880);
  or g6692__2398(n_1920 ,n_3 ,n_879);
  or g6693__5107(n_1918 ,n_847 ,n_881);
  and g6694__6260(n_917 ,in4[5] ,n_886);
  or g6695__4319(n_1916 ,n_812 ,n_863);
  or g6696__8428(n_1915 ,n_772 ,n_877);
  or g6697__5526(n_1914 ,n_808 ,n_876);
  or g6698__6783(n_1913 ,n_806 ,n_875);
  or g6699__3680(n_1911 ,n_801 ,n_874);
  or g6700__1617(n_1910 ,n_828 ,n_873);
  and g6701__2802(n_916 ,n_265 ,n_891);
  and g6702__1705(n_915 ,n_51 ,n_884);
  and g6703__5122(n_914 ,n_134 ,n_890);
  and g6704__8246(n_913 ,n_61 ,n_886);
  and g6705__7098(n_912 ,n_134 ,n_887);
  and g6706__6131(n_911 ,n_265 ,n_888);
  and g6707__1881(n_910 ,n_134 ,n_893);
  and g6708__5115(n_909 ,n_42 ,n_892);
  and g6709__7482(n_908 ,in4[5] ,n_887);
  and g6710__4733(n_907 ,n_134 ,n_889);
  and g6711__6161(n_906 ,n_265 ,n_885);
  and g6712__9315(n_905 ,in4[5] ,n_888);
  and g6713__9945(n_904 ,in4[5] ,n_893);
  and g6714__2883(n_903 ,in4[5] ,n_892);
  and g6715__2346(n_902 ,in4[5] ,n_890);
  and g6716__1666(n_901 ,in4[5] ,n_889);
  or g6717__7410(n_1924 ,n_830 ,n_852);
  or g6718__6417(n_1909 ,n_834 ,n_872);
  and g6719__5477(n_900 ,n_134 ,n_864);
  and g6720__2398(n_899 ,n_265 ,n_865);
  or g6721__5107(n_1912 ,n_2 ,n_862);
  nor g6722__6260(n_898 ,n_134 ,n_870);
  or g6723__4319(n_1917 ,n_853 ,n_883);
  or g6724__8428(n_1922 ,n_850 ,n_871);
  or g6725__5526(n_1919 ,n_848 ,n_878);
  and g6726__6783(n_897 ,n_134 ,n_867);
  and g6727__3680(n_896 ,n_71 ,n_869);
  and g6728__1617(n_895 ,n_134 ,n_866);
  and g6729__2802(n_894 ,n_265 ,n_868);
  or g6730__1705(n_883 ,n_715 ,n_813);
  or g6731__5122(n_882 ,n_524 ,n_826);
  or g6732__8246(n_881 ,n_724 ,n_814);
  or g6733__7098(n_880 ,n_654 ,n_823);
  or g6734__6131(n_879 ,n_641 ,n_820);
  or g6735__1881(n_878 ,n_744 ,n_817);
  or g6736__5115(n_877 ,n_809 ,n_810);
  or g6737__7482(n_876 ,n_1 ,n_807);
  or g6738__4733(n_875 ,n_816 ,n_777);
  or g6739__6161(n_874 ,n_716 ,n_827);
  or g6740__9315(n_873 ,n_699 ,n_781);
  or g6741__9945(n_872 ,n_0 ,n_775);
  or g6742__2883(n_871 ,n_599 ,n_825);
  or g6743__2346(n_893 ,n_794 ,n_793);
  or g6744__1666(n_892 ,n_779 ,n_792);
  or g6745__7410(n_891 ,n_822 ,n_821);
  or g6746__6417(n_890 ,n_787 ,n_829);
  or g6747__5477(n_889 ,n_650 ,n_785);
  or g6748__2398(n_888 ,n_796 ,n_795);
  or g6749__5107(n_887 ,n_780 ,n_797);
  or g6750__6260(n_886 ,n_815 ,n_819);
  or g6751__4319(n_885 ,n_589 ,n_831);
  or g6752__8428(n_884 ,n_818 ,n_798);
  not g6753(n_870 ,n_869);
  or g6754__5526(n_863 ,n_745 ,n_811);
  or g6755__6783(n_862 ,n_720 ,n_824);
  and g6756__3680(n_861 ,n_134 ,n_803);
  and g6757__1617(n_860 ,n_42 ,n_804);
  and g6758__2802(n_859 ,n_134 ,n_836);
  and g6759__1705(n_858 ,n_265 ,n_838);
  and g6760__5122(n_857 ,n_134 ,n_840);
  and g6761__8246(n_856 ,n_265 ,n_842);
  and g6762__7098(n_855 ,n_134 ,n_844);
  and g6763__6131(n_854 ,n_51 ,n_846);
  nor g6764__1881(n_853 ,n_265 ,n_805);
  nor g6765__5115(n_852 ,n_134 ,n_835);
  nor g6766__7482(n_851 ,n_134 ,n_837);
  nor g6767__4733(n_850 ,n_134 ,n_839);
  nor g6768__6161(n_849 ,n_265 ,n_841);
  nor g6769__9315(n_848 ,n_134 ,n_843);
  nor g6770__9945(n_847 ,n_52 ,n_845);
  or g6771__2883(n_869 ,n_719 ,n_786);
  or g6772__2346(n_868 ,n_718 ,n_790);
  or g6773__1666(n_867 ,n_717 ,n_791);
  or g6774__7410(n_866 ,n_598 ,n_833);
  or g6775__6417(n_865 ,n_722 ,n_788);
  or g6776__5477(n_864 ,n_643 ,n_782);
  not g6777(n_846 ,n_845);
  not g6778(n_844 ,n_843);
  not g6779(n_842 ,n_841);
  not g6780(n_840 ,n_839);
  not g6781(n_838 ,n_837);
  not g6782(n_836 ,n_835);
  nor g6783__2398(n_834 ,n_237 ,n_771);
  nor g6784__5107(n_833 ,in4[4] ,n_757);
  nor g6785__6260(n_832 ,n_237 ,n_748);
  nor g6786__4319(n_831 ,in4[4] ,n_771);
  nor g6787__8428(n_830 ,n_237 ,n_767);
  nor g6788__5526(n_829 ,in4[4] ,n_763);
  nor g6789__6783(n_828 ,n_237 ,n_757);
  and g6790__3680(n_827 ,n_197 ,n_736);
  nor g6791__1617(n_826 ,n_237 ,n_756);
  nor g6792__2802(n_825 ,n_237 ,n_763);
  nor g6793__1705(n_824 ,n_342 ,n_735);
  nor g6794__5122(n_823 ,n_342 ,n_759);
  and g6795__8246(n_822 ,in4[4] ,n_752);
  nor g6796__7098(n_821 ,in4[4] ,n_767);
  nor g6797__6131(n_820 ,n_237 ,n_758);
  nor g6798__1881(n_819 ,in4[4] ,n_759);
  and g6799__5115(n_818 ,in4[4] ,n_768);
  nor g6800__7482(n_817 ,n_237 ,n_754);
  and g6801__4733(n_816 ,in4[5] ,n_770);
  and g6802__6161(n_815 ,in4[4] ,n_765);
  nor g6803__9315(n_814 ,n_342 ,n_750);
  nor g6804__9945(n_813 ,n_237 ,n_749);
  and g6805__2883(n_812 ,in4[5] ,n_764);
  nor g6806__2346(n_811 ,n_237 ,n_747);
  nor g6807__1666(n_810 ,n_237 ,n_742);
  and g6808__7410(n_809 ,in4[5] ,n_762);
  and g6809__6417(n_808 ,n_197 ,n_727);
  nor g6810__5477(n_807 ,n_237 ,n_728);
  nor g6811__2398(n_806 ,n_237 ,n_733);
  or g6812__5107(n_845 ,in4[4] ,n_751);
  or g6813__6260(n_843 ,in4[4] ,n_755);
  or g6814__4319(n_841 ,in4[4] ,n_766);
  or g6815__8428(n_839 ,in4[4] ,n_731);
  or g6816__5526(n_837 ,in4[4] ,n_769);
  or g6817__6783(n_835 ,in4[4] ,n_753);
  not g6818(n_805 ,n_804);
  nor g6819__3680(n_802 ,n_237 ,n_734);
  nor g6820__1617(n_801 ,n_237 ,n_741);
  and g6821__2802(n_800 ,n_265 ,n_762);
  and g6822__1705(n_799 ,n_134 ,n_770);
  nor g6823__5122(n_798 ,in4[4] ,n_756);
  nor g6824__8246(n_797 ,in4[4] ,n_758);
  nor g6825__7098(n_796 ,n_216 ,n_755);
  nor g6826__6131(n_795 ,in4[4] ,n_754);
  nor g6827__1881(n_794 ,n_148 ,n_751);
  nor g6828__5115(n_793 ,in4[4] ,n_750);
  nor g6829__7482(n_792 ,in4[4] ,n_749);
  nor g6830__4733(n_791 ,in4[4] ,n_747);
  nor g6831__6161(n_790 ,in4[4] ,n_742);
  and g6832__9315(n_789 ,n_213 ,n_727);
  nor g6833__9945(n_788 ,in4[4] ,n_728);
  nor g6834__2883(n_787 ,n_148 ,n_731);
  nor g6835__2346(n_786 ,in4[4] ,n_733);
  nor g6836__1666(n_785 ,in4[4] ,n_735);
  and g6837__7410(n_784 ,n_213 ,n_736);
  and g6838__6417(n_783 ,n_265 ,n_764);
  nor g6839__5477(n_782 ,in4[4] ,n_741);
  and g6840__2398(n_781 ,n_197 ,n_760);
  nor g6841__5107(n_780 ,n_189 ,n_740);
  nor g6842__6260(n_779 ,n_148 ,n_738);
  nor g6843__4319(n_778 ,n_237 ,n_761);
  and g6844__8428(n_777 ,n_197 ,n_729);
  and g6845__5526(n_776 ,n_134 ,n_732);
  nor g6846__6783(n_775 ,n_195 ,n_748);
  nor g6847__3680(n_774 ,n_237 ,n_725);
  nor g6848__1617(n_773 ,n_237 ,n_730);
  and g6849__2802(n_772 ,n_197 ,n_726);
  and g6850__1705(n_804 ,n_148 ,n_737);
  and g6851__5122(n_803 ,n_148 ,n_739);
  not g6852(n_769 ,n_768);
  not g6853(n_766 ,n_765);
  not g6854(n_761 ,n_760);
  not g6855(n_753 ,n_752);
  nor g6856__8246(n_746 ,n_237 ,n_712);
  nor g6857__7098(n_745 ,n_195 ,n_713);
  nor g6858__6131(n_744 ,n_199 ,n_712);
  nor g6859__1881(n_743 ,n_237 ,n_713);
  and g6860__5115(n_771 ,n_705 ,n_703);
  and g6861__7482(n_770 ,n_148 ,n_668);
  or g6862__4733(n_768 ,n_706 ,n_696);
  and g6863__6161(n_767 ,n_702 ,n_685);
  or g6864__9315(n_765 ,n_701 ,n_700);
  and g6865__9945(n_764 ,n_148 ,n_669);
  and g6866__2883(n_763 ,n_709 ,n_707);
  and g6867__2346(n_762 ,n_148 ,n_667);
  or g6868__1666(n_760 ,n_648 ,n_693);
  and g6869__7410(n_759 ,n_697 ,n_704);
  and g6870__6417(n_758 ,n_711 ,n_692);
  and g6871__5477(n_757 ,n_710 ,n_698);
  and g6872__2398(n_756 ,n_686 ,n_681);
  and g6873__5107(n_755 ,n_596 ,n_689);
  and g6874__6260(n_754 ,n_688 ,n_687);
  or g6875__4319(n_752 ,n_655 ,n_690);
  and g6876__8428(n_751 ,n_548 ,n_684);
  and g6877__5526(n_750 ,n_682 ,n_683);
  and g6878__6783(n_749 ,n_679 ,n_678);
  and g6879__3680(n_748 ,n_639 ,n_708);
  and g6880__1617(n_747 ,n_665 ,n_664);
  not g6881(n_740 ,n_739);
  not g6882(n_738 ,n_737);
  not g6883(n_730 ,n_729);
  not g6884(n_726 ,n_725);
  and g6885__2802(n_1880 ,n_61 ,n_676);
  nor g6886__1705(n_724 ,n_219 ,n_677);
  nor g6887__5122(n_723 ,n_237 ,n_677);
  nor g6888__8246(n_722 ,n_216 ,n_673);
  and g6889__7098(n_721 ,n_134 ,n_670);
  nor g6890__6131(n_720 ,n_134 ,n_675);
  and g6891__1881(n_719 ,in4[4] ,n_668);
  and g6892__5115(n_718 ,in4[4] ,n_667);
  and g6893__7482(n_717 ,in4[4] ,n_669);
  nor g6894__4733(n_716 ,n_71 ,n_671);
  nor g6895__6161(n_715 ,n_195 ,n_672);
  nor g6896__9315(n_714 ,n_342 ,n_672);
  and g6897__9945(n_742 ,n_661 ,n_660);
  and g6898__2883(n_741 ,n_691 ,n_644);
  or g6899__2346(n_739 ,n_597 ,n_694);
  or g6900__1666(n_737 ,n_483 ,n_680);
  or g6901__7410(n_736 ,n_645 ,n_646);
  and g6902__6417(n_735 ,n_649 ,n_647);
  and g6903__5477(n_734 ,n_594 ,n_651);
  and g6904__2398(n_733 ,n_653 ,n_652);
  and g6905__5107(n_732 ,n_37 ,n_674);
  and g6906__6260(n_731 ,n_642 ,n_666);
  or g6907__4319(n_729 ,n_595 ,n_656);
  and g6908__8428(n_728 ,n_658 ,n_657);
  or g6909__5526(n_727 ,n_525 ,n_659);
  and g6910__6783(n_725 ,n_482 ,n_663);
  or g6911__3680(n_711 ,n_18 ,n_638);
  or g6912__1617(n_710 ,n_178 ,n_619);
  or g6913__2802(n_709 ,n_18 ,n_637);
  or g6914__1705(n_708 ,n_18 ,n_607);
  or g6915__5122(n_707 ,in4[3] ,n_635);
  and g6916__8246(n_706 ,in4[3] ,n_636);
  or g6917__7098(n_705 ,n_178 ,n_610);
  or g6918__6131(n_704 ,in4[3] ,n_631);
  or g6919__1881(n_703 ,in4[3] ,n_609);
  or g6920__5115(n_702 ,n_178 ,n_633);
  and g6921__7482(n_701 ,in4[3] ,n_615);
  nor g6922__4733(n_700 ,in4[3] ,n_618);
  and g6923__6161(n_699 ,in4[5] ,n_606);
  or g6924__9315(n_698 ,in4[3] ,n_617);
  or g6925__9945(n_697 ,n_178 ,n_632);
  nor g6926__2883(n_696 ,in4[3] ,n_630);
  and g6927__2346(n_695 ,n_134 ,n_606);
  nor g6928__1666(n_694 ,in4[3] ,n_628);
  and g6929__7410(n_693 ,in4[3] ,n_601);
  or g6930__6417(n_692 ,in4[3] ,n_626);
  or g6931__5477(n_691 ,n_178 ,n_624);
  nor g6932__2398(n_690 ,in4[3] ,n_634);
  or g6933__5107(n_689 ,in4[3] ,n_624);
  or g6934__6260(n_688 ,n_178 ,n_623);
  or g6935__4319(n_687 ,in4[3] ,n_621);
  or g6936__8428(n_686 ,n_178 ,n_622);
  or g6937__5526(n_685 ,in4[3] ,n_613);
  or g6938__6783(n_684 ,in4[3] ,n_619);
  or g6939__3680(n_683 ,in4[3] ,n_602);
  or g6940__1617(n_682 ,n_178 ,n_617);
  or g6941__2802(n_681 ,in4[3] ,n_611);
  nor g6942__1705(n_680 ,in4[3] ,n_610);
  or g6943__5122(n_679 ,n_178 ,n_609);
  or g6944__8246(n_678 ,in4[3] ,n_607);
  or g6945__7098(n_713 ,n_18 ,n_613);
  or g6946__6131(n_712 ,n_178 ,n_625);
  not g6947(n_676 ,n_675);
  not g6948(n_674 ,n_673);
  not g6949(n_671 ,n_670);
  or g6950__1881(n_666 ,in4[3] ,n_616);
  or g6951__5115(n_665 ,n_178 ,n_634);
  or g6952__7482(n_664 ,in4[3] ,n_633);
  or g6953__4733(n_663 ,n_178 ,n_611);
  nor g6954__6161(n_662 ,n_237 ,n_605);
  or g6955__9315(n_661 ,n_18 ,n_630);
  or g6956__9945(n_660 ,in4[3] ,n_622);
  nor g6957__2883(n_659 ,n_178 ,n_635);
  or g6958__2346(n_658 ,n_178 ,n_616);
  or g6959__1666(n_657 ,in4[3] ,n_637);
  nor g6960__7410(n_656 ,n_178 ,n_631);
  and g6961__6417(n_655 ,in4[3] ,n_627);
  nor g6962__5477(n_654 ,n_199 ,n_605);
  or g6963__2398(n_653 ,n_178 ,n_618);
  or g6964__5107(n_652 ,in4[3] ,n_632);
  or g6965__6260(n_651 ,n_18 ,n_626);
  nor g6966__4319(n_650 ,n_148 ,n_612);
  or g6967__8428(n_649 ,n_178 ,n_628);
  nor g6968__5526(n_648 ,in4[3] ,n_620);
  or g6969__6783(n_647 ,in4[3] ,n_638);
  nor g6970__3680(n_646 ,n_178 ,n_621);
  nor g6971__1617(n_645 ,in4[3] ,n_625);
  or g6972__2802(n_644 ,in4[3] ,n_623);
  nor g6973__1705(n_643 ,n_188 ,n_603);
  or g6974__5122(n_642 ,n_18 ,n_608);
  nor g6975__8246(n_641 ,n_218 ,n_629);
  nor g6976__7098(n_640 ,n_237 ,n_629);
  or g6977__6131(n_639 ,in4[3] ,n_614);
  or g6978__1881(n_677 ,n_178 ,n_620);
  or g6979__5115(n_675 ,in4[4] ,n_612);
  or g6980__7482(n_673 ,in4[3] ,n_608);
  or g6981__4733(n_672 ,n_18 ,n_614);
  and g6982__6161(n_670 ,n_148 ,n_604);
  and g6983__9315(n_669 ,n_178 ,n_627);
  and g6984__9945(n_668 ,n_178 ,n_615);
  and g6985__2883(n_667 ,n_18 ,n_636);
  and g6986__2346(n_638 ,n_565 ,n_564);
  and g6987__1666(n_637 ,n_581 ,n_587);
  or g6988__7410(n_636 ,n_526 ,n_580);
  and g6989__6417(n_635 ,n_586 ,n_584);
  and g6990__5477(n_634 ,n_567 ,n_532);
  and g6991__2398(n_633 ,n_585 ,n_559);
  and g6992__5107(n_632 ,n_577 ,n_576);
  and g6993__6260(n_631 ,n_575 ,n_573);
  and g6994__4319(n_630 ,n_572 ,n_563);
  or g6995__8428(n_629 ,n_178 ,n_592);
  and g6996__5526(n_628 ,n_566 ,n_568);
  or g6997__6783(n_627 ,n_570 ,n_538);
  and g6998__3680(n_626 ,n_562 ,n_561);
  and g6999__1617(n_625 ,n_428 ,n_560);
  and g7000__2802(n_624 ,n_569 ,n_571);
  and g7001__1705(n_623 ,n_591 ,n_530);
  and g7002__5122(n_622 ,n_550 ,n_545);
  and g7003__8246(n_621 ,n_527 ,n_551);
  and g7004__7098(n_620 ,n_485 ,n_549);
  and g7005__6131(n_619 ,n_546 ,n_547);
  and g7006__1881(n_618 ,n_574 ,n_579);
  and g7007__5115(n_617 ,n_544 ,n_539);
  not g7008(n_604 ,n_603);
  not g7009(n_602 ,n_601);
  nor g7010__7482(n_600 ,n_237 ,n_557);
  nor g7011__4733(n_599 ,n_218 ,n_557);
  and g7012__6161(n_1877 ,n_134 ,n_555);
  nor g7013__9315(n_598 ,n_148 ,n_553);
  nor g7014__9945(n_597 ,n_178 ,n_593);
  or g7015__2883(n_596 ,n_178 ,n_558);
  nor g7016__2346(n_595 ,in4[3] ,n_556);
  or g7017__1666(n_594 ,in4[3] ,n_592);
  and g7018__7410(n_616 ,n_529 ,n_528);
  or g7019__6417(n_615 ,n_423 ,n_583);
  and g7020__5477(n_614 ,n_552 ,n_540);
  and g7021__2398(n_613 ,n_537 ,n_543);
  or g7022__5107(n_612 ,in4[3] ,n_593);
  and g7023__6260(n_611 ,n_536 ,n_534);
  and g7024__4319(n_610 ,n_582 ,n_578);
  and g7025__8428(n_609 ,n_588 ,n_535);
  and g7026__5526(n_608 ,n_484 ,n_531);
  and g7027__6783(n_607 ,n_533 ,n_590);
  and g7028__3680(n_606 ,n_188 ,n_554);
  or g7029__1617(n_605 ,n_18 ,n_556);
  or g7030__2802(n_603 ,in4[3] ,n_558);
  or g7031__1705(n_601 ,n_542 ,n_541);
  or g7032__5122(n_591 ,n_125 ,n_507);
  or g7033__8246(n_590 ,in4[2] ,n_521);
  nor g7034__7098(n_589 ,n_216 ,n_491);
  or g7035__6131(n_588 ,n_10 ,n_514);
  or g7036__1881(n_587 ,in4[2] ,n_520);
  or g7037__5115(n_586 ,n_125 ,n_519);
  or g7038__7482(n_585 ,n_125 ,n_516);
  or g7039__4733(n_584 ,in4[2] ,n_510);
  nor g7040__6161(n_583 ,in4[2] ,n_515);
  or g7041__9315(n_582 ,n_125 ,n_515);
  or g7042__9945(n_581 ,n_125 ,n_517);
  nor g7043__2883(n_580 ,in4[2] ,n_497);
  or g7044__2346(n_579 ,in4[2] ,n_514);
  or g7045__1666(n_578 ,in4[2] ,n_508);
  or g7046__7410(n_577 ,n_125 ,n_511);
  or g7047__6417(n_576 ,in4[2] ,n_522);
  or g7048__5477(n_575 ,n_125 ,n_521);
  or g7049__2398(n_574 ,n_125 ,n_508);
  or g7050__5107(n_573 ,in4[2] ,n_486);
  or g7051__6260(n_572 ,n_125 ,n_487);
  or g7052__4319(n_571 ,in4[2] ,n_487);
  and g7053__8428(n_570 ,in4[2] ,n_502);
  or g7054__5526(n_569 ,n_125 ,n_497);
  or g7055__6783(n_568 ,in4[2] ,n_506);
  or g7056__3680(n_567 ,n_125 ,n_506);
  or g7057__1617(n_566 ,n_125 ,n_499);
  or g7058__2802(n_565 ,n_125 ,n_496);
  or g7059__1705(n_564 ,in4[2] ,n_516);
  or g7060__5122(n_563 ,in4[2] ,n_507);
  or g7061__8246(n_562 ,n_125 ,n_504);
  or g7062__7098(n_561 ,in4[2] ,n_518);
  or g7063__6131(n_560 ,n_125 ,n_500);
  or g7064__1881(n_559 ,in4[2] ,n_504);
  or g7065__5115(n_593 ,in4[2] ,n_503);
  or g7066__7482(n_592 ,n_10 ,n_495);
  not g7067(n_554 ,n_553);
  or g7068__4733(n_552 ,in4[2] ,n_509);
  or g7069__6161(n_551 ,in4[2] ,n_489);
  or g7070(n_550 ,n_10 ,n_494);
  or g7071(n_549 ,n_125 ,n_510);
  or g7072(n_548 ,n_18 ,n_492);
  or g7073(n_547 ,in4[2] ,n_498);
  or g7074(n_546 ,n_125 ,n_512);
  or g7075(n_545 ,in4[2] ,n_501);
  or g7076(n_544 ,n_125 ,n_513);
  or g7077(n_543 ,in4[2] ,n_495);
  nor g7078(n_542 ,n_125 ,n_520);
  nor g7079(n_541 ,in4[2] ,n_519);
  or g7080(n_540 ,n_125 ,n_486);
  or g7081(n_539 ,in4[2] ,n_517);
  nor g7082(n_538 ,in4[2] ,n_499);
  or g7083(n_537 ,n_125 ,n_518);
  or g7084(n_536 ,n_125 ,n_489);
  or g7085(n_535 ,in4[2] ,n_511);
  or g7086(n_534 ,in4[2] ,n_500);
  or g7087(n_533 ,n_125 ,n_522);
  or g7088(n_532 ,in4[2] ,n_496);
  or g7089(n_531 ,in4[2] ,n_512);
  or g7090(n_530 ,in4[2] ,n_494);
  or g7091(n_529 ,n_125 ,n_498);
  or g7092(n_528 ,in4[2] ,n_513);
  or g7093(n_527 ,n_125 ,n_501);
  nor g7094(n_526 ,n_125 ,n_488);
  nor g7095(n_525 ,in4[3] ,n_505);
  nor g7096(n_524 ,n_219 ,n_493);
  nor g7097(n_523 ,n_237 ,n_493);
  or g7098(n_558 ,in4[2] ,n_488);
  or g7099(n_557 ,n_18 ,n_505);
  or g7100(n_556 ,n_125 ,n_509);
  and g7101(n_555 ,n_37 ,n_490);
  or g7102(n_553 ,in4[3] ,n_492);
  and g7103(n_522 ,n_472 ,n_460);
  and g7104(n_521 ,n_477 ,n_415);
  and g7105(n_520 ,n_469 ,n_437);
  and g7106(n_519 ,n_473 ,n_432);
  and g7107(n_518 ,n_420 ,n_425);
  and g7108(n_517 ,n_464 ,n_457);
  and g7109(n_516 ,n_421 ,n_429);
  and g7110(n_515 ,n_463 ,n_478);
  and g7111(n_514 ,n_454 ,n_433);
  and g7112(n_513 ,n_451 ,n_448);
  and g7113(n_512 ,n_418 ,n_449);
  and g7114(n_511 ,n_458 ,n_476);
  and g7115(n_510 ,n_426 ,n_468);
  and g7116(n_509 ,n_396 ,n_455);
  and g7117(n_508 ,n_470 ,n_434);
  and g7118(n_507 ,n_461 ,n_442);
  and g7119(n_506 ,n_444 ,n_435);
  or g7120(n_505 ,n_10 ,n_479);
  and g7121(n_504 ,n_462 ,n_440);
  not g7122(n_503 ,n_502);
  not g7123(n_491 ,n_490);
  or g7124(n_485 ,in4[2] ,n_479);
  or g7125(n_484 ,n_125 ,n_446);
  nor g7126(n_483 ,n_178 ,n_480);
  or g7127(n_482 ,in4[3] ,n_447);
  or g7128(n_502 ,n_427 ,n_431);
  and g7129(n_501 ,n_436 ,n_417);
  and g7130(n_500 ,n_445 ,n_424);
  and g7131(n_499 ,n_422 ,n_475);
  and g7132(n_498 ,n_439 ,n_467);
  and g7133(n_497 ,n_453 ,n_459);
  and g7134(n_496 ,n_465 ,n_466);
  and g7135(n_495 ,n_471 ,n_416);
  and g7136(n_494 ,n_441 ,n_438);
  or g7137(n_493 ,n_18 ,n_447);
  or g7138(n_492 ,in4[2] ,n_446);
  and g7139(n_490 ,n_18 ,n_481);
  and g7140(n_489 ,n_474 ,n_430);
  and g7141(n_488 ,n_397 ,n_443);
  and g7142(n_487 ,n_452 ,n_450);
  and g7143(n_486 ,n_456 ,n_419);
  not g7144(n_481 ,n_480);
  or g7145(n_478 ,in4[1] ,n_402);
  or g7146(n_477 ,n_110 ,n_393);
  or g7147(n_476 ,in4[1] ,n_378);
  or g7148(n_475 ,in4[1] ,n_404);
  or g7149(n_474 ,n_110 ,n_405);
  or g7150(n_473 ,n_110 ,n_385);
  or g7151(n_472 ,n_110 ,n_400);
  or g7152(n_471 ,n_110 ,n_407);
  or g7153(n_470 ,n_110 ,n_383);
  or g7154(n_469 ,n_110 ,n_388);
  or g7155(n_468 ,in4[1] ,n_407);
  or g7156(n_467 ,in4[1] ,n_392);
  or g7157(n_466 ,in4[1] ,n_406);
  or g7158(n_465 ,n_110 ,n_410);
  or g7159(n_464 ,n_110 ,n_406);
  or g7160(n_463 ,n_110 ,n_389);
  or g7161(n_462 ,n_110 ,n_403);
  or g7162(n_461 ,n_110 ,n_414);
  or g7163(n_460 ,in4[1] ,n_380);
  or g7164(n_459 ,in4[1] ,n_383);
  or g7165(n_458 ,n_110 ,n_394);
  or g7166(n_457 ,in4[1] ,n_401);
  or g7167(n_456 ,n_110 ,n_386);
  or g7168(n_455 ,n_110 ,n_381);
  or g7169(n_454 ,n_110 ,n_399);
  or g7170(n_453 ,n_30 ,n_402);
  or g7171(n_452 ,n_110 ,n_387);
  or g7172(n_451 ,n_110 ,n_398);
  or g7173(n_450 ,in4[1] ,n_399);
  or g7174(n_449 ,in4[1] ,n_390);
  or g7175(n_448 ,in4[1] ,n_410);
  or g7176(n_480 ,in4[2] ,n_411);
  or g7177(n_479 ,n_110 ,n_379);
  or g7178(n_445 ,n_110 ,n_382);
  or g7179(n_444 ,n_110 ,n_392);
  or g7180(n_443 ,in4[1] ,n_389);
  or g7181(n_442 ,in4[1] ,n_394);
  or g7182(n_441 ,n_110 ,n_378);
  or g7183(n_440 ,in4[1] ,n_385);
  or g7184(n_439 ,n_110 ,n_404);
  or g7185(n_438 ,in4[1] ,n_400);
  or g7186(n_437 ,in4[1] ,n_403);
  or g7187(n_436 ,n_110 ,n_380);
  or g7188(n_435 ,in4[1] ,n_398);
  or g7189(n_434 ,in4[1] ,n_387);
  or g7190(n_433 ,in4[1] ,n_414);
  or g7191(n_432 ,in4[1] ,n_395);
  and g7192(n_431 ,n_110 ,n_412);
  or g7193(n_430 ,in4[1] ,n_386);
  or g7194(n_429 ,in4[1] ,n_388);
  or g7195(n_428 ,in4[2] ,n_391);
  and g7196(n_427 ,in4[1] ,n_408);
  or g7197(n_426 ,n_110 ,n_384);
  or g7198(n_425 ,in4[1] ,n_384);
  or g7199(n_424 ,in4[1] ,n_381);
  nor g7200(n_423 ,n_125 ,n_411);
  or g7201(n_422 ,n_110 ,n_390);
  or g7202(n_421 ,n_110 ,n_401);
  or g7203(n_420 ,n_110 ,n_395);
  or g7204(n_419 ,in4[1] ,n_382);
  or g7205(n_418 ,n_110 ,n_413);
  or g7206(n_417 ,in4[1] ,n_393);
  or g7207(n_416 ,in4[1] ,n_379);
  or g7208(n_415 ,in4[1] ,n_405);
  or g7209(n_447 ,n_125 ,n_391);
  or g7210(n_446 ,in4[1] ,n_409);
  not g7211(n_413 ,n_412);
  not g7212(n_409 ,n_408);
  or g7213(n_397 ,n_110 ,n_377);
  or g7214(n_396 ,in4[1] ,n_344);
  and g7215(n_414 ,n_335 ,n_374);
  or g7216(n_412 ,n_324 ,n_357);
  or g7217(n_411 ,in4[1] ,n_377);
  and g7218(n_410 ,n_337 ,n_366);
  or g7219(n_408 ,n_339 ,n_367);
  and g7220(n_407 ,n_319 ,n_349);
  and g7221(n_406 ,n_323 ,n_371);
  and g7222(n_405 ,n_321 ,n_347);
  and g7223(n_404 ,n_322 ,n_354);
  and g7224(n_403 ,n_310 ,n_345);
  and g7225(n_402 ,n_313 ,n_368);
  and g7226(n_401 ,n_318 ,n_358);
  and g7227(n_400 ,n_311 ,n_348);
  and g7228(n_399 ,n_332 ,n_364);
  and g7229(n_398 ,n_330 ,n_362);
  and g7230(n_395 ,n_312 ,n_373);
  and g7231(n_394 ,n_334 ,n_375);
  and g7232(n_393 ,n_336 ,n_351);
  and g7233(n_392 ,n_326 ,n_369);
  or g7234(n_391 ,n_30 ,n_344);
  and g7235(n_390 ,n_333 ,n_372);
  and g7236(n_389 ,n_320 ,n_370);
  and g7237(n_388 ,n_327 ,n_376);
  and g7238(n_387 ,n_329 ,n_361);
  and g7239(n_386 ,n_315 ,n_350);
  and g7240(n_385 ,n_317 ,n_356);
  and g7241(n_384 ,n_360 ,n_353);
  and g7242(n_383 ,n_328 ,n_359);
  and g7243(n_382 ,n_331 ,n_346);
  and g7244(n_381 ,n_316 ,n_352);
  and g7245(n_380 ,n_325 ,n_363);
  and g7246(n_379 ,n_338 ,n_365);
  and g7247(n_378 ,n_314 ,n_355);
  or g7248(n_376 ,n_280 ,in4[0]);
  or g7249(n_375 ,n_309 ,in4[0]);
  or g7250(n_374 ,n_290 ,in4[0]);
  or g7251(n_373 ,n_302 ,in4[0]);
  or g7252(n_372 ,n_294 ,in4[0]);
  or g7253(n_371 ,n_279 ,in4[0]);
  or g7254(n_370 ,n_305 ,in4[0]);
  or g7255(n_369 ,n_301 ,in4[0]);
  or g7256(n_368 ,n_285 ,in4[0]);
  and g7257(n_367 ,in1[1] ,n_119);
  or g7258(n_366 ,n_283 ,in4[0]);
  or g7259(n_365 ,n_293 ,in4[0]);
  or g7260(n_364 ,n_288 ,in4[0]);
  or g7261(n_363 ,n_284 ,in4[0]);
  or g7262(n_362 ,n_287 ,in4[0]);
  or g7263(n_361 ,n_286 ,in4[0]);
  or g7264(n_360 ,n_307 ,n_119);
  or g7265(n_359 ,n_306 ,in4[0]);
  or g7266(n_358 ,n_282 ,in4[0]);
  and g7267(n_357 ,in1[3] ,n_119);
  or g7268(n_356 ,n_295 ,in4[0]);
  or g7269(n_355 ,n_303 ,in4[0]);
  or g7270(n_354 ,n_308 ,in4[0]);
  or g7271(n_353 ,n_281 ,in4[0]);
  or g7272(n_352 ,n_304 ,in4[0]);
  or g7273(n_351 ,n_297 ,in4[0]);
  or g7274(n_350 ,n_307 ,in4[0]);
  or g7275(n_349 ,n_277 ,in4[0]);
  or g7276(n_348 ,n_299 ,in4[0]);
  or g7277(n_347 ,n_298 ,in4[0]);
  or g7278(n_346 ,n_296 ,in4[0]);
  or g7279(n_345 ,n_300 ,in4[0]);
  or g7280(n_377 ,n_289 ,in4[0]);
  not g7281(n_343 ,n_271);
  not g7282(n_342 ,n_213);
  nor g7286(n_339 ,n_119 ,n_289);
  or g7287(n_338 ,n_304 ,n_119);
  or g7288(n_337 ,n_290 ,n_119);
  or g7289(n_336 ,n_300 ,n_119);
  or g7290(n_335 ,n_287 ,n_119);
  or g7291(n_334 ,n_283 ,n_119);
  or g7292(n_333 ,n_285 ,n_119);
  or g7293(n_332 ,n_301 ,n_119);
  or g7294(n_331 ,n_281 ,n_119);
  or g7295(n_330 ,n_288 ,n_119);
  or g7296(n_329 ,n_308 ,n_119);
  or g7297(n_328 ,n_294 ,n_119);
  or g7298(n_327 ,n_299 ,n_119);
  or g7299(n_326 ,n_286 ,n_28);
  or g7300(n_325 ,n_280 ,n_28);
  nor g7301(n_324 ,n_119 ,n_305);
  or g7302(n_323 ,n_309 ,n_119);
  or g7303(n_322 ,n_306 ,n_119);
  or g7304(n_321 ,n_295 ,n_119);
  or g7305(n_320 ,n_278 ,n_119);
  or g7306(n_319 ,n_296 ,n_119);
  or g7307(n_318 ,n_303 ,n_119);
  or g7308(n_317 ,n_297 ,n_119);
  or g7309(n_316 ,n_277 ,n_119);
  or g7310(n_315 ,n_302 ,n_119);
  or g7311(n_314 ,n_279 ,n_119);
  or g7312(n_313 ,n_276 ,n_119);
  or g7313(n_312 ,n_298 ,n_28);
  or g7314(n_311 ,n_282 ,n_28);
  or g7315(n_310 ,n_284 ,n_119);
  or g7316(n_344 ,n_293 ,n_119);
  or g7317(n_271 ,in4[5] ,in4[4]);
  and g7318(n_341 ,in4[4] ,n_134);
  not g7319(n_309 ,in1[14]);
  not g7320(n_308 ,in1[7]);
  not g7321(n_307 ,in1[26]);
  not g7322(n_306 ,in1[6]);
  not g7323(n_305 ,in1[2]);
  not g7324(n_304 ,in1[30]);
  not g7325(n_303 ,in1[16]);
  not g7326(n_302 ,in1[25]);
  not g7327(n_301 ,in1[9]);
  not g7328(n_300 ,in1[21]);
  not g7329(n_299 ,in1[18]);
  not g7330(n_298 ,in1[24]);
  not g7331(n_297 ,in1[22]);
  not g7332(n_296 ,in1[28]);
  not g7333(n_295 ,in1[23]);
  not g7334(n_294 ,in1[5]);
  not g7335(n_293 ,in1[31]);
  not g7336(n_292 ,in4[1]);
  not g7337(n_291 ,in4[2]);
  not g7338(n_290 ,in1[12]);
  not g7339(n_289 ,in1[0]);
  not g7340(n_288 ,in1[10]);
  not g7341(n_287 ,in1[11]);
  not g7342(n_286 ,in1[8]);
  not g7343(n_285 ,in1[4]);
  not g7344(n_284 ,in1[20]);
  not g7345(n_283 ,in1[13]);
  not g7346(n_282 ,in1[17]);
  not g7347(n_281 ,in1[27]);
  not g7348(n_280 ,in1[19]);
  not g7349(n_279 ,in1[15]);
  not g7350(n_278 ,in1[1]);
  not g7351(n_277 ,in1[29]);
  not g7352(n_276 ,in1[3]);
  not g7353(n_275 ,in4[4]);
  not g7354(n_274 ,in4[0]);
  not g7355(n_273 ,in4[5]);
  not g7356(n_272 ,in4[3]);
  not drc_bufs7358(n_266 ,n_144);
  not drc_bufs7359(n_265 ,n_143);
  not drc_bufs7362(n_262 ,n_144);
  not drc_bufs7365(n_259 ,n_273);
  not drc_bufs7367(n_257 ,n_204);
  not drc_bufs7371(n_253 ,n_210);
  not drc_bufs7375(n_249 ,n_206);
  not drc_bufs7379(n_245 ,n_208);
  not drc_bufs7387(n_237 ,n_235);
  not drc_bufs7389(n_235 ,n_342);
  not drc_bufs7405(n_219 ,n_217);
  not drc_bufs7406(n_218 ,n_217);
  not drc_bufs7407(n_217 ,n_271);
  buf drc_bufs7408(n_1878 ,n_695);
  buf drc_bufs7409(n_1887 ,n_855);
  buf drc_bufs7410(n_1889 ,n_856);
  buf drc_bufs6217(n_1890 ,n_857);
  buf drc_bufs6218(n_1898 ,n_899);
  buf drc_bufs6219(n_1895 ,n_900);
  buf drc_bufs6220(n_1906 ,n_914);
  buf drc_bufs6221(n_1903 ,n_911);
  buf drc_bufs6222(n_1891 ,n_858);
  buf drc_bufs6223(n_1904 ,n_912);
  buf drc_bufs6224(n_1886 ,n_854);
  buf drc_bufs6225(n_1881 ,n_799);
  buf drc_bufs6226(n_1892 ,n_859);
  buf drc_bufs6227(n_1901 ,n_909);
  buf drc_bufs6228(n_1908 ,n_916);
  buf drc_bufs6229(n_1884 ,n_783);
  buf drc_bufs6230(n_1882 ,n_776);
  buf drc_bufs6231(n_1883 ,n_800);
  buf drc_bufs6232(n_1894 ,n_895);
  buf drc_bufs6233(n_1879 ,n_721);
  buf drc_bufs6234(n_1896 ,n_907);
  buf drc_bufs6235(n_1902 ,n_910);
  buf drc_bufs6236(n_1897 ,n_896);
  buf drc_bufs6237(n_1907 ,n_915);
  buf drc_bufs6238(n_1899 ,n_894);
  buf drc_bufs6239(n_1888 ,n_861);
  buf drc_bufs6240(n_1900 ,n_897);
  buf drc_bufs6241(n_1893 ,n_906);
  buf drc_bufs7411(n_1885 ,n_860);
  buf drc_bufs7412(n_1905 ,n_913);
  not drc_bufs6269(n_216 ,n_214);
  not drc_bufs6271(n_214 ,n_275);
  not drc_bufs6371(n_213 ,n_212);
  not drc_bufs7413(n_212 ,n_341);
  not drc_bufs6379(n_210 ,n_291);
  not drc_bufs6383(n_208 ,n_292);
  not drc_bufs6387(n_206 ,n_274);
  not drc_bufs6391(n_204 ,n_272);
  not drc_bufs6399(n_199 ,n_197);
  not drc_bufs6403(n_197 ,n_195);
  not drc_bufs7421(n_195 ,n_343);
  not drc_bufs6415(n_189 ,n_187);
  not drc_bufs7425(n_188 ,n_187);
  not drc_bufs7426(n_187 ,n_275);
  not drc_bufs6431(n_178 ,n_176);
  not drc_bufs7434(n_176 ,n_257);
  not drc_bufs6471(n_148 ,n_146);
  not drc_bufs7454(n_146 ,n_216);
  not drc_bufs7455(n_144 ,n_273);
  not drc_bufs6479(n_143 ,n_141);
  not drc_bufs7457(n_141 ,n_259);
  not drc_bufs6491(n_134 ,n_132);
  not drc_bufs7463(n_132 ,n_265);
  not drc_bufs6503(n_125 ,n_123);
  not drc_bufs7469(n_123 ,n_253);
  not drc_bufs6511(n_119 ,n_117);
  not drc_bufs7473(n_117 ,n_249);
  not drc_bufs6523(n_110 ,n_108);
  not drc_bufs7479(n_108 ,n_245);
  not drc_bufs6575(n_71 ,n_70);
  not drc_bufs7500(n_70 ,n_266);
  not drc_bufs6592(n_61 ,n_60);
  not drc_bufs7505(n_60 ,n_266);
  not drc_bufs6607(n_52 ,n_50);
  not drc_bufs6608(n_51 ,n_50);
  not drc_bufs7509(n_50 ,n_262);
  not drc_bufs7514(n_42 ,n_41);
  not drc_bufs6625(n_41 ,n_262);
  not drc_bufs7517(n_37 ,n_36);
  not drc_bufs6637(n_36 ,n_189);
  not drc_bufs6647(n_30 ,n_29);
  not drc_bufs6649(n_29 ,n_110);
  not drc_bufs6651(n_28 ,n_27);
  not drc_bufs6653(n_27 ,n_119);
  not drc_bufs6671(n_18 ,n_17);
  not drc_bufs6673(n_17 ,n_178);
  not drc_bufs6687(n_10 ,n_9);
  not drc_bufs6689(n_9 ,n_125);
  and g7519(n_8 ,n_41 ,n_868);
  and g7520(n_7 ,n_132 ,n_867);
  and g7521(n_6 ,n_143 ,n_866);
  and g7522(n_5 ,n_70 ,n_865);
  and g7523(n_4 ,n_132 ,n_864);
  and g7524(n_3 ,n_132 ,n_803);
  nor g7525(n_2 ,n_195 ,n_734);
  and g7526(n_1 ,n_143 ,n_732);
  and g7527(n_0 ,n_60 ,n_555);
  xnor csa_tree_add_8_49_groupi_g2217(out1[63] ,csa_tree_add_8_49_groupi_n_419 ,csa_tree_add_8_49_groupi_n_753);
  or csa_tree_add_8_49_groupi_g2218(csa_tree_add_8_49_groupi_n_753 ,csa_tree_add_8_49_groupi_n_336 ,csa_tree_add_8_49_groupi_n_751);
  xnor csa_tree_add_8_49_groupi_g2219(out1[62] ,csa_tree_add_8_49_groupi_n_750 ,csa_tree_add_8_49_groupi_n_438);
  and csa_tree_add_8_49_groupi_g2220(csa_tree_add_8_49_groupi_n_751 ,csa_tree_add_8_49_groupi_n_379 ,csa_tree_add_8_49_groupi_n_750);
  or csa_tree_add_8_49_groupi_g2221(csa_tree_add_8_49_groupi_n_750 ,csa_tree_add_8_49_groupi_n_333 ,csa_tree_add_8_49_groupi_n_748);
  xnor csa_tree_add_8_49_groupi_g2222(out1[61] ,csa_tree_add_8_49_groupi_n_747 ,csa_tree_add_8_49_groupi_n_437);
  and csa_tree_add_8_49_groupi_g2223(csa_tree_add_8_49_groupi_n_748 ,csa_tree_add_8_49_groupi_n_387 ,csa_tree_add_8_49_groupi_n_747);
  or csa_tree_add_8_49_groupi_g2224(csa_tree_add_8_49_groupi_n_747 ,csa_tree_add_8_49_groupi_n_378 ,csa_tree_add_8_49_groupi_n_745);
  xnor csa_tree_add_8_49_groupi_g2225(out1[60] ,csa_tree_add_8_49_groupi_n_744 ,csa_tree_add_8_49_groupi_n_436);
  and csa_tree_add_8_49_groupi_g2226(csa_tree_add_8_49_groupi_n_745 ,csa_tree_add_8_49_groupi_n_367 ,csa_tree_add_8_49_groupi_n_744);
  or csa_tree_add_8_49_groupi_g2227(csa_tree_add_8_49_groupi_n_744 ,csa_tree_add_8_49_groupi_n_386 ,csa_tree_add_8_49_groupi_n_742);
  xnor csa_tree_add_8_49_groupi_g2228(out1[59] ,csa_tree_add_8_49_groupi_n_741 ,csa_tree_add_8_49_groupi_n_435);
  and csa_tree_add_8_49_groupi_g2229(csa_tree_add_8_49_groupi_n_742 ,csa_tree_add_8_49_groupi_n_328 ,csa_tree_add_8_49_groupi_n_741);
  or csa_tree_add_8_49_groupi_g2230(csa_tree_add_8_49_groupi_n_741 ,csa_tree_add_8_49_groupi_n_319 ,csa_tree_add_8_49_groupi_n_739);
  xnor csa_tree_add_8_49_groupi_g2231(out1[58] ,csa_tree_add_8_49_groupi_n_738 ,csa_tree_add_8_49_groupi_n_434);
  and csa_tree_add_8_49_groupi_g2232(csa_tree_add_8_49_groupi_n_739 ,csa_tree_add_8_49_groupi_n_340 ,csa_tree_add_8_49_groupi_n_738);
  or csa_tree_add_8_49_groupi_g2233(csa_tree_add_8_49_groupi_n_738 ,csa_tree_add_8_49_groupi_n_384 ,csa_tree_add_8_49_groupi_n_736);
  xnor csa_tree_add_8_49_groupi_g2234(out1[57] ,csa_tree_add_8_49_groupi_n_735 ,csa_tree_add_8_49_groupi_n_433);
  and csa_tree_add_8_49_groupi_g2235(csa_tree_add_8_49_groupi_n_736 ,csa_tree_add_8_49_groupi_n_321 ,csa_tree_add_8_49_groupi_n_735);
  or csa_tree_add_8_49_groupi_g2236(csa_tree_add_8_49_groupi_n_735 ,csa_tree_add_8_49_groupi_n_374 ,csa_tree_add_8_49_groupi_n_733);
  xnor csa_tree_add_8_49_groupi_g2237(out1[56] ,csa_tree_add_8_49_groupi_n_732 ,csa_tree_add_8_49_groupi_n_432);
  and csa_tree_add_8_49_groupi_g2238(csa_tree_add_8_49_groupi_n_733 ,csa_tree_add_8_49_groupi_n_364 ,csa_tree_add_8_49_groupi_n_732);
  or csa_tree_add_8_49_groupi_g2239(csa_tree_add_8_49_groupi_n_732 ,csa_tree_add_8_49_groupi_n_368 ,csa_tree_add_8_49_groupi_n_730);
  xnor csa_tree_add_8_49_groupi_g2240(out1[55] ,csa_tree_add_8_49_groupi_n_729 ,csa_tree_add_8_49_groupi_n_431);
  and csa_tree_add_8_49_groupi_g2241(csa_tree_add_8_49_groupi_n_730 ,csa_tree_add_8_49_groupi_n_347 ,csa_tree_add_8_49_groupi_n_729);
  or csa_tree_add_8_49_groupi_g2242(csa_tree_add_8_49_groupi_n_729 ,csa_tree_add_8_49_groupi_n_342 ,csa_tree_add_8_49_groupi_n_727);
  xnor csa_tree_add_8_49_groupi_g2243(out1[54] ,csa_tree_add_8_49_groupi_n_726 ,csa_tree_add_8_49_groupi_n_430);
  and csa_tree_add_8_49_groupi_g2244(csa_tree_add_8_49_groupi_n_727 ,csa_tree_add_8_49_groupi_n_383 ,csa_tree_add_8_49_groupi_n_726);
  or csa_tree_add_8_49_groupi_g2245(csa_tree_add_8_49_groupi_n_726 ,csa_tree_add_8_49_groupi_n_326 ,csa_tree_add_8_49_groupi_n_724);
  xnor csa_tree_add_8_49_groupi_g2246(out1[53] ,csa_tree_add_8_49_groupi_n_723 ,csa_tree_add_8_49_groupi_n_429);
  and csa_tree_add_8_49_groupi_g2247(csa_tree_add_8_49_groupi_n_724 ,csa_tree_add_8_49_groupi_n_320 ,csa_tree_add_8_49_groupi_n_723);
  or csa_tree_add_8_49_groupi_g2248(csa_tree_add_8_49_groupi_n_723 ,csa_tree_add_8_49_groupi_n_329 ,csa_tree_add_8_49_groupi_n_721);
  xnor csa_tree_add_8_49_groupi_g2249(out1[52] ,csa_tree_add_8_49_groupi_n_720 ,csa_tree_add_8_49_groupi_n_428);
  and csa_tree_add_8_49_groupi_g2250(csa_tree_add_8_49_groupi_n_721 ,csa_tree_add_8_49_groupi_n_331 ,csa_tree_add_8_49_groupi_n_720);
  or csa_tree_add_8_49_groupi_g2251(csa_tree_add_8_49_groupi_n_720 ,csa_tree_add_8_49_groupi_n_337 ,csa_tree_add_8_49_groupi_n_718);
  xnor csa_tree_add_8_49_groupi_g2252(out1[51] ,csa_tree_add_8_49_groupi_n_717 ,csa_tree_add_8_49_groupi_n_427);
  and csa_tree_add_8_49_groupi_g2253(csa_tree_add_8_49_groupi_n_718 ,csa_tree_add_8_49_groupi_n_345 ,csa_tree_add_8_49_groupi_n_717);
  or csa_tree_add_8_49_groupi_g2254(csa_tree_add_8_49_groupi_n_717 ,csa_tree_add_8_49_groupi_n_389 ,csa_tree_add_8_49_groupi_n_715);
  xnor csa_tree_add_8_49_groupi_g2255(out1[50] ,csa_tree_add_8_49_groupi_n_714 ,csa_tree_add_8_49_groupi_n_426);
  and csa_tree_add_8_49_groupi_g2256(csa_tree_add_8_49_groupi_n_715 ,csa_tree_add_8_49_groupi_n_344 ,csa_tree_add_8_49_groupi_n_714);
  or csa_tree_add_8_49_groupi_g2257(csa_tree_add_8_49_groupi_n_714 ,csa_tree_add_8_49_groupi_n_373 ,csa_tree_add_8_49_groupi_n_712);
  xnor csa_tree_add_8_49_groupi_g2258(out1[49] ,csa_tree_add_8_49_groupi_n_711 ,csa_tree_add_8_49_groupi_n_441);
  and csa_tree_add_8_49_groupi_g2259(csa_tree_add_8_49_groupi_n_712 ,csa_tree_add_8_49_groupi_n_372 ,csa_tree_add_8_49_groupi_n_711);
  or csa_tree_add_8_49_groupi_g2260(csa_tree_add_8_49_groupi_n_711 ,csa_tree_add_8_49_groupi_n_393 ,csa_tree_add_8_49_groupi_n_709);
  xnor csa_tree_add_8_49_groupi_g2261(out1[48] ,csa_tree_add_8_49_groupi_n_708 ,csa_tree_add_8_49_groupi_n_424);
  and csa_tree_add_8_49_groupi_g2262(csa_tree_add_8_49_groupi_n_709 ,csa_tree_add_8_49_groupi_n_365 ,csa_tree_add_8_49_groupi_n_708);
  or csa_tree_add_8_49_groupi_g2263(csa_tree_add_8_49_groupi_n_708 ,csa_tree_add_8_49_groupi_n_366 ,csa_tree_add_8_49_groupi_n_706);
  xnor csa_tree_add_8_49_groupi_g2264(out1[47] ,csa_tree_add_8_49_groupi_n_705 ,csa_tree_add_8_49_groupi_n_423);
  and csa_tree_add_8_49_groupi_g2265(csa_tree_add_8_49_groupi_n_706 ,csa_tree_add_8_49_groupi_n_371 ,csa_tree_add_8_49_groupi_n_705);
  or csa_tree_add_8_49_groupi_g2266(csa_tree_add_8_49_groupi_n_705 ,csa_tree_add_8_49_groupi_n_376 ,csa_tree_add_8_49_groupi_n_703);
  xnor csa_tree_add_8_49_groupi_g2267(out1[46] ,csa_tree_add_8_49_groupi_n_702 ,csa_tree_add_8_49_groupi_n_422);
  and csa_tree_add_8_49_groupi_g2268(csa_tree_add_8_49_groupi_n_703 ,csa_tree_add_8_49_groupi_n_388 ,csa_tree_add_8_49_groupi_n_702);
  or csa_tree_add_8_49_groupi_g2269(csa_tree_add_8_49_groupi_n_702 ,csa_tree_add_8_49_groupi_n_346 ,csa_tree_add_8_49_groupi_n_700);
  xnor csa_tree_add_8_49_groupi_g2270(out1[45] ,csa_tree_add_8_49_groupi_n_699 ,csa_tree_add_8_49_groupi_n_421);
  and csa_tree_add_8_49_groupi_g2271(csa_tree_add_8_49_groupi_n_700 ,csa_tree_add_8_49_groupi_n_339 ,csa_tree_add_8_49_groupi_n_699);
  or csa_tree_add_8_49_groupi_g2272(csa_tree_add_8_49_groupi_n_699 ,csa_tree_add_8_49_groupi_n_338 ,csa_tree_add_8_49_groupi_n_697);
  xnor csa_tree_add_8_49_groupi_g2273(out1[44] ,csa_tree_add_8_49_groupi_n_696 ,csa_tree_add_8_49_groupi_n_420);
  and csa_tree_add_8_49_groupi_g2274(csa_tree_add_8_49_groupi_n_697 ,csa_tree_add_8_49_groupi_n_334 ,csa_tree_add_8_49_groupi_n_696);
  or csa_tree_add_8_49_groupi_g2275(csa_tree_add_8_49_groupi_n_696 ,csa_tree_add_8_49_groupi_n_332 ,csa_tree_add_8_49_groupi_n_694);
  xnor csa_tree_add_8_49_groupi_g2276(out1[43] ,csa_tree_add_8_49_groupi_n_693 ,csa_tree_add_8_49_groupi_n_418);
  and csa_tree_add_8_49_groupi_g2277(csa_tree_add_8_49_groupi_n_694 ,csa_tree_add_8_49_groupi_n_348 ,csa_tree_add_8_49_groupi_n_693);
  or csa_tree_add_8_49_groupi_g2278(csa_tree_add_8_49_groupi_n_693 ,csa_tree_add_8_49_groupi_n_323 ,csa_tree_add_8_49_groupi_n_691);
  xnor csa_tree_add_8_49_groupi_g2279(out1[42] ,csa_tree_add_8_49_groupi_n_690 ,csa_tree_add_8_49_groupi_n_417);
  and csa_tree_add_8_49_groupi_g2280(csa_tree_add_8_49_groupi_n_691 ,csa_tree_add_8_49_groupi_n_390 ,csa_tree_add_8_49_groupi_n_690);
  or csa_tree_add_8_49_groupi_g2281(csa_tree_add_8_49_groupi_n_690 ,csa_tree_add_8_49_groupi_n_317 ,csa_tree_add_8_49_groupi_n_688);
  xnor csa_tree_add_8_49_groupi_g2282(out1[41] ,csa_tree_add_8_49_groupi_n_687 ,csa_tree_add_8_49_groupi_n_416);
  and csa_tree_add_8_49_groupi_g2283(csa_tree_add_8_49_groupi_n_688 ,csa_tree_add_8_49_groupi_n_325 ,csa_tree_add_8_49_groupi_n_687);
  or csa_tree_add_8_49_groupi_g2284(csa_tree_add_8_49_groupi_n_687 ,csa_tree_add_8_49_groupi_n_327 ,csa_tree_add_8_49_groupi_n_685);
  xnor csa_tree_add_8_49_groupi_g2285(out1[40] ,csa_tree_add_8_49_groupi_n_684 ,csa_tree_add_8_49_groupi_n_415);
  and csa_tree_add_8_49_groupi_g2286(csa_tree_add_8_49_groupi_n_685 ,csa_tree_add_8_49_groupi_n_377 ,csa_tree_add_8_49_groupi_n_684);
  or csa_tree_add_8_49_groupi_g2287(csa_tree_add_8_49_groupi_n_684 ,csa_tree_add_8_49_groupi_n_380 ,csa_tree_add_8_49_groupi_n_682);
  xnor csa_tree_add_8_49_groupi_g2288(out1[39] ,csa_tree_add_8_49_groupi_n_681 ,csa_tree_add_8_49_groupi_n_414);
  and csa_tree_add_8_49_groupi_g2289(csa_tree_add_8_49_groupi_n_682 ,csa_tree_add_8_49_groupi_n_381 ,csa_tree_add_8_49_groupi_n_681);
  or csa_tree_add_8_49_groupi_g2290(csa_tree_add_8_49_groupi_n_681 ,csa_tree_add_8_49_groupi_n_341 ,csa_tree_add_8_49_groupi_n_679);
  xnor csa_tree_add_8_49_groupi_g2291(out1[38] ,csa_tree_add_8_49_groupi_n_678 ,csa_tree_add_8_49_groupi_n_413);
  and csa_tree_add_8_49_groupi_g2292(csa_tree_add_8_49_groupi_n_679 ,csa_tree_add_8_49_groupi_n_385 ,csa_tree_add_8_49_groupi_n_678);
  or csa_tree_add_8_49_groupi_g2293(csa_tree_add_8_49_groupi_n_678 ,csa_tree_add_8_49_groupi_n_391 ,csa_tree_add_8_49_groupi_n_676);
  xnor csa_tree_add_8_49_groupi_g2294(out1[37] ,csa_tree_add_8_49_groupi_n_675 ,csa_tree_add_8_49_groupi_n_412);
  and csa_tree_add_8_49_groupi_g2295(csa_tree_add_8_49_groupi_n_676 ,csa_tree_add_8_49_groupi_n_330 ,csa_tree_add_8_49_groupi_n_675);
  or csa_tree_add_8_49_groupi_g2296(csa_tree_add_8_49_groupi_n_675 ,csa_tree_add_8_49_groupi_n_335 ,csa_tree_add_8_49_groupi_n_673);
  xnor csa_tree_add_8_49_groupi_g2297(out1[36] ,csa_tree_add_8_49_groupi_n_672 ,csa_tree_add_8_49_groupi_n_411);
  and csa_tree_add_8_49_groupi_g2298(csa_tree_add_8_49_groupi_n_673 ,csa_tree_add_8_49_groupi_n_318 ,csa_tree_add_8_49_groupi_n_672);
  or csa_tree_add_8_49_groupi_g2299(csa_tree_add_8_49_groupi_n_672 ,csa_tree_add_8_49_groupi_n_382 ,csa_tree_add_8_49_groupi_n_670);
  xnor csa_tree_add_8_49_groupi_g2300(out1[35] ,csa_tree_add_8_49_groupi_n_669 ,csa_tree_add_8_49_groupi_n_425);
  and csa_tree_add_8_49_groupi_g2301(csa_tree_add_8_49_groupi_n_670 ,csa_tree_add_8_49_groupi_n_343 ,csa_tree_add_8_49_groupi_n_669);
  or csa_tree_add_8_49_groupi_g2302(csa_tree_add_8_49_groupi_n_669 ,csa_tree_add_8_49_groupi_n_375 ,csa_tree_add_8_49_groupi_n_667);
  xnor csa_tree_add_8_49_groupi_g2303(out1[34] ,csa_tree_add_8_49_groupi_n_666 ,csa_tree_add_8_49_groupi_n_440);
  and csa_tree_add_8_49_groupi_g2304(csa_tree_add_8_49_groupi_n_667 ,csa_tree_add_8_49_groupi_n_324 ,csa_tree_add_8_49_groupi_n_666);
  or csa_tree_add_8_49_groupi_g2305(csa_tree_add_8_49_groupi_n_666 ,csa_tree_add_8_49_groupi_n_322 ,csa_tree_add_8_49_groupi_n_664);
  xnor csa_tree_add_8_49_groupi_g2306(out1[33] ,csa_tree_add_8_49_groupi_n_663 ,csa_tree_add_8_49_groupi_n_439);
  and csa_tree_add_8_49_groupi_g2307(csa_tree_add_8_49_groupi_n_664 ,csa_tree_add_8_49_groupi_n_369 ,csa_tree_add_8_49_groupi_n_663);
  or csa_tree_add_8_49_groupi_g2308(csa_tree_add_8_49_groupi_n_663 ,csa_tree_add_8_49_groupi_n_445 ,csa_tree_add_8_49_groupi_n_661);
  xor csa_tree_add_8_49_groupi_g2309(out1[32] ,csa_tree_add_8_49_groupi_n_660 ,csa_tree_add_8_49_groupi_n_478);
  and csa_tree_add_8_49_groupi_g2310(csa_tree_add_8_49_groupi_n_661 ,csa_tree_add_8_49_groupi_n_447 ,csa_tree_add_8_49_groupi_n_660);
  or csa_tree_add_8_49_groupi_g2311(csa_tree_add_8_49_groupi_n_660 ,csa_tree_add_8_49_groupi_n_524 ,csa_tree_add_8_49_groupi_n_658);
  xnor csa_tree_add_8_49_groupi_g2312(out1[31] ,csa_tree_add_8_49_groupi_n_657 ,csa_tree_add_8_49_groupi_n_569);
  and csa_tree_add_8_49_groupi_g2313(csa_tree_add_8_49_groupi_n_658 ,csa_tree_add_8_49_groupi_n_519 ,csa_tree_add_8_49_groupi_n_657);
  or csa_tree_add_8_49_groupi_g2314(csa_tree_add_8_49_groupi_n_657 ,csa_tree_add_8_49_groupi_n_518 ,csa_tree_add_8_49_groupi_n_655);
  xnor csa_tree_add_8_49_groupi_g2315(out1[30] ,csa_tree_add_8_49_groupi_n_654 ,csa_tree_add_8_49_groupi_n_568);
  and csa_tree_add_8_49_groupi_g2316(csa_tree_add_8_49_groupi_n_655 ,csa_tree_add_8_49_groupi_n_513 ,csa_tree_add_8_49_groupi_n_654);
  or csa_tree_add_8_49_groupi_g2317(csa_tree_add_8_49_groupi_n_654 ,csa_tree_add_8_49_groupi_n_512 ,csa_tree_add_8_49_groupi_n_652);
  xnor csa_tree_add_8_49_groupi_g2318(out1[29] ,csa_tree_add_8_49_groupi_n_651 ,csa_tree_add_8_49_groupi_n_567);
  and csa_tree_add_8_49_groupi_g2319(csa_tree_add_8_49_groupi_n_652 ,csa_tree_add_8_49_groupi_n_506 ,csa_tree_add_8_49_groupi_n_651);
  or csa_tree_add_8_49_groupi_g2320(csa_tree_add_8_49_groupi_n_651 ,csa_tree_add_8_49_groupi_n_505 ,csa_tree_add_8_49_groupi_n_649);
  xnor csa_tree_add_8_49_groupi_g2321(out1[28] ,csa_tree_add_8_49_groupi_n_648 ,csa_tree_add_8_49_groupi_n_566);
  and csa_tree_add_8_49_groupi_g2322(csa_tree_add_8_49_groupi_n_649 ,csa_tree_add_8_49_groupi_n_502 ,csa_tree_add_8_49_groupi_n_648);
  or csa_tree_add_8_49_groupi_g2323(csa_tree_add_8_49_groupi_n_648 ,csa_tree_add_8_49_groupi_n_499 ,csa_tree_add_8_49_groupi_n_646);
  xnor csa_tree_add_8_49_groupi_g2324(out1[27] ,csa_tree_add_8_49_groupi_n_645 ,csa_tree_add_8_49_groupi_n_565);
  and csa_tree_add_8_49_groupi_g2325(csa_tree_add_8_49_groupi_n_646 ,csa_tree_add_8_49_groupi_n_494 ,csa_tree_add_8_49_groupi_n_645);
  or csa_tree_add_8_49_groupi_g2326(csa_tree_add_8_49_groupi_n_645 ,csa_tree_add_8_49_groupi_n_493 ,csa_tree_add_8_49_groupi_n_643);
  xnor csa_tree_add_8_49_groupi_g2327(out1[26] ,csa_tree_add_8_49_groupi_n_642 ,csa_tree_add_8_49_groupi_n_564);
  and csa_tree_add_8_49_groupi_g2328(csa_tree_add_8_49_groupi_n_643 ,csa_tree_add_8_49_groupi_n_490 ,csa_tree_add_8_49_groupi_n_642);
  or csa_tree_add_8_49_groupi_g2329(csa_tree_add_8_49_groupi_n_642 ,csa_tree_add_8_49_groupi_n_489 ,csa_tree_add_8_49_groupi_n_640);
  xnor csa_tree_add_8_49_groupi_g2330(out1[25] ,csa_tree_add_8_49_groupi_n_639 ,csa_tree_add_8_49_groupi_n_563);
  and csa_tree_add_8_49_groupi_g2331(csa_tree_add_8_49_groupi_n_640 ,csa_tree_add_8_49_groupi_n_488 ,csa_tree_add_8_49_groupi_n_639);
  or csa_tree_add_8_49_groupi_g2332(csa_tree_add_8_49_groupi_n_639 ,csa_tree_add_8_49_groupi_n_487 ,csa_tree_add_8_49_groupi_n_637);
  xnor csa_tree_add_8_49_groupi_g2333(out1[24] ,csa_tree_add_8_49_groupi_n_636 ,csa_tree_add_8_49_groupi_n_562);
  and csa_tree_add_8_49_groupi_g2334(csa_tree_add_8_49_groupi_n_637 ,csa_tree_add_8_49_groupi_n_486 ,csa_tree_add_8_49_groupi_n_636);
  or csa_tree_add_8_49_groupi_g2335(csa_tree_add_8_49_groupi_n_636 ,csa_tree_add_8_49_groupi_n_485 ,csa_tree_add_8_49_groupi_n_634);
  xnor csa_tree_add_8_49_groupi_g2336(out1[23] ,csa_tree_add_8_49_groupi_n_633 ,csa_tree_add_8_49_groupi_n_561);
  and csa_tree_add_8_49_groupi_g2337(csa_tree_add_8_49_groupi_n_634 ,csa_tree_add_8_49_groupi_n_484 ,csa_tree_add_8_49_groupi_n_633);
  or csa_tree_add_8_49_groupi_g2338(csa_tree_add_8_49_groupi_n_633 ,csa_tree_add_8_49_groupi_n_483 ,csa_tree_add_8_49_groupi_n_631);
  xnor csa_tree_add_8_49_groupi_g2339(out1[22] ,csa_tree_add_8_49_groupi_n_630 ,csa_tree_add_8_49_groupi_n_560);
  and csa_tree_add_8_49_groupi_g2340(csa_tree_add_8_49_groupi_n_631 ,csa_tree_add_8_49_groupi_n_480 ,csa_tree_add_8_49_groupi_n_630);
  or csa_tree_add_8_49_groupi_g2341(csa_tree_add_8_49_groupi_n_630 ,csa_tree_add_8_49_groupi_n_479 ,csa_tree_add_8_49_groupi_n_628);
  xnor csa_tree_add_8_49_groupi_g2342(out1[21] ,csa_tree_add_8_49_groupi_n_627 ,csa_tree_add_8_49_groupi_n_559);
  and csa_tree_add_8_49_groupi_g2343(csa_tree_add_8_49_groupi_n_628 ,csa_tree_add_8_49_groupi_n_539 ,csa_tree_add_8_49_groupi_n_627);
  or csa_tree_add_8_49_groupi_g2344(csa_tree_add_8_49_groupi_n_627 ,csa_tree_add_8_49_groupi_n_538 ,csa_tree_add_8_49_groupi_n_625);
  xnor csa_tree_add_8_49_groupi_g2345(out1[20] ,csa_tree_add_8_49_groupi_n_624 ,csa_tree_add_8_49_groupi_n_558);
  and csa_tree_add_8_49_groupi_g2346(csa_tree_add_8_49_groupi_n_625 ,csa_tree_add_8_49_groupi_n_537 ,csa_tree_add_8_49_groupi_n_624);
  or csa_tree_add_8_49_groupi_g2347(csa_tree_add_8_49_groupi_n_624 ,csa_tree_add_8_49_groupi_n_536 ,csa_tree_add_8_49_groupi_n_622);
  xnor csa_tree_add_8_49_groupi_g2348(out1[19] ,csa_tree_add_8_49_groupi_n_621 ,csa_tree_add_8_49_groupi_n_557);
  and csa_tree_add_8_49_groupi_g2349(csa_tree_add_8_49_groupi_n_622 ,csa_tree_add_8_49_groupi_n_491 ,csa_tree_add_8_49_groupi_n_621);
  or csa_tree_add_8_49_groupi_g2350(csa_tree_add_8_49_groupi_n_621 ,csa_tree_add_8_49_groupi_n_535 ,csa_tree_add_8_49_groupi_n_619);
  xnor csa_tree_add_8_49_groupi_g2351(out1[18] ,csa_tree_add_8_49_groupi_n_618 ,csa_tree_add_8_49_groupi_n_556);
  and csa_tree_add_8_49_groupi_g2352(csa_tree_add_8_49_groupi_n_619 ,csa_tree_add_8_49_groupi_n_482 ,csa_tree_add_8_49_groupi_n_618);
  or csa_tree_add_8_49_groupi_g2353(csa_tree_add_8_49_groupi_n_618 ,csa_tree_add_8_49_groupi_n_481 ,csa_tree_add_8_49_groupi_n_616);
  xnor csa_tree_add_8_49_groupi_g2354(out1[17] ,csa_tree_add_8_49_groupi_n_615 ,csa_tree_add_8_49_groupi_n_541);
  and csa_tree_add_8_49_groupi_g2355(csa_tree_add_8_49_groupi_n_616 ,csa_tree_add_8_49_groupi_n_534 ,csa_tree_add_8_49_groupi_n_615);
  or csa_tree_add_8_49_groupi_g2356(csa_tree_add_8_49_groupi_n_615 ,csa_tree_add_8_49_groupi_n_533 ,csa_tree_add_8_49_groupi_n_613);
  xnor csa_tree_add_8_49_groupi_g2357(out1[16] ,csa_tree_add_8_49_groupi_n_612 ,csa_tree_add_8_49_groupi_n_540);
  and csa_tree_add_8_49_groupi_g2358(csa_tree_add_8_49_groupi_n_613 ,csa_tree_add_8_49_groupi_n_532 ,csa_tree_add_8_49_groupi_n_612);
  or csa_tree_add_8_49_groupi_g2359(csa_tree_add_8_49_groupi_n_612 ,csa_tree_add_8_49_groupi_n_531 ,csa_tree_add_8_49_groupi_n_610);
  xnor csa_tree_add_8_49_groupi_g2360(out1[15] ,csa_tree_add_8_49_groupi_n_609 ,csa_tree_add_8_49_groupi_n_547);
  and csa_tree_add_8_49_groupi_g2361(csa_tree_add_8_49_groupi_n_610 ,csa_tree_add_8_49_groupi_n_530 ,csa_tree_add_8_49_groupi_n_609);
  or csa_tree_add_8_49_groupi_g2362(csa_tree_add_8_49_groupi_n_609 ,csa_tree_add_8_49_groupi_n_529 ,csa_tree_add_8_49_groupi_n_607);
  xnor csa_tree_add_8_49_groupi_g2363(out1[14] ,csa_tree_add_8_49_groupi_n_606 ,csa_tree_add_8_49_groupi_n_553);
  and csa_tree_add_8_49_groupi_g2364(csa_tree_add_8_49_groupi_n_607 ,csa_tree_add_8_49_groupi_n_528 ,csa_tree_add_8_49_groupi_n_606);
  or csa_tree_add_8_49_groupi_g2365(csa_tree_add_8_49_groupi_n_606 ,csa_tree_add_8_49_groupi_n_527 ,csa_tree_add_8_49_groupi_n_604);
  xnor csa_tree_add_8_49_groupi_g2366(out1[13] ,csa_tree_add_8_49_groupi_n_603 ,csa_tree_add_8_49_groupi_n_552);
  and csa_tree_add_8_49_groupi_g2367(csa_tree_add_8_49_groupi_n_604 ,csa_tree_add_8_49_groupi_n_526 ,csa_tree_add_8_49_groupi_n_603);
  or csa_tree_add_8_49_groupi_g2368(csa_tree_add_8_49_groupi_n_603 ,csa_tree_add_8_49_groupi_n_525 ,csa_tree_add_8_49_groupi_n_601);
  xnor csa_tree_add_8_49_groupi_g2369(out1[12] ,csa_tree_add_8_49_groupi_n_600 ,csa_tree_add_8_49_groupi_n_551);
  and csa_tree_add_8_49_groupi_g2370(csa_tree_add_8_49_groupi_n_601 ,csa_tree_add_8_49_groupi_n_523 ,csa_tree_add_8_49_groupi_n_600);
  or csa_tree_add_8_49_groupi_g2371(csa_tree_add_8_49_groupi_n_600 ,csa_tree_add_8_49_groupi_n_522 ,csa_tree_add_8_49_groupi_n_598);
  xnor csa_tree_add_8_49_groupi_g2372(out1[11] ,csa_tree_add_8_49_groupi_n_597 ,csa_tree_add_8_49_groupi_n_550);
  and csa_tree_add_8_49_groupi_g2373(csa_tree_add_8_49_groupi_n_598 ,csa_tree_add_8_49_groupi_n_521 ,csa_tree_add_8_49_groupi_n_597);
  or csa_tree_add_8_49_groupi_g2374(csa_tree_add_8_49_groupi_n_597 ,csa_tree_add_8_49_groupi_n_520 ,csa_tree_add_8_49_groupi_n_595);
  xnor csa_tree_add_8_49_groupi_g2375(out1[10] ,csa_tree_add_8_49_groupi_n_594 ,csa_tree_add_8_49_groupi_n_549);
  and csa_tree_add_8_49_groupi_g2376(csa_tree_add_8_49_groupi_n_595 ,csa_tree_add_8_49_groupi_n_517 ,csa_tree_add_8_49_groupi_n_594);
  or csa_tree_add_8_49_groupi_g2377(csa_tree_add_8_49_groupi_n_594 ,csa_tree_add_8_49_groupi_n_516 ,csa_tree_add_8_49_groupi_n_592);
  xnor csa_tree_add_8_49_groupi_g2378(out1[9] ,csa_tree_add_8_49_groupi_n_591 ,csa_tree_add_8_49_groupi_n_548);
  and csa_tree_add_8_49_groupi_g2379(csa_tree_add_8_49_groupi_n_592 ,csa_tree_add_8_49_groupi_n_515 ,csa_tree_add_8_49_groupi_n_591);
  or csa_tree_add_8_49_groupi_g2380(csa_tree_add_8_49_groupi_n_591 ,csa_tree_add_8_49_groupi_n_514 ,csa_tree_add_8_49_groupi_n_589);
  xnor csa_tree_add_8_49_groupi_g2381(out1[8] ,csa_tree_add_8_49_groupi_n_588 ,csa_tree_add_8_49_groupi_n_554);
  and csa_tree_add_8_49_groupi_g2382(csa_tree_add_8_49_groupi_n_589 ,csa_tree_add_8_49_groupi_n_511 ,csa_tree_add_8_49_groupi_n_588);
  or csa_tree_add_8_49_groupi_g2383(csa_tree_add_8_49_groupi_n_588 ,csa_tree_add_8_49_groupi_n_510 ,csa_tree_add_8_49_groupi_n_586);
  xnor csa_tree_add_8_49_groupi_g2384(out1[7] ,csa_tree_add_8_49_groupi_n_585 ,csa_tree_add_8_49_groupi_n_546);
  and csa_tree_add_8_49_groupi_g2385(csa_tree_add_8_49_groupi_n_586 ,csa_tree_add_8_49_groupi_n_509 ,csa_tree_add_8_49_groupi_n_585);
  or csa_tree_add_8_49_groupi_g2386(csa_tree_add_8_49_groupi_n_585 ,csa_tree_add_8_49_groupi_n_507 ,csa_tree_add_8_49_groupi_n_583);
  xnor csa_tree_add_8_49_groupi_g2387(out1[6] ,csa_tree_add_8_49_groupi_n_582 ,csa_tree_add_8_49_groupi_n_545);
  and csa_tree_add_8_49_groupi_g2388(csa_tree_add_8_49_groupi_n_583 ,csa_tree_add_8_49_groupi_n_504 ,csa_tree_add_8_49_groupi_n_582);
  or csa_tree_add_8_49_groupi_g2389(csa_tree_add_8_49_groupi_n_582 ,csa_tree_add_8_49_groupi_n_503 ,csa_tree_add_8_49_groupi_n_580);
  xnor csa_tree_add_8_49_groupi_g2390(out1[5] ,csa_tree_add_8_49_groupi_n_579 ,csa_tree_add_8_49_groupi_n_544);
  and csa_tree_add_8_49_groupi_g2391(csa_tree_add_8_49_groupi_n_580 ,csa_tree_add_8_49_groupi_n_501 ,csa_tree_add_8_49_groupi_n_579);
  or csa_tree_add_8_49_groupi_g2392(csa_tree_add_8_49_groupi_n_579 ,csa_tree_add_8_49_groupi_n_500 ,csa_tree_add_8_49_groupi_n_577);
  xnor csa_tree_add_8_49_groupi_g2393(out1[4] ,csa_tree_add_8_49_groupi_n_576 ,csa_tree_add_8_49_groupi_n_543);
  and csa_tree_add_8_49_groupi_g2394(csa_tree_add_8_49_groupi_n_577 ,csa_tree_add_8_49_groupi_n_498 ,csa_tree_add_8_49_groupi_n_576);
  or csa_tree_add_8_49_groupi_g2395(csa_tree_add_8_49_groupi_n_576 ,csa_tree_add_8_49_groupi_n_497 ,csa_tree_add_8_49_groupi_n_574);
  xnor csa_tree_add_8_49_groupi_g2396(out1[3] ,csa_tree_add_8_49_groupi_n_572 ,csa_tree_add_8_49_groupi_n_542);
  and csa_tree_add_8_49_groupi_g2397(csa_tree_add_8_49_groupi_n_574 ,csa_tree_add_8_49_groupi_n_496 ,csa_tree_add_8_49_groupi_n_572);
  xor csa_tree_add_8_49_groupi_g2398(out1[2] ,csa_tree_add_8_49_groupi_n_508 ,csa_tree_add_8_49_groupi_n_570);
  or csa_tree_add_8_49_groupi_g2399(csa_tree_add_8_49_groupi_n_572 ,csa_tree_add_8_49_groupi_n_495 ,csa_tree_add_8_49_groupi_n_571);
  and csa_tree_add_8_49_groupi_g2400(csa_tree_add_8_49_groupi_n_571 ,csa_tree_add_8_49_groupi_n_492 ,csa_tree_add_8_49_groupi_n_508);
  xnor csa_tree_add_8_49_groupi_g2401(csa_tree_add_8_49_groupi_n_570 ,csa_tree_add_8_49_groupi_n_173 ,csa_tree_add_8_49_groupi_n_456);
  xnor csa_tree_add_8_49_groupi_g2402(csa_tree_add_8_49_groupi_n_569 ,csa_tree_add_8_49_groupi_n_394 ,csa_tree_add_8_49_groupi_n_469);
  xnor csa_tree_add_8_49_groupi_g2403(csa_tree_add_8_49_groupi_n_568 ,csa_tree_add_8_49_groupi_n_403 ,csa_tree_add_8_49_groupi_n_475);
  xnor csa_tree_add_8_49_groupi_g2404(csa_tree_add_8_49_groupi_n_567 ,csa_tree_add_8_49_groupi_n_396 ,csa_tree_add_8_49_groupi_n_464);
  xnor csa_tree_add_8_49_groupi_g2405(csa_tree_add_8_49_groupi_n_566 ,csa_tree_add_8_49_groupi_n_349 ,csa_tree_add_8_49_groupi_n_461);
  xnor csa_tree_add_8_49_groupi_g2406(csa_tree_add_8_49_groupi_n_565 ,csa_tree_add_8_49_groupi_n_353 ,csa_tree_add_8_49_groupi_n_458);
  xnor csa_tree_add_8_49_groupi_g2407(csa_tree_add_8_49_groupi_n_564 ,csa_tree_add_8_49_groupi_n_357 ,csa_tree_add_8_49_groupi_n_454);
  xnor csa_tree_add_8_49_groupi_g2408(csa_tree_add_8_49_groupi_n_563 ,csa_tree_add_8_49_groupi_n_359 ,csa_tree_add_8_49_groupi_n_453);
  xnor csa_tree_add_8_49_groupi_g2409(csa_tree_add_8_49_groupi_n_562 ,csa_tree_add_8_49_groupi_n_356 ,csa_tree_add_8_49_groupi_n_451);
  xnor csa_tree_add_8_49_groupi_g2410(csa_tree_add_8_49_groupi_n_561 ,csa_tree_add_8_49_groupi_n_360 ,csa_tree_add_8_49_groupi_n_450);
  xnor csa_tree_add_8_49_groupi_g2411(csa_tree_add_8_49_groupi_n_560 ,csa_tree_add_8_49_groupi_n_400 ,csa_tree_add_8_49_groupi_n_449);
  xnor csa_tree_add_8_49_groupi_g2412(csa_tree_add_8_49_groupi_n_559 ,csa_tree_add_8_49_groupi_n_398 ,csa_tree_add_8_49_groupi_n_442);
  xnor csa_tree_add_8_49_groupi_g2413(csa_tree_add_8_49_groupi_n_558 ,csa_tree_add_8_49_groupi_n_397 ,csa_tree_add_8_49_groupi_n_474);
  xnor csa_tree_add_8_49_groupi_g2414(csa_tree_add_8_49_groupi_n_557 ,csa_tree_add_8_49_groupi_n_395 ,csa_tree_add_8_49_groupi_n_466);
  xnor csa_tree_add_8_49_groupi_g2415(csa_tree_add_8_49_groupi_n_556 ,csa_tree_add_8_49_groupi_n_352 ,csa_tree_add_8_49_groupi_n_443);
  xor csa_tree_add_8_49_groupi_g2416(out1[1] ,csa_tree_add_8_49_groupi_n_363 ,csa_tree_add_8_49_groupi_n_444);
  xnor csa_tree_add_8_49_groupi_g2417(csa_tree_add_8_49_groupi_n_554 ,csa_tree_add_8_49_groupi_n_399 ,csa_tree_add_8_49_groupi_n_465);
  xnor csa_tree_add_8_49_groupi_g2418(csa_tree_add_8_49_groupi_n_553 ,csa_tree_add_8_49_groupi_n_402 ,csa_tree_add_8_49_groupi_n_473);
  xnor csa_tree_add_8_49_groupi_g2419(csa_tree_add_8_49_groupi_n_552 ,csa_tree_add_8_49_groupi_n_406 ,csa_tree_add_8_49_groupi_n_472);
  xnor csa_tree_add_8_49_groupi_g2420(csa_tree_add_8_49_groupi_n_551 ,csa_tree_add_8_49_groupi_n_407 ,csa_tree_add_8_49_groupi_n_471);
  xnor csa_tree_add_8_49_groupi_g2421(csa_tree_add_8_49_groupi_n_550 ,csa_tree_add_8_49_groupi_n_409 ,csa_tree_add_8_49_groupi_n_470);
  xnor csa_tree_add_8_49_groupi_g2422(csa_tree_add_8_49_groupi_n_549 ,csa_tree_add_8_49_groupi_n_410 ,csa_tree_add_8_49_groupi_n_468);
  xnor csa_tree_add_8_49_groupi_g2423(csa_tree_add_8_49_groupi_n_548 ,csa_tree_add_8_49_groupi_n_401 ,csa_tree_add_8_49_groupi_n_467);
  xnor csa_tree_add_8_49_groupi_g2424(csa_tree_add_8_49_groupi_n_547 ,csa_tree_add_8_49_groupi_n_361 ,csa_tree_add_8_49_groupi_n_476);
  xnor csa_tree_add_8_49_groupi_g2425(csa_tree_add_8_49_groupi_n_546 ,csa_tree_add_8_49_groupi_n_358 ,csa_tree_add_8_49_groupi_n_463);
  xnor csa_tree_add_8_49_groupi_g2426(csa_tree_add_8_49_groupi_n_545 ,csa_tree_add_8_49_groupi_n_408 ,csa_tree_add_8_49_groupi_n_462);
  xnor csa_tree_add_8_49_groupi_g2427(csa_tree_add_8_49_groupi_n_544 ,csa_tree_add_8_49_groupi_n_350 ,csa_tree_add_8_49_groupi_n_460);
  xnor csa_tree_add_8_49_groupi_g2428(csa_tree_add_8_49_groupi_n_543 ,csa_tree_add_8_49_groupi_n_351 ,csa_tree_add_8_49_groupi_n_459);
  xnor csa_tree_add_8_49_groupi_g2429(csa_tree_add_8_49_groupi_n_542 ,csa_tree_add_8_49_groupi_n_354 ,csa_tree_add_8_49_groupi_n_457);
  xnor csa_tree_add_8_49_groupi_g2430(csa_tree_add_8_49_groupi_n_541 ,csa_tree_add_8_49_groupi_n_355 ,csa_tree_add_8_49_groupi_n_477);
  xnor csa_tree_add_8_49_groupi_g2431(csa_tree_add_8_49_groupi_n_540 ,csa_tree_add_8_49_groupi_n_362 ,csa_tree_add_8_49_groupi_n_452);
  or csa_tree_add_8_49_groupi_g2432(csa_tree_add_8_49_groupi_n_539 ,csa_tree_add_8_49_groupi_n_398 ,csa_tree_add_8_49_groupi_n_442);
  and csa_tree_add_8_49_groupi_g2433(csa_tree_add_8_49_groupi_n_538 ,csa_tree_add_8_49_groupi_n_397 ,csa_tree_add_8_49_groupi_n_474);
  or csa_tree_add_8_49_groupi_g2434(csa_tree_add_8_49_groupi_n_537 ,csa_tree_add_8_49_groupi_n_397 ,csa_tree_add_8_49_groupi_n_474);
  and csa_tree_add_8_49_groupi_g2435(csa_tree_add_8_49_groupi_n_536 ,csa_tree_add_8_49_groupi_n_395 ,csa_tree_add_8_49_groupi_n_466);
  and csa_tree_add_8_49_groupi_g2436(csa_tree_add_8_49_groupi_n_535 ,csa_tree_add_8_49_groupi_n_352 ,csa_tree_add_8_49_groupi_n_443);
  or csa_tree_add_8_49_groupi_g2437(csa_tree_add_8_49_groupi_n_534 ,csa_tree_add_8_49_groupi_n_355 ,csa_tree_add_8_49_groupi_n_477);
  and csa_tree_add_8_49_groupi_g2438(csa_tree_add_8_49_groupi_n_533 ,csa_tree_add_8_49_groupi_n_362 ,csa_tree_add_8_49_groupi_n_452);
  or csa_tree_add_8_49_groupi_g2439(csa_tree_add_8_49_groupi_n_532 ,csa_tree_add_8_49_groupi_n_362 ,csa_tree_add_8_49_groupi_n_452);
  and csa_tree_add_8_49_groupi_g2440(csa_tree_add_8_49_groupi_n_531 ,csa_tree_add_8_49_groupi_n_361 ,csa_tree_add_8_49_groupi_n_476);
  or csa_tree_add_8_49_groupi_g2441(csa_tree_add_8_49_groupi_n_530 ,csa_tree_add_8_49_groupi_n_361 ,csa_tree_add_8_49_groupi_n_476);
  and csa_tree_add_8_49_groupi_g2442(csa_tree_add_8_49_groupi_n_529 ,csa_tree_add_8_49_groupi_n_402 ,csa_tree_add_8_49_groupi_n_473);
  or csa_tree_add_8_49_groupi_g2443(csa_tree_add_8_49_groupi_n_528 ,csa_tree_add_8_49_groupi_n_402 ,csa_tree_add_8_49_groupi_n_473);
  and csa_tree_add_8_49_groupi_g2444(csa_tree_add_8_49_groupi_n_527 ,csa_tree_add_8_49_groupi_n_406 ,csa_tree_add_8_49_groupi_n_472);
  or csa_tree_add_8_49_groupi_g2445(csa_tree_add_8_49_groupi_n_526 ,csa_tree_add_8_49_groupi_n_406 ,csa_tree_add_8_49_groupi_n_472);
  and csa_tree_add_8_49_groupi_g2446(csa_tree_add_8_49_groupi_n_525 ,csa_tree_add_8_49_groupi_n_407 ,csa_tree_add_8_49_groupi_n_471);
  and csa_tree_add_8_49_groupi_g2447(csa_tree_add_8_49_groupi_n_524 ,csa_tree_add_8_49_groupi_n_394 ,csa_tree_add_8_49_groupi_n_469);
  or csa_tree_add_8_49_groupi_g2448(csa_tree_add_8_49_groupi_n_523 ,csa_tree_add_8_49_groupi_n_407 ,csa_tree_add_8_49_groupi_n_471);
  and csa_tree_add_8_49_groupi_g2449(csa_tree_add_8_49_groupi_n_522 ,csa_tree_add_8_49_groupi_n_409 ,csa_tree_add_8_49_groupi_n_470);
  or csa_tree_add_8_49_groupi_g2450(csa_tree_add_8_49_groupi_n_521 ,csa_tree_add_8_49_groupi_n_409 ,csa_tree_add_8_49_groupi_n_470);
  and csa_tree_add_8_49_groupi_g2451(csa_tree_add_8_49_groupi_n_520 ,csa_tree_add_8_49_groupi_n_410 ,csa_tree_add_8_49_groupi_n_468);
  or csa_tree_add_8_49_groupi_g2452(csa_tree_add_8_49_groupi_n_519 ,csa_tree_add_8_49_groupi_n_394 ,csa_tree_add_8_49_groupi_n_469);
  and csa_tree_add_8_49_groupi_g2453(csa_tree_add_8_49_groupi_n_518 ,csa_tree_add_8_49_groupi_n_403 ,csa_tree_add_8_49_groupi_n_475);
  or csa_tree_add_8_49_groupi_g2454(csa_tree_add_8_49_groupi_n_517 ,csa_tree_add_8_49_groupi_n_410 ,csa_tree_add_8_49_groupi_n_468);
  and csa_tree_add_8_49_groupi_g2455(csa_tree_add_8_49_groupi_n_516 ,csa_tree_add_8_49_groupi_n_401 ,csa_tree_add_8_49_groupi_n_467);
  or csa_tree_add_8_49_groupi_g2456(csa_tree_add_8_49_groupi_n_515 ,csa_tree_add_8_49_groupi_n_401 ,csa_tree_add_8_49_groupi_n_467);
  and csa_tree_add_8_49_groupi_g2457(csa_tree_add_8_49_groupi_n_514 ,csa_tree_add_8_49_groupi_n_399 ,csa_tree_add_8_49_groupi_n_465);
  or csa_tree_add_8_49_groupi_g2458(csa_tree_add_8_49_groupi_n_513 ,csa_tree_add_8_49_groupi_n_403 ,csa_tree_add_8_49_groupi_n_475);
  and csa_tree_add_8_49_groupi_g2459(csa_tree_add_8_49_groupi_n_512 ,csa_tree_add_8_49_groupi_n_396 ,csa_tree_add_8_49_groupi_n_464);
  or csa_tree_add_8_49_groupi_g2460(csa_tree_add_8_49_groupi_n_511 ,csa_tree_add_8_49_groupi_n_399 ,csa_tree_add_8_49_groupi_n_465);
  and csa_tree_add_8_49_groupi_g2461(csa_tree_add_8_49_groupi_n_510 ,csa_tree_add_8_49_groupi_n_358 ,csa_tree_add_8_49_groupi_n_463);
  or csa_tree_add_8_49_groupi_g2462(csa_tree_add_8_49_groupi_n_509 ,csa_tree_add_8_49_groupi_n_358 ,csa_tree_add_8_49_groupi_n_463);
  and csa_tree_add_8_49_groupi_g2463(csa_tree_add_8_49_groupi_n_507 ,csa_tree_add_8_49_groupi_n_408 ,csa_tree_add_8_49_groupi_n_462);
  or csa_tree_add_8_49_groupi_g2464(csa_tree_add_8_49_groupi_n_506 ,csa_tree_add_8_49_groupi_n_396 ,csa_tree_add_8_49_groupi_n_464);
  and csa_tree_add_8_49_groupi_g2465(csa_tree_add_8_49_groupi_n_505 ,csa_tree_add_8_49_groupi_n_349 ,csa_tree_add_8_49_groupi_n_461);
  or csa_tree_add_8_49_groupi_g2466(csa_tree_add_8_49_groupi_n_504 ,csa_tree_add_8_49_groupi_n_408 ,csa_tree_add_8_49_groupi_n_462);
  and csa_tree_add_8_49_groupi_g2467(csa_tree_add_8_49_groupi_n_503 ,csa_tree_add_8_49_groupi_n_350 ,csa_tree_add_8_49_groupi_n_460);
  or csa_tree_add_8_49_groupi_g2468(csa_tree_add_8_49_groupi_n_502 ,csa_tree_add_8_49_groupi_n_349 ,csa_tree_add_8_49_groupi_n_461);
  or csa_tree_add_8_49_groupi_g2469(csa_tree_add_8_49_groupi_n_501 ,csa_tree_add_8_49_groupi_n_350 ,csa_tree_add_8_49_groupi_n_460);
  and csa_tree_add_8_49_groupi_g2470(csa_tree_add_8_49_groupi_n_500 ,csa_tree_add_8_49_groupi_n_351 ,csa_tree_add_8_49_groupi_n_459);
  and csa_tree_add_8_49_groupi_g2471(csa_tree_add_8_49_groupi_n_499 ,csa_tree_add_8_49_groupi_n_353 ,csa_tree_add_8_49_groupi_n_458);
  or csa_tree_add_8_49_groupi_g2472(csa_tree_add_8_49_groupi_n_498 ,csa_tree_add_8_49_groupi_n_351 ,csa_tree_add_8_49_groupi_n_459);
  and csa_tree_add_8_49_groupi_g2473(csa_tree_add_8_49_groupi_n_497 ,csa_tree_add_8_49_groupi_n_354 ,csa_tree_add_8_49_groupi_n_457);
  or csa_tree_add_8_49_groupi_g2474(csa_tree_add_8_49_groupi_n_496 ,csa_tree_add_8_49_groupi_n_354 ,csa_tree_add_8_49_groupi_n_457);
  nor csa_tree_add_8_49_groupi_g2475(csa_tree_add_8_49_groupi_n_495 ,csa_tree_add_8_49_groupi_n_173 ,csa_tree_add_8_49_groupi_n_455);
  or csa_tree_add_8_49_groupi_g2476(csa_tree_add_8_49_groupi_n_494 ,csa_tree_add_8_49_groupi_n_353 ,csa_tree_add_8_49_groupi_n_458);
  and csa_tree_add_8_49_groupi_g2477(csa_tree_add_8_49_groupi_n_493 ,csa_tree_add_8_49_groupi_n_357 ,csa_tree_add_8_49_groupi_n_454);
  or csa_tree_add_8_49_groupi_g2478(csa_tree_add_8_49_groupi_n_492 ,csa_tree_add_8_49_groupi_n_172 ,csa_tree_add_8_49_groupi_n_456);
  or csa_tree_add_8_49_groupi_g2479(csa_tree_add_8_49_groupi_n_491 ,csa_tree_add_8_49_groupi_n_395 ,csa_tree_add_8_49_groupi_n_466);
  or csa_tree_add_8_49_groupi_g2480(csa_tree_add_8_49_groupi_n_490 ,csa_tree_add_8_49_groupi_n_357 ,csa_tree_add_8_49_groupi_n_454);
  and csa_tree_add_8_49_groupi_g2481(csa_tree_add_8_49_groupi_n_489 ,csa_tree_add_8_49_groupi_n_359 ,csa_tree_add_8_49_groupi_n_453);
  or csa_tree_add_8_49_groupi_g2482(csa_tree_add_8_49_groupi_n_488 ,csa_tree_add_8_49_groupi_n_359 ,csa_tree_add_8_49_groupi_n_453);
  and csa_tree_add_8_49_groupi_g2483(csa_tree_add_8_49_groupi_n_487 ,csa_tree_add_8_49_groupi_n_356 ,csa_tree_add_8_49_groupi_n_451);
  or csa_tree_add_8_49_groupi_g2484(csa_tree_add_8_49_groupi_n_486 ,csa_tree_add_8_49_groupi_n_356 ,csa_tree_add_8_49_groupi_n_451);
  and csa_tree_add_8_49_groupi_g2485(csa_tree_add_8_49_groupi_n_485 ,csa_tree_add_8_49_groupi_n_360 ,csa_tree_add_8_49_groupi_n_450);
  or csa_tree_add_8_49_groupi_g2486(csa_tree_add_8_49_groupi_n_484 ,csa_tree_add_8_49_groupi_n_360 ,csa_tree_add_8_49_groupi_n_450);
  and csa_tree_add_8_49_groupi_g2487(csa_tree_add_8_49_groupi_n_483 ,csa_tree_add_8_49_groupi_n_400 ,csa_tree_add_8_49_groupi_n_449);
  or csa_tree_add_8_49_groupi_g2488(csa_tree_add_8_49_groupi_n_482 ,csa_tree_add_8_49_groupi_n_352 ,csa_tree_add_8_49_groupi_n_443);
  and csa_tree_add_8_49_groupi_g2489(csa_tree_add_8_49_groupi_n_481 ,csa_tree_add_8_49_groupi_n_355 ,csa_tree_add_8_49_groupi_n_477);
  or csa_tree_add_8_49_groupi_g2490(csa_tree_add_8_49_groupi_n_480 ,csa_tree_add_8_49_groupi_n_400 ,csa_tree_add_8_49_groupi_n_449);
  and csa_tree_add_8_49_groupi_g2491(csa_tree_add_8_49_groupi_n_479 ,csa_tree_add_8_49_groupi_n_398 ,csa_tree_add_8_49_groupi_n_442);
  xnor csa_tree_add_8_49_groupi_g2492(csa_tree_add_8_49_groupi_n_478 ,csa_tree_add_8_49_groupi_n_245 ,csa_tree_add_8_49_groupi_n_405);
  or csa_tree_add_8_49_groupi_g2493(csa_tree_add_8_49_groupi_n_508 ,csa_tree_add_8_49_groupi_n_370 ,csa_tree_add_8_49_groupi_n_446);
  not csa_tree_add_8_49_groupi_g2494(csa_tree_add_8_49_groupi_n_455 ,csa_tree_add_8_49_groupi_n_456);
  xnor csa_tree_add_8_49_groupi_g2495(out1[0] ,csa_tree_add_8_49_groupi_n_213 ,in3[0]);
  or csa_tree_add_8_49_groupi_g2496(csa_tree_add_8_49_groupi_n_447 ,csa_tree_add_8_49_groupi_n_244 ,csa_tree_add_8_49_groupi_n_405);
  and csa_tree_add_8_49_groupi_g2497(csa_tree_add_8_49_groupi_n_446 ,csa_tree_add_8_49_groupi_n_363 ,csa_tree_add_8_49_groupi_n_392);
  nor csa_tree_add_8_49_groupi_g2498(csa_tree_add_8_49_groupi_n_445 ,csa_tree_add_8_49_groupi_n_245 ,csa_tree_add_8_49_groupi_n_404);
  xnor csa_tree_add_8_49_groupi_g2499(csa_tree_add_8_49_groupi_n_444 ,csa_tree_add_8_49_groupi_n_235 ,n_1878);
  xnor csa_tree_add_8_49_groupi_g2500(csa_tree_add_8_49_groupi_n_477 ,csa_tree_add_8_49_groupi_n_265 ,n_1830);
  xnor csa_tree_add_8_49_groupi_g2501(csa_tree_add_8_49_groupi_n_476 ,csa_tree_add_8_49_groupi_n_264 ,n_1828);
  xnor csa_tree_add_8_49_groupi_g2502(csa_tree_add_8_49_groupi_n_475 ,csa_tree_add_8_49_groupi_n_204 ,n_1843);
  xnor csa_tree_add_8_49_groupi_g2503(csa_tree_add_8_49_groupi_n_474 ,csa_tree_add_8_49_groupi_n_195 ,n_1833);
  xnor csa_tree_add_8_49_groupi_g2504(csa_tree_add_8_49_groupi_n_473 ,csa_tree_add_8_49_groupi_n_212 ,n_1827);
  xnor csa_tree_add_8_49_groupi_g2505(csa_tree_add_8_49_groupi_n_472 ,csa_tree_add_8_49_groupi_n_209 ,n_1826);
  xnor csa_tree_add_8_49_groupi_g2506(csa_tree_add_8_49_groupi_n_471 ,csa_tree_add_8_49_groupi_n_207 ,n_1825);
  xnor csa_tree_add_8_49_groupi_g2507(csa_tree_add_8_49_groupi_n_470 ,csa_tree_add_8_49_groupi_n_269 ,n_1824);
  xnor csa_tree_add_8_49_groupi_g2508(csa_tree_add_8_49_groupi_n_469 ,csa_tree_add_8_49_groupi_n_206 ,n_1844);
  xnor csa_tree_add_8_49_groupi_g2509(csa_tree_add_8_49_groupi_n_468 ,csa_tree_add_8_49_groupi_n_205 ,n_1823);
  xnor csa_tree_add_8_49_groupi_g2510(csa_tree_add_8_49_groupi_n_467 ,csa_tree_add_8_49_groupi_n_203 ,n_1822);
  xnor csa_tree_add_8_49_groupi_g2511(csa_tree_add_8_49_groupi_n_466 ,csa_tree_add_8_49_groupi_n_210 ,n_1832);
  xnor csa_tree_add_8_49_groupi_g2512(csa_tree_add_8_49_groupi_n_465 ,csa_tree_add_8_49_groupi_n_202 ,n_1821);
  xnor csa_tree_add_8_49_groupi_g2513(csa_tree_add_8_49_groupi_n_464 ,csa_tree_add_8_49_groupi_n_201 ,n_1842);
  xnor csa_tree_add_8_49_groupi_g2514(csa_tree_add_8_49_groupi_n_463 ,csa_tree_add_8_49_groupi_n_200 ,n_1820);
  xnor csa_tree_add_8_49_groupi_g2515(csa_tree_add_8_49_groupi_n_462 ,csa_tree_add_8_49_groupi_n_199 ,n_1819);
  xnor csa_tree_add_8_49_groupi_g2516(csa_tree_add_8_49_groupi_n_461 ,csa_tree_add_8_49_groupi_n_191 ,n_1841);
  xnor csa_tree_add_8_49_groupi_g2517(csa_tree_add_8_49_groupi_n_460 ,csa_tree_add_8_49_groupi_n_190 ,n_1818);
  xnor csa_tree_add_8_49_groupi_g2518(csa_tree_add_8_49_groupi_n_459 ,csa_tree_add_8_49_groupi_n_196 ,n_1817);
  xnor csa_tree_add_8_49_groupi_g2519(csa_tree_add_8_49_groupi_n_458 ,csa_tree_add_8_49_groupi_n_197 ,n_1840);
  xnor csa_tree_add_8_49_groupi_g2520(csa_tree_add_8_49_groupi_n_457 ,csa_tree_add_8_49_groupi_n_193 ,n_1816);
  xnor csa_tree_add_8_49_groupi_g2521(csa_tree_add_8_49_groupi_n_456 ,csa_tree_add_8_49_groupi_n_194 ,n_1815);
  xnor csa_tree_add_8_49_groupi_g2522(csa_tree_add_8_49_groupi_n_454 ,csa_tree_add_8_49_groupi_n_263 ,n_1839);
  xnor csa_tree_add_8_49_groupi_g2523(csa_tree_add_8_49_groupi_n_453 ,csa_tree_add_8_49_groupi_n_192 ,n_1838);
  xnor csa_tree_add_8_49_groupi_g2524(csa_tree_add_8_49_groupi_n_452 ,csa_tree_add_8_49_groupi_n_208 ,n_1829);
  xnor csa_tree_add_8_49_groupi_g2525(csa_tree_add_8_49_groupi_n_451 ,csa_tree_add_8_49_groupi_n_267 ,n_1837);
  xnor csa_tree_add_8_49_groupi_g2526(csa_tree_add_8_49_groupi_n_450 ,csa_tree_add_8_49_groupi_n_262 ,n_1836);
  xnor csa_tree_add_8_49_groupi_g2527(csa_tree_add_8_49_groupi_n_449 ,csa_tree_add_8_49_groupi_n_211 ,n_1835);
  xnor csa_tree_add_8_49_groupi_g2528(csa_tree_add_8_49_groupi_n_441 ,csa_tree_add_8_49_groupi_n_112 ,csa_tree_add_8_49_groupi_n_314);
  xnor csa_tree_add_8_49_groupi_g2529(csa_tree_add_8_49_groupi_n_440 ,csa_tree_add_8_49_groupi_n_102 ,csa_tree_add_8_49_groupi_n_241);
  xnor csa_tree_add_8_49_groupi_g2530(csa_tree_add_8_49_groupi_n_439 ,csa_tree_add_8_49_groupi_n_161 ,csa_tree_add_8_49_groupi_n_261);
  xnor csa_tree_add_8_49_groupi_g2531(csa_tree_add_8_49_groupi_n_438 ,csa_tree_add_8_49_groupi_n_159 ,csa_tree_add_8_49_groupi_n_221);
  xnor csa_tree_add_8_49_groupi_g2532(csa_tree_add_8_49_groupi_n_437 ,csa_tree_add_8_49_groupi_n_185 ,csa_tree_add_8_49_groupi_n_223);
  xnor csa_tree_add_8_49_groupi_g2533(csa_tree_add_8_49_groupi_n_436 ,csa_tree_add_8_49_groupi_n_181 ,csa_tree_add_8_49_groupi_n_233);
  xnor csa_tree_add_8_49_groupi_g2534(csa_tree_add_8_49_groupi_n_435 ,csa_tree_add_8_49_groupi_n_118 ,csa_tree_add_8_49_groupi_n_253);
  xnor csa_tree_add_8_49_groupi_g2535(csa_tree_add_8_49_groupi_n_434 ,csa_tree_add_8_49_groupi_n_163 ,csa_tree_add_8_49_groupi_n_257);
  xnor csa_tree_add_8_49_groupi_g2536(csa_tree_add_8_49_groupi_n_433 ,csa_tree_add_8_49_groupi_n_124 ,csa_tree_add_8_49_groupi_n_306);
  xnor csa_tree_add_8_49_groupi_g2537(csa_tree_add_8_49_groupi_n_432 ,csa_tree_add_8_49_groupi_n_179 ,csa_tree_add_8_49_groupi_n_259);
  xnor csa_tree_add_8_49_groupi_g2538(csa_tree_add_8_49_groupi_n_431 ,csa_tree_add_8_49_groupi_n_165 ,csa_tree_add_8_49_groupi_n_231);
  xnor csa_tree_add_8_49_groupi_g2539(csa_tree_add_8_49_groupi_n_430 ,csa_tree_add_8_49_groupi_n_106 ,csa_tree_add_8_49_groupi_n_249);
  xnor csa_tree_add_8_49_groupi_g2540(csa_tree_add_8_49_groupi_n_429 ,csa_tree_add_8_49_groupi_n_110 ,csa_tree_add_8_49_groupi_n_229);
  xnor csa_tree_add_8_49_groupi_g2541(csa_tree_add_8_49_groupi_n_428 ,csa_tree_add_8_49_groupi_n_116 ,csa_tree_add_8_49_groupi_n_225);
  xnor csa_tree_add_8_49_groupi_g2542(csa_tree_add_8_49_groupi_n_427 ,csa_tree_add_8_49_groupi_n_189 ,csa_tree_add_8_49_groupi_n_304);
  xnor csa_tree_add_8_49_groupi_g2543(csa_tree_add_8_49_groupi_n_426 ,csa_tree_add_8_49_groupi_n_171 ,csa_tree_add_8_49_groupi_n_310);
  xnor csa_tree_add_8_49_groupi_g2544(csa_tree_add_8_49_groupi_n_425 ,csa_tree_add_8_49_groupi_n_175 ,csa_tree_add_8_49_groupi_n_255);
  xnor csa_tree_add_8_49_groupi_g2545(csa_tree_add_8_49_groupi_n_424 ,csa_tree_add_8_49_groupi_n_169 ,csa_tree_add_8_49_groupi_n_219);
  xnor csa_tree_add_8_49_groupi_g2546(csa_tree_add_8_49_groupi_n_423 ,csa_tree_add_8_49_groupi_n_177 ,csa_tree_add_8_49_groupi_n_251);
  xnor csa_tree_add_8_49_groupi_g2547(csa_tree_add_8_49_groupi_n_422 ,csa_tree_add_8_49_groupi_n_108 ,csa_tree_add_8_49_groupi_n_217);
  xnor csa_tree_add_8_49_groupi_g2548(csa_tree_add_8_49_groupi_n_421 ,csa_tree_add_8_49_groupi_n_183 ,csa_tree_add_8_49_groupi_n_243);
  xnor csa_tree_add_8_49_groupi_g2549(csa_tree_add_8_49_groupi_n_420 ,csa_tree_add_8_49_groupi_n_126 ,csa_tree_add_8_49_groupi_n_247);
  xnor csa_tree_add_8_49_groupi_g2550(csa_tree_add_8_49_groupi_n_419 ,csa_tree_add_8_49_groupi_n_127 ,csa_tree_add_8_49_groupi_n_268);
  xnor csa_tree_add_8_49_groupi_g2551(csa_tree_add_8_49_groupi_n_418 ,csa_tree_add_8_49_groupi_n_114 ,csa_tree_add_8_49_groupi_n_237);
  xnor csa_tree_add_8_49_groupi_g2552(csa_tree_add_8_49_groupi_n_417 ,csa_tree_add_8_49_groupi_n_98 ,csa_tree_add_8_49_groupi_n_227);
  xnor csa_tree_add_8_49_groupi_g2553(csa_tree_add_8_49_groupi_n_416 ,csa_tree_add_8_49_groupi_n_122 ,csa_tree_add_8_49_groupi_n_308);
  xnor csa_tree_add_8_49_groupi_g2554(csa_tree_add_8_49_groupi_n_415 ,csa_tree_add_8_49_groupi_n_104 ,csa_tree_add_8_49_groupi_n_239);
  xnor csa_tree_add_8_49_groupi_g2555(csa_tree_add_8_49_groupi_n_414 ,csa_tree_add_8_49_groupi_n_187 ,csa_tree_add_8_49_groupi_n_215);
  xnor csa_tree_add_8_49_groupi_g2556(csa_tree_add_8_49_groupi_n_413 ,csa_tree_add_8_49_groupi_n_167 ,csa_tree_add_8_49_groupi_n_316);
  xnor csa_tree_add_8_49_groupi_g2557(csa_tree_add_8_49_groupi_n_412 ,csa_tree_add_8_49_groupi_n_120 ,csa_tree_add_8_49_groupi_n_302);
  xnor csa_tree_add_8_49_groupi_g2558(csa_tree_add_8_49_groupi_n_411 ,csa_tree_add_8_49_groupi_n_100 ,csa_tree_add_8_49_groupi_n_312);
  xnor csa_tree_add_8_49_groupi_g2559(csa_tree_add_8_49_groupi_n_443 ,csa_tree_add_8_49_groupi_n_198 ,n_1831);
  xnor csa_tree_add_8_49_groupi_g2560(csa_tree_add_8_49_groupi_n_442 ,csa_tree_add_8_49_groupi_n_266 ,n_1834);
  not csa_tree_add_8_49_groupi_g2561(csa_tree_add_8_49_groupi_n_404 ,csa_tree_add_8_49_groupi_n_405);
  nor csa_tree_add_8_49_groupi_g2562(csa_tree_add_8_49_groupi_n_393 ,csa_tree_add_8_49_groupi_n_169 ,csa_tree_add_8_49_groupi_n_219);
  or csa_tree_add_8_49_groupi_g2563(csa_tree_add_8_49_groupi_n_392 ,n_1878 ,csa_tree_add_8_49_groupi_n_234);
  nor csa_tree_add_8_49_groupi_g2564(csa_tree_add_8_49_groupi_n_391 ,csa_tree_add_8_49_groupi_n_120 ,csa_tree_add_8_49_groupi_n_302);
  or csa_tree_add_8_49_groupi_g2565(csa_tree_add_8_49_groupi_n_390 ,csa_tree_add_8_49_groupi_n_97 ,csa_tree_add_8_49_groupi_n_226);
  nor csa_tree_add_8_49_groupi_g2566(csa_tree_add_8_49_groupi_n_389 ,csa_tree_add_8_49_groupi_n_171 ,csa_tree_add_8_49_groupi_n_310);
  or csa_tree_add_8_49_groupi_g2567(csa_tree_add_8_49_groupi_n_388 ,csa_tree_add_8_49_groupi_n_107 ,csa_tree_add_8_49_groupi_n_216);
  or csa_tree_add_8_49_groupi_g2568(csa_tree_add_8_49_groupi_n_387 ,csa_tree_add_8_49_groupi_n_184 ,csa_tree_add_8_49_groupi_n_222);
  nor csa_tree_add_8_49_groupi_g2569(csa_tree_add_8_49_groupi_n_386 ,csa_tree_add_8_49_groupi_n_118 ,csa_tree_add_8_49_groupi_n_253);
  or csa_tree_add_8_49_groupi_g2570(csa_tree_add_8_49_groupi_n_385 ,csa_tree_add_8_49_groupi_n_166 ,csa_tree_add_8_49_groupi_n_315);
  nor csa_tree_add_8_49_groupi_g2571(csa_tree_add_8_49_groupi_n_384 ,csa_tree_add_8_49_groupi_n_124 ,csa_tree_add_8_49_groupi_n_306);
  or csa_tree_add_8_49_groupi_g2572(csa_tree_add_8_49_groupi_n_383 ,csa_tree_add_8_49_groupi_n_105 ,csa_tree_add_8_49_groupi_n_248);
  nor csa_tree_add_8_49_groupi_g2573(csa_tree_add_8_49_groupi_n_382 ,csa_tree_add_8_49_groupi_n_175 ,csa_tree_add_8_49_groupi_n_255);
  or csa_tree_add_8_49_groupi_g2574(csa_tree_add_8_49_groupi_n_381 ,csa_tree_add_8_49_groupi_n_186 ,csa_tree_add_8_49_groupi_n_214);
  nor csa_tree_add_8_49_groupi_g2575(csa_tree_add_8_49_groupi_n_380 ,csa_tree_add_8_49_groupi_n_187 ,csa_tree_add_8_49_groupi_n_215);
  or csa_tree_add_8_49_groupi_g2576(csa_tree_add_8_49_groupi_n_379 ,csa_tree_add_8_49_groupi_n_158 ,csa_tree_add_8_49_groupi_n_220);
  nor csa_tree_add_8_49_groupi_g2577(csa_tree_add_8_49_groupi_n_378 ,csa_tree_add_8_49_groupi_n_181 ,csa_tree_add_8_49_groupi_n_233);
  or csa_tree_add_8_49_groupi_g2578(csa_tree_add_8_49_groupi_n_377 ,csa_tree_add_8_49_groupi_n_103 ,csa_tree_add_8_49_groupi_n_238);
  nor csa_tree_add_8_49_groupi_g2579(csa_tree_add_8_49_groupi_n_376 ,csa_tree_add_8_49_groupi_n_108 ,csa_tree_add_8_49_groupi_n_217);
  nor csa_tree_add_8_49_groupi_g2580(csa_tree_add_8_49_groupi_n_375 ,csa_tree_add_8_49_groupi_n_102 ,csa_tree_add_8_49_groupi_n_241);
  nor csa_tree_add_8_49_groupi_g2581(csa_tree_add_8_49_groupi_n_374 ,csa_tree_add_8_49_groupi_n_179 ,csa_tree_add_8_49_groupi_n_259);
  nor csa_tree_add_8_49_groupi_g2582(csa_tree_add_8_49_groupi_n_373 ,csa_tree_add_8_49_groupi_n_112 ,csa_tree_add_8_49_groupi_n_314);
  or csa_tree_add_8_49_groupi_g2583(csa_tree_add_8_49_groupi_n_372 ,csa_tree_add_8_49_groupi_n_111 ,csa_tree_add_8_49_groupi_n_313);
  or csa_tree_add_8_49_groupi_g2584(csa_tree_add_8_49_groupi_n_371 ,csa_tree_add_8_49_groupi_n_176 ,csa_tree_add_8_49_groupi_n_250);
  nor csa_tree_add_8_49_groupi_g2585(csa_tree_add_8_49_groupi_n_370 ,csa_tree_add_8_49_groupi_n_0 ,csa_tree_add_8_49_groupi_n_235);
  or csa_tree_add_8_49_groupi_g2586(csa_tree_add_8_49_groupi_n_369 ,csa_tree_add_8_49_groupi_n_160 ,csa_tree_add_8_49_groupi_n_260);
  nor csa_tree_add_8_49_groupi_g2587(csa_tree_add_8_49_groupi_n_368 ,csa_tree_add_8_49_groupi_n_165 ,csa_tree_add_8_49_groupi_n_231);
  or csa_tree_add_8_49_groupi_g2588(csa_tree_add_8_49_groupi_n_367 ,csa_tree_add_8_49_groupi_n_180 ,csa_tree_add_8_49_groupi_n_232);
  nor csa_tree_add_8_49_groupi_g2589(csa_tree_add_8_49_groupi_n_366 ,csa_tree_add_8_49_groupi_n_177 ,csa_tree_add_8_49_groupi_n_251);
  or csa_tree_add_8_49_groupi_g2590(csa_tree_add_8_49_groupi_n_365 ,csa_tree_add_8_49_groupi_n_168 ,csa_tree_add_8_49_groupi_n_218);
  or csa_tree_add_8_49_groupi_g2591(csa_tree_add_8_49_groupi_n_364 ,csa_tree_add_8_49_groupi_n_178 ,csa_tree_add_8_49_groupi_n_258);
  or csa_tree_add_8_49_groupi_g2592(csa_tree_add_8_49_groupi_n_410 ,csa_tree_add_8_49_groupi_n_152 ,csa_tree_add_8_49_groupi_n_288);
  or csa_tree_add_8_49_groupi_g2593(csa_tree_add_8_49_groupi_n_409 ,csa_tree_add_8_49_groupi_n_87 ,csa_tree_add_8_49_groupi_n_290);
  or csa_tree_add_8_49_groupi_g2594(csa_tree_add_8_49_groupi_n_408 ,csa_tree_add_8_49_groupi_n_84 ,csa_tree_add_8_49_groupi_n_282);
  or csa_tree_add_8_49_groupi_g2595(csa_tree_add_8_49_groupi_n_407 ,csa_tree_add_8_49_groupi_n_135 ,csa_tree_add_8_49_groupi_n_292);
  or csa_tree_add_8_49_groupi_g2596(csa_tree_add_8_49_groupi_n_406 ,csa_tree_add_8_49_groupi_n_146 ,csa_tree_add_8_49_groupi_n_293);
  or csa_tree_add_8_49_groupi_g2597(csa_tree_add_8_49_groupi_n_405 ,csa_tree_add_8_49_groupi_n_131 ,csa_tree_add_8_49_groupi_n_294);
  or csa_tree_add_8_49_groupi_g2598(csa_tree_add_8_49_groupi_n_403 ,csa_tree_add_8_49_groupi_n_78 ,csa_tree_add_8_49_groupi_n_287);
  or csa_tree_add_8_49_groupi_g2599(csa_tree_add_8_49_groupi_n_402 ,csa_tree_add_8_49_groupi_n_154 ,csa_tree_add_8_49_groupi_n_295);
  or csa_tree_add_8_49_groupi_g2600(csa_tree_add_8_49_groupi_n_401 ,csa_tree_add_8_49_groupi_n_93 ,csa_tree_add_8_49_groupi_n_286);
  or csa_tree_add_8_49_groupi_g2601(csa_tree_add_8_49_groupi_n_400 ,csa_tree_add_8_49_groupi_n_156 ,csa_tree_add_8_49_groupi_n_289);
  or csa_tree_add_8_49_groupi_g2602(csa_tree_add_8_49_groupi_n_399 ,csa_tree_add_8_49_groupi_n_70 ,csa_tree_add_8_49_groupi_n_285);
  or csa_tree_add_8_49_groupi_g2603(csa_tree_add_8_49_groupi_n_398 ,csa_tree_add_8_49_groupi_n_66 ,csa_tree_add_8_49_groupi_n_297);
  or csa_tree_add_8_49_groupi_g2604(csa_tree_add_8_49_groupi_n_397 ,csa_tree_add_8_49_groupi_n_82 ,csa_tree_add_8_49_groupi_n_277);
  or csa_tree_add_8_49_groupi_g2605(csa_tree_add_8_49_groupi_n_396 ,csa_tree_add_8_49_groupi_n_65 ,csa_tree_add_8_49_groupi_n_284);
  or csa_tree_add_8_49_groupi_g2606(csa_tree_add_8_49_groupi_n_395 ,csa_tree_add_8_49_groupi_n_81 ,csa_tree_add_8_49_groupi_n_299);
  or csa_tree_add_8_49_groupi_g2607(csa_tree_add_8_49_groupi_n_394 ,csa_tree_add_8_49_groupi_n_157 ,csa_tree_add_8_49_groupi_n_291);
  or csa_tree_add_8_49_groupi_g2608(csa_tree_add_8_49_groupi_n_348 ,csa_tree_add_8_49_groupi_n_113 ,csa_tree_add_8_49_groupi_n_236);
  or csa_tree_add_8_49_groupi_g2609(csa_tree_add_8_49_groupi_n_347 ,csa_tree_add_8_49_groupi_n_164 ,csa_tree_add_8_49_groupi_n_230);
  nor csa_tree_add_8_49_groupi_g2610(csa_tree_add_8_49_groupi_n_346 ,csa_tree_add_8_49_groupi_n_183 ,csa_tree_add_8_49_groupi_n_243);
  or csa_tree_add_8_49_groupi_g2611(csa_tree_add_8_49_groupi_n_345 ,csa_tree_add_8_49_groupi_n_188 ,csa_tree_add_8_49_groupi_n_303);
  or csa_tree_add_8_49_groupi_g2612(csa_tree_add_8_49_groupi_n_344 ,csa_tree_add_8_49_groupi_n_170 ,csa_tree_add_8_49_groupi_n_309);
  or csa_tree_add_8_49_groupi_g2613(csa_tree_add_8_49_groupi_n_343 ,csa_tree_add_8_49_groupi_n_174 ,csa_tree_add_8_49_groupi_n_254);
  nor csa_tree_add_8_49_groupi_g2614(csa_tree_add_8_49_groupi_n_342 ,csa_tree_add_8_49_groupi_n_106 ,csa_tree_add_8_49_groupi_n_249);
  nor csa_tree_add_8_49_groupi_g2615(csa_tree_add_8_49_groupi_n_341 ,csa_tree_add_8_49_groupi_n_167 ,csa_tree_add_8_49_groupi_n_316);
  or csa_tree_add_8_49_groupi_g2616(csa_tree_add_8_49_groupi_n_340 ,csa_tree_add_8_49_groupi_n_162 ,csa_tree_add_8_49_groupi_n_256);
  or csa_tree_add_8_49_groupi_g2617(csa_tree_add_8_49_groupi_n_339 ,csa_tree_add_8_49_groupi_n_182 ,csa_tree_add_8_49_groupi_n_242);
  nor csa_tree_add_8_49_groupi_g2618(csa_tree_add_8_49_groupi_n_338 ,csa_tree_add_8_49_groupi_n_126 ,csa_tree_add_8_49_groupi_n_247);
  nor csa_tree_add_8_49_groupi_g2619(csa_tree_add_8_49_groupi_n_337 ,csa_tree_add_8_49_groupi_n_189 ,csa_tree_add_8_49_groupi_n_304);
  nor csa_tree_add_8_49_groupi_g2620(csa_tree_add_8_49_groupi_n_336 ,csa_tree_add_8_49_groupi_n_159 ,csa_tree_add_8_49_groupi_n_221);
  nor csa_tree_add_8_49_groupi_g2621(csa_tree_add_8_49_groupi_n_335 ,csa_tree_add_8_49_groupi_n_100 ,csa_tree_add_8_49_groupi_n_312);
  or csa_tree_add_8_49_groupi_g2622(csa_tree_add_8_49_groupi_n_334 ,csa_tree_add_8_49_groupi_n_125 ,csa_tree_add_8_49_groupi_n_246);
  nor csa_tree_add_8_49_groupi_g2623(csa_tree_add_8_49_groupi_n_333 ,csa_tree_add_8_49_groupi_n_185 ,csa_tree_add_8_49_groupi_n_223);
  nor csa_tree_add_8_49_groupi_g2624(csa_tree_add_8_49_groupi_n_332 ,csa_tree_add_8_49_groupi_n_114 ,csa_tree_add_8_49_groupi_n_237);
  or csa_tree_add_8_49_groupi_g2625(csa_tree_add_8_49_groupi_n_331 ,csa_tree_add_8_49_groupi_n_115 ,csa_tree_add_8_49_groupi_n_224);
  or csa_tree_add_8_49_groupi_g2626(csa_tree_add_8_49_groupi_n_330 ,csa_tree_add_8_49_groupi_n_119 ,csa_tree_add_8_49_groupi_n_301);
  nor csa_tree_add_8_49_groupi_g2627(csa_tree_add_8_49_groupi_n_329 ,csa_tree_add_8_49_groupi_n_116 ,csa_tree_add_8_49_groupi_n_225);
  or csa_tree_add_8_49_groupi_g2628(csa_tree_add_8_49_groupi_n_328 ,csa_tree_add_8_49_groupi_n_117 ,csa_tree_add_8_49_groupi_n_252);
  nor csa_tree_add_8_49_groupi_g2629(csa_tree_add_8_49_groupi_n_327 ,csa_tree_add_8_49_groupi_n_104 ,csa_tree_add_8_49_groupi_n_239);
  nor csa_tree_add_8_49_groupi_g2630(csa_tree_add_8_49_groupi_n_326 ,csa_tree_add_8_49_groupi_n_110 ,csa_tree_add_8_49_groupi_n_229);
  or csa_tree_add_8_49_groupi_g2631(csa_tree_add_8_49_groupi_n_325 ,csa_tree_add_8_49_groupi_n_121 ,csa_tree_add_8_49_groupi_n_307);
  or csa_tree_add_8_49_groupi_g2632(csa_tree_add_8_49_groupi_n_324 ,csa_tree_add_8_49_groupi_n_101 ,csa_tree_add_8_49_groupi_n_240);
  nor csa_tree_add_8_49_groupi_g2633(csa_tree_add_8_49_groupi_n_323 ,csa_tree_add_8_49_groupi_n_98 ,csa_tree_add_8_49_groupi_n_227);
  nor csa_tree_add_8_49_groupi_g2634(csa_tree_add_8_49_groupi_n_322 ,csa_tree_add_8_49_groupi_n_161 ,csa_tree_add_8_49_groupi_n_261);
  or csa_tree_add_8_49_groupi_g2635(csa_tree_add_8_49_groupi_n_321 ,csa_tree_add_8_49_groupi_n_123 ,csa_tree_add_8_49_groupi_n_305);
  or csa_tree_add_8_49_groupi_g2636(csa_tree_add_8_49_groupi_n_320 ,csa_tree_add_8_49_groupi_n_109 ,csa_tree_add_8_49_groupi_n_228);
  nor csa_tree_add_8_49_groupi_g2637(csa_tree_add_8_49_groupi_n_319 ,csa_tree_add_8_49_groupi_n_163 ,csa_tree_add_8_49_groupi_n_257);
  or csa_tree_add_8_49_groupi_g2638(csa_tree_add_8_49_groupi_n_318 ,csa_tree_add_8_49_groupi_n_99 ,csa_tree_add_8_49_groupi_n_311);
  nor csa_tree_add_8_49_groupi_g2639(csa_tree_add_8_49_groupi_n_317 ,csa_tree_add_8_49_groupi_n_122 ,csa_tree_add_8_49_groupi_n_308);
  or csa_tree_add_8_49_groupi_g2640(csa_tree_add_8_49_groupi_n_363 ,csa_tree_add_8_49_groupi_n_130 ,csa_tree_add_8_49_groupi_n_275);
  or csa_tree_add_8_49_groupi_g2641(csa_tree_add_8_49_groupi_n_362 ,csa_tree_add_8_49_groupi_n_79 ,csa_tree_add_8_49_groupi_n_272);
  or csa_tree_add_8_49_groupi_g2642(csa_tree_add_8_49_groupi_n_361 ,csa_tree_add_8_49_groupi_n_71 ,csa_tree_add_8_49_groupi_n_298);
  or csa_tree_add_8_49_groupi_g2643(csa_tree_add_8_49_groupi_n_360 ,csa_tree_add_8_49_groupi_n_94 ,csa_tree_add_8_49_groupi_n_296);
  or csa_tree_add_8_49_groupi_g2644(csa_tree_add_8_49_groupi_n_359 ,csa_tree_add_8_49_groupi_n_144 ,csa_tree_add_8_49_groupi_n_274);
  or csa_tree_add_8_49_groupi_g2645(csa_tree_add_8_49_groupi_n_358 ,csa_tree_add_8_49_groupi_n_92 ,csa_tree_add_8_49_groupi_n_283);
  or csa_tree_add_8_49_groupi_g2646(csa_tree_add_8_49_groupi_n_357 ,csa_tree_add_8_49_groupi_n_134 ,csa_tree_add_8_49_groupi_n_276);
  or csa_tree_add_8_49_groupi_g2647(csa_tree_add_8_49_groupi_n_356 ,csa_tree_add_8_49_groupi_n_86 ,csa_tree_add_8_49_groupi_n_273);
  or csa_tree_add_8_49_groupi_g2648(csa_tree_add_8_49_groupi_n_355 ,csa_tree_add_8_49_groupi_n_151 ,csa_tree_add_8_49_groupi_n_271);
  or csa_tree_add_8_49_groupi_g2649(csa_tree_add_8_49_groupi_n_354 ,csa_tree_add_8_49_groupi_n_96 ,csa_tree_add_8_49_groupi_n_300);
  or csa_tree_add_8_49_groupi_g2650(csa_tree_add_8_49_groupi_n_353 ,csa_tree_add_8_49_groupi_n_148 ,csa_tree_add_8_49_groupi_n_278);
  or csa_tree_add_8_49_groupi_g2651(csa_tree_add_8_49_groupi_n_352 ,csa_tree_add_8_49_groupi_n_85 ,csa_tree_add_8_49_groupi_n_270);
  or csa_tree_add_8_49_groupi_g2652(csa_tree_add_8_49_groupi_n_351 ,csa_tree_add_8_49_groupi_n_83 ,csa_tree_add_8_49_groupi_n_279);
  or csa_tree_add_8_49_groupi_g2653(csa_tree_add_8_49_groupi_n_350 ,csa_tree_add_8_49_groupi_n_67 ,csa_tree_add_8_49_groupi_n_280);
  or csa_tree_add_8_49_groupi_g2654(csa_tree_add_8_49_groupi_n_349 ,csa_tree_add_8_49_groupi_n_137 ,csa_tree_add_8_49_groupi_n_281);
  not csa_tree_add_8_49_groupi_g2655(csa_tree_add_8_49_groupi_n_315 ,csa_tree_add_8_49_groupi_n_316);
  not csa_tree_add_8_49_groupi_g2656(csa_tree_add_8_49_groupi_n_313 ,csa_tree_add_8_49_groupi_n_314);
  not csa_tree_add_8_49_groupi_g2657(csa_tree_add_8_49_groupi_n_311 ,csa_tree_add_8_49_groupi_n_312);
  not csa_tree_add_8_49_groupi_g2658(csa_tree_add_8_49_groupi_n_309 ,csa_tree_add_8_49_groupi_n_310);
  not csa_tree_add_8_49_groupi_g2659(csa_tree_add_8_49_groupi_n_307 ,csa_tree_add_8_49_groupi_n_308);
  not csa_tree_add_8_49_groupi_g2660(csa_tree_add_8_49_groupi_n_305 ,csa_tree_add_8_49_groupi_n_306);
  not csa_tree_add_8_49_groupi_g2661(csa_tree_add_8_49_groupi_n_303 ,csa_tree_add_8_49_groupi_n_304);
  not csa_tree_add_8_49_groupi_g2662(csa_tree_add_8_49_groupi_n_301 ,csa_tree_add_8_49_groupi_n_302);
  and csa_tree_add_8_49_groupi_g2663(csa_tree_add_8_49_groupi_n_300 ,n_1815 ,csa_tree_add_8_49_groupi_n_75);
  and csa_tree_add_8_49_groupi_g2664(csa_tree_add_8_49_groupi_n_299 ,n_1831 ,csa_tree_add_8_49_groupi_n_68);
  and csa_tree_add_8_49_groupi_g2665(csa_tree_add_8_49_groupi_n_298 ,n_1827 ,csa_tree_add_8_49_groupi_n_132);
  and csa_tree_add_8_49_groupi_g2666(csa_tree_add_8_49_groupi_n_297 ,n_1833 ,csa_tree_add_8_49_groupi_n_140);
  and csa_tree_add_8_49_groupi_g2667(csa_tree_add_8_49_groupi_n_296 ,n_1835 ,csa_tree_add_8_49_groupi_n_89);
  and csa_tree_add_8_49_groupi_g2668(csa_tree_add_8_49_groupi_n_295 ,n_1826 ,csa_tree_add_8_49_groupi_n_128);
  and csa_tree_add_8_49_groupi_g2669(csa_tree_add_8_49_groupi_n_294 ,n_1844 ,csa_tree_add_8_49_groupi_n_150);
  and csa_tree_add_8_49_groupi_g2670(csa_tree_add_8_49_groupi_n_293 ,n_1825 ,csa_tree_add_8_49_groupi_n_149);
  and csa_tree_add_8_49_groupi_g2671(csa_tree_add_8_49_groupi_n_292 ,n_1824 ,csa_tree_add_8_49_groupi_n_139);
  and csa_tree_add_8_49_groupi_g2672(csa_tree_add_8_49_groupi_n_291 ,n_1843 ,csa_tree_add_8_49_groupi_n_143);
  and csa_tree_add_8_49_groupi_g2673(csa_tree_add_8_49_groupi_n_290 ,n_1823 ,csa_tree_add_8_49_groupi_n_147);
  and csa_tree_add_8_49_groupi_g2674(csa_tree_add_8_49_groupi_n_289 ,n_1834 ,csa_tree_add_8_49_groupi_n_138);
  and csa_tree_add_8_49_groupi_g2675(csa_tree_add_8_49_groupi_n_288 ,n_1822 ,csa_tree_add_8_49_groupi_n_153);
  and csa_tree_add_8_49_groupi_g2676(csa_tree_add_8_49_groupi_n_287 ,n_1842 ,csa_tree_add_8_49_groupi_n_73);
  and csa_tree_add_8_49_groupi_g2677(csa_tree_add_8_49_groupi_n_286 ,n_1821 ,csa_tree_add_8_49_groupi_n_90);
  and csa_tree_add_8_49_groupi_g2678(csa_tree_add_8_49_groupi_n_285 ,n_1820 ,csa_tree_add_8_49_groupi_n_142);
  and csa_tree_add_8_49_groupi_g2679(csa_tree_add_8_49_groupi_n_284 ,n_1841 ,csa_tree_add_8_49_groupi_n_91);
  and csa_tree_add_8_49_groupi_g2680(csa_tree_add_8_49_groupi_n_283 ,n_1819 ,csa_tree_add_8_49_groupi_n_88);
  and csa_tree_add_8_49_groupi_g2681(csa_tree_add_8_49_groupi_n_282 ,n_1818 ,csa_tree_add_8_49_groupi_n_155);
  and csa_tree_add_8_49_groupi_g2682(csa_tree_add_8_49_groupi_n_281 ,n_1840 ,csa_tree_add_8_49_groupi_n_80);
  and csa_tree_add_8_49_groupi_g2683(csa_tree_add_8_49_groupi_n_280 ,in3[4] ,csa_tree_add_8_49_groupi_n_95);
  and csa_tree_add_8_49_groupi_g2684(csa_tree_add_8_49_groupi_n_279 ,n_1880 ,csa_tree_add_8_49_groupi_n_72);
  and csa_tree_add_8_49_groupi_g2685(csa_tree_add_8_49_groupi_n_278 ,n_1839 ,csa_tree_add_8_49_groupi_n_74);
  and csa_tree_add_8_49_groupi_g2686(csa_tree_add_8_49_groupi_n_277 ,n_1832 ,csa_tree_add_8_49_groupi_n_69);
  and csa_tree_add_8_49_groupi_g2687(csa_tree_add_8_49_groupi_n_276 ,n_1838 ,csa_tree_add_8_49_groupi_n_136);
  and csa_tree_add_8_49_groupi_g2688(csa_tree_add_8_49_groupi_n_275 ,n_1877 ,csa_tree_add_8_49_groupi_n_129);
  and csa_tree_add_8_49_groupi_g2689(csa_tree_add_8_49_groupi_n_274 ,n_1837 ,csa_tree_add_8_49_groupi_n_133);
  and csa_tree_add_8_49_groupi_g2690(csa_tree_add_8_49_groupi_n_273 ,n_1836 ,csa_tree_add_8_49_groupi_n_145);
  and csa_tree_add_8_49_groupi_g2691(csa_tree_add_8_49_groupi_n_272 ,n_1828 ,csa_tree_add_8_49_groupi_n_76);
  and csa_tree_add_8_49_groupi_g2692(csa_tree_add_8_49_groupi_n_271 ,n_1829 ,csa_tree_add_8_49_groupi_n_77);
  and csa_tree_add_8_49_groupi_g2693(csa_tree_add_8_49_groupi_n_270 ,n_1830 ,csa_tree_add_8_49_groupi_n_141);
  xnor csa_tree_add_8_49_groupi_g2694(csa_tree_add_8_49_groupi_n_269 ,n_1888 ,in3[11]);
  xnor csa_tree_add_8_49_groupi_g2695(csa_tree_add_8_49_groupi_n_268 ,n_1940 ,n_1876);
  xnor csa_tree_add_8_49_groupi_g2696(csa_tree_add_8_49_groupi_n_267 ,n_1901 ,in3[24]);
  xnor csa_tree_add_8_49_groupi_g2697(csa_tree_add_8_49_groupi_n_266 ,n_1898 ,in3[21]);
  xnor csa_tree_add_8_49_groupi_g2698(csa_tree_add_8_49_groupi_n_265 ,n_1894 ,in3[17]);
  xnor csa_tree_add_8_49_groupi_g2699(csa_tree_add_8_49_groupi_n_264 ,n_1892 ,in3[15]);
  xnor csa_tree_add_8_49_groupi_g2700(csa_tree_add_8_49_groupi_n_263 ,n_1903 ,in3[26]);
  xnor csa_tree_add_8_49_groupi_g2701(csa_tree_add_8_49_groupi_n_262 ,n_1900 ,in3[23]);
  xnor csa_tree_add_8_49_groupi_g2702(csa_tree_add_8_49_groupi_n_316 ,n_1915 ,n_1851);
  xnor csa_tree_add_8_49_groupi_g2703(csa_tree_add_8_49_groupi_n_314 ,n_1926 ,n_1862);
  xnor csa_tree_add_8_49_groupi_g2704(csa_tree_add_8_49_groupi_n_312 ,n_1913 ,n_1849);
  xnor csa_tree_add_8_49_groupi_g2705(csa_tree_add_8_49_groupi_n_310 ,n_1927 ,n_1863);
  xnor csa_tree_add_8_49_groupi_g2706(csa_tree_add_8_49_groupi_n_308 ,n_1918 ,n_1854);
  xnor csa_tree_add_8_49_groupi_g2707(csa_tree_add_8_49_groupi_n_306 ,n_1934 ,n_1870);
  xnor csa_tree_add_8_49_groupi_g2708(csa_tree_add_8_49_groupi_n_304 ,n_1928 ,n_1864);
  xnor csa_tree_add_8_49_groupi_g2709(csa_tree_add_8_49_groupi_n_302 ,n_1914 ,n_1850);
  not csa_tree_add_8_49_groupi_g2710(csa_tree_add_8_49_groupi_n_260 ,csa_tree_add_8_49_groupi_n_261);
  not csa_tree_add_8_49_groupi_g2711(csa_tree_add_8_49_groupi_n_258 ,csa_tree_add_8_49_groupi_n_259);
  not csa_tree_add_8_49_groupi_g2712(csa_tree_add_8_49_groupi_n_256 ,csa_tree_add_8_49_groupi_n_257);
  not csa_tree_add_8_49_groupi_g2713(csa_tree_add_8_49_groupi_n_254 ,csa_tree_add_8_49_groupi_n_255);
  not csa_tree_add_8_49_groupi_g2714(csa_tree_add_8_49_groupi_n_252 ,csa_tree_add_8_49_groupi_n_253);
  not csa_tree_add_8_49_groupi_g2715(csa_tree_add_8_49_groupi_n_250 ,csa_tree_add_8_49_groupi_n_251);
  not csa_tree_add_8_49_groupi_g2716(csa_tree_add_8_49_groupi_n_248 ,csa_tree_add_8_49_groupi_n_249);
  not csa_tree_add_8_49_groupi_g2717(csa_tree_add_8_49_groupi_n_246 ,csa_tree_add_8_49_groupi_n_247);
  not csa_tree_add_8_49_groupi_g2718(csa_tree_add_8_49_groupi_n_244 ,csa_tree_add_8_49_groupi_n_245);
  not csa_tree_add_8_49_groupi_g2719(csa_tree_add_8_49_groupi_n_242 ,csa_tree_add_8_49_groupi_n_243);
  not csa_tree_add_8_49_groupi_g2720(csa_tree_add_8_49_groupi_n_240 ,csa_tree_add_8_49_groupi_n_241);
  not csa_tree_add_8_49_groupi_g2721(csa_tree_add_8_49_groupi_n_238 ,csa_tree_add_8_49_groupi_n_239);
  not csa_tree_add_8_49_groupi_g2722(csa_tree_add_8_49_groupi_n_236 ,csa_tree_add_8_49_groupi_n_237);
  not csa_tree_add_8_49_groupi_g2723(csa_tree_add_8_49_groupi_n_234 ,csa_tree_add_8_49_groupi_n_235);
  not csa_tree_add_8_49_groupi_g2724(csa_tree_add_8_49_groupi_n_232 ,csa_tree_add_8_49_groupi_n_233);
  not csa_tree_add_8_49_groupi_g2725(csa_tree_add_8_49_groupi_n_230 ,csa_tree_add_8_49_groupi_n_231);
  not csa_tree_add_8_49_groupi_g2726(csa_tree_add_8_49_groupi_n_228 ,csa_tree_add_8_49_groupi_n_229);
  not csa_tree_add_8_49_groupi_g2727(csa_tree_add_8_49_groupi_n_226 ,csa_tree_add_8_49_groupi_n_227);
  not csa_tree_add_8_49_groupi_g2728(csa_tree_add_8_49_groupi_n_224 ,csa_tree_add_8_49_groupi_n_225);
  not csa_tree_add_8_49_groupi_g2729(csa_tree_add_8_49_groupi_n_222 ,csa_tree_add_8_49_groupi_n_223);
  not csa_tree_add_8_49_groupi_g2730(csa_tree_add_8_49_groupi_n_220 ,csa_tree_add_8_49_groupi_n_221);
  not csa_tree_add_8_49_groupi_g2731(csa_tree_add_8_49_groupi_n_218 ,csa_tree_add_8_49_groupi_n_219);
  not csa_tree_add_8_49_groupi_g2732(csa_tree_add_8_49_groupi_n_216 ,csa_tree_add_8_49_groupi_n_217);
  not csa_tree_add_8_49_groupi_g2733(csa_tree_add_8_49_groupi_n_214 ,csa_tree_add_8_49_groupi_n_215);
  xnor csa_tree_add_8_49_groupi_g2734(csa_tree_add_8_49_groupi_n_213 ,n_1877 ,n_1813);
  xnor csa_tree_add_8_49_groupi_g2735(csa_tree_add_8_49_groupi_n_212 ,n_1891 ,in3[14]);
  xnor csa_tree_add_8_49_groupi_g2736(csa_tree_add_8_49_groupi_n_211 ,n_1899 ,in3[22]);
  xnor csa_tree_add_8_49_groupi_g2737(csa_tree_add_8_49_groupi_n_210 ,n_1896 ,in3[19]);
  xnor csa_tree_add_8_49_groupi_g2738(csa_tree_add_8_49_groupi_n_209 ,n_1890 ,in3[13]);
  xnor csa_tree_add_8_49_groupi_g2739(csa_tree_add_8_49_groupi_n_208 ,n_1893 ,in3[16]);
  xnor csa_tree_add_8_49_groupi_g2740(csa_tree_add_8_49_groupi_n_207 ,n_1889 ,in3[12]);
  xnor csa_tree_add_8_49_groupi_g2741(csa_tree_add_8_49_groupi_n_206 ,n_1908 ,in3[31]);
  xnor csa_tree_add_8_49_groupi_g2742(csa_tree_add_8_49_groupi_n_205 ,n_1887 ,in3[10]);
  xnor csa_tree_add_8_49_groupi_g2743(csa_tree_add_8_49_groupi_n_204 ,n_1907 ,in3[30]);
  xnor csa_tree_add_8_49_groupi_g2744(csa_tree_add_8_49_groupi_n_203 ,n_1886 ,in3[9]);
  xnor csa_tree_add_8_49_groupi_g2745(csa_tree_add_8_49_groupi_n_202 ,n_1885 ,in3[8]);
  xnor csa_tree_add_8_49_groupi_g2746(csa_tree_add_8_49_groupi_n_201 ,n_1906 ,in3[29]);
  xnor csa_tree_add_8_49_groupi_g2747(csa_tree_add_8_49_groupi_n_200 ,n_1884 ,in3[7]);
  xnor csa_tree_add_8_49_groupi_g2748(csa_tree_add_8_49_groupi_n_199 ,n_1883 ,in3[6]);
  xnor csa_tree_add_8_49_groupi_g2749(csa_tree_add_8_49_groupi_n_198 ,n_1895 ,in3[18]);
  xnor csa_tree_add_8_49_groupi_g2750(csa_tree_add_8_49_groupi_n_197 ,n_1904 ,in3[27]);
  xnor csa_tree_add_8_49_groupi_g2751(csa_tree_add_8_49_groupi_n_196 ,n_1881 ,in3[4]);
  xnor csa_tree_add_8_49_groupi_g2752(csa_tree_add_8_49_groupi_n_195 ,n_1897 ,in3[20]);
  xnor csa_tree_add_8_49_groupi_g2753(csa_tree_add_8_49_groupi_n_194 ,n_1879 ,in3[2]);
  xnor csa_tree_add_8_49_groupi_g2754(csa_tree_add_8_49_groupi_n_193 ,n_1880 ,in3[3]);
  xnor csa_tree_add_8_49_groupi_g2755(csa_tree_add_8_49_groupi_n_192 ,n_1902 ,in3[25]);
  xnor csa_tree_add_8_49_groupi_g2756(csa_tree_add_8_49_groupi_n_191 ,n_1905 ,in3[28]);
  xnor csa_tree_add_8_49_groupi_g2757(csa_tree_add_8_49_groupi_n_190 ,n_1882 ,in3[5]);
  xnor csa_tree_add_8_49_groupi_g2758(csa_tree_add_8_49_groupi_n_261 ,n_1910 ,n_1846);
  xnor csa_tree_add_8_49_groupi_g2759(csa_tree_add_8_49_groupi_n_259 ,n_1933 ,n_1869);
  xnor csa_tree_add_8_49_groupi_g2760(csa_tree_add_8_49_groupi_n_257 ,n_1935 ,n_1871);
  xnor csa_tree_add_8_49_groupi_g2761(csa_tree_add_8_49_groupi_n_255 ,n_1912 ,n_1848);
  xnor csa_tree_add_8_49_groupi_g2762(csa_tree_add_8_49_groupi_n_253 ,n_1936 ,n_1872);
  xnor csa_tree_add_8_49_groupi_g2763(csa_tree_add_8_49_groupi_n_251 ,n_1924 ,n_1860);
  xnor csa_tree_add_8_49_groupi_g2764(csa_tree_add_8_49_groupi_n_249 ,n_1931 ,n_1867);
  xnor csa_tree_add_8_49_groupi_g2765(csa_tree_add_8_49_groupi_n_247 ,n_1921 ,n_1857);
  xnor csa_tree_add_8_49_groupi_g2766(csa_tree_add_8_49_groupi_n_245 ,n_1909 ,n_1845);
  xnor csa_tree_add_8_49_groupi_g2767(csa_tree_add_8_49_groupi_n_243 ,n_1922 ,n_1858);
  xnor csa_tree_add_8_49_groupi_g2768(csa_tree_add_8_49_groupi_n_241 ,n_1911 ,n_1847);
  xnor csa_tree_add_8_49_groupi_g2769(csa_tree_add_8_49_groupi_n_239 ,n_1917 ,n_1853);
  xnor csa_tree_add_8_49_groupi_g2770(csa_tree_add_8_49_groupi_n_237 ,n_1920 ,n_1856);
  xnor csa_tree_add_8_49_groupi_g2771(csa_tree_add_8_49_groupi_n_235 ,n_1814 ,in3[1]);
  xnor csa_tree_add_8_49_groupi_g2772(csa_tree_add_8_49_groupi_n_233 ,n_1937 ,n_1873);
  xnor csa_tree_add_8_49_groupi_g2773(csa_tree_add_8_49_groupi_n_231 ,n_1932 ,n_1868);
  xnor csa_tree_add_8_49_groupi_g2774(csa_tree_add_8_49_groupi_n_229 ,n_1930 ,n_1866);
  xnor csa_tree_add_8_49_groupi_g2775(csa_tree_add_8_49_groupi_n_227 ,n_1919 ,n_1855);
  xnor csa_tree_add_8_49_groupi_g2776(csa_tree_add_8_49_groupi_n_225 ,n_1929 ,n_1865);
  xnor csa_tree_add_8_49_groupi_g2777(csa_tree_add_8_49_groupi_n_223 ,n_1938 ,n_1874);
  xnor csa_tree_add_8_49_groupi_g2778(csa_tree_add_8_49_groupi_n_221 ,n_1939 ,n_1875);
  xnor csa_tree_add_8_49_groupi_g2779(csa_tree_add_8_49_groupi_n_219 ,n_1925 ,n_1861);
  xnor csa_tree_add_8_49_groupi_g2780(csa_tree_add_8_49_groupi_n_217 ,n_1923 ,n_1859);
  xnor csa_tree_add_8_49_groupi_g2781(csa_tree_add_8_49_groupi_n_215 ,n_1916 ,n_1852);
  not csa_tree_add_8_49_groupi_g2782(csa_tree_add_8_49_groupi_n_188 ,csa_tree_add_8_49_groupi_n_189);
  not csa_tree_add_8_49_groupi_g2783(csa_tree_add_8_49_groupi_n_186 ,csa_tree_add_8_49_groupi_n_187);
  not csa_tree_add_8_49_groupi_g2784(csa_tree_add_8_49_groupi_n_184 ,csa_tree_add_8_49_groupi_n_185);
  not csa_tree_add_8_49_groupi_g2785(csa_tree_add_8_49_groupi_n_182 ,csa_tree_add_8_49_groupi_n_183);
  not csa_tree_add_8_49_groupi_g2786(csa_tree_add_8_49_groupi_n_180 ,csa_tree_add_8_49_groupi_n_181);
  not csa_tree_add_8_49_groupi_g2787(csa_tree_add_8_49_groupi_n_178 ,csa_tree_add_8_49_groupi_n_179);
  not csa_tree_add_8_49_groupi_g2788(csa_tree_add_8_49_groupi_n_176 ,csa_tree_add_8_49_groupi_n_177);
  not csa_tree_add_8_49_groupi_g2789(csa_tree_add_8_49_groupi_n_174 ,csa_tree_add_8_49_groupi_n_175);
  not csa_tree_add_8_49_groupi_g2790(csa_tree_add_8_49_groupi_n_172 ,csa_tree_add_8_49_groupi_n_173);
  not csa_tree_add_8_49_groupi_g2791(csa_tree_add_8_49_groupi_n_170 ,csa_tree_add_8_49_groupi_n_171);
  not csa_tree_add_8_49_groupi_g2792(csa_tree_add_8_49_groupi_n_168 ,csa_tree_add_8_49_groupi_n_169);
  not csa_tree_add_8_49_groupi_g2793(csa_tree_add_8_49_groupi_n_166 ,csa_tree_add_8_49_groupi_n_167);
  not csa_tree_add_8_49_groupi_g2794(csa_tree_add_8_49_groupi_n_164 ,csa_tree_add_8_49_groupi_n_165);
  not csa_tree_add_8_49_groupi_g2795(csa_tree_add_8_49_groupi_n_162 ,csa_tree_add_8_49_groupi_n_163);
  not csa_tree_add_8_49_groupi_g2796(csa_tree_add_8_49_groupi_n_160 ,csa_tree_add_8_49_groupi_n_161);
  not csa_tree_add_8_49_groupi_g2797(csa_tree_add_8_49_groupi_n_158 ,csa_tree_add_8_49_groupi_n_159);
  and csa_tree_add_8_49_groupi_g2798(csa_tree_add_8_49_groupi_n_157 ,in3[30] ,n_1907);
  and csa_tree_add_8_49_groupi_g2799(csa_tree_add_8_49_groupi_n_156 ,in3[21] ,n_1898);
  or csa_tree_add_8_49_groupi_g2800(csa_tree_add_8_49_groupi_n_155 ,in3[5] ,n_1882);
  and csa_tree_add_8_49_groupi_g2801(csa_tree_add_8_49_groupi_n_154 ,in3[13] ,n_1890);
  or csa_tree_add_8_49_groupi_g2802(csa_tree_add_8_49_groupi_n_153 ,in3[9] ,n_1886);
  and csa_tree_add_8_49_groupi_g2803(csa_tree_add_8_49_groupi_n_152 ,in3[9] ,n_1886);
  and csa_tree_add_8_49_groupi_g2804(csa_tree_add_8_49_groupi_n_151 ,in3[16] ,n_1893);
  or csa_tree_add_8_49_groupi_g2805(csa_tree_add_8_49_groupi_n_150 ,in3[31] ,n_1908);
  or csa_tree_add_8_49_groupi_g2806(csa_tree_add_8_49_groupi_n_149 ,in3[12] ,n_1889);
  and csa_tree_add_8_49_groupi_g2807(csa_tree_add_8_49_groupi_n_148 ,in3[26] ,n_1903);
  or csa_tree_add_8_49_groupi_g2808(csa_tree_add_8_49_groupi_n_147 ,in3[10] ,n_1887);
  and csa_tree_add_8_49_groupi_g2809(csa_tree_add_8_49_groupi_n_146 ,in3[12] ,n_1889);
  or csa_tree_add_8_49_groupi_g2810(csa_tree_add_8_49_groupi_n_145 ,in3[23] ,n_1900);
  and csa_tree_add_8_49_groupi_g2811(csa_tree_add_8_49_groupi_n_144 ,in3[24] ,n_1901);
  or csa_tree_add_8_49_groupi_g2812(csa_tree_add_8_49_groupi_n_143 ,in3[30] ,n_1907);
  or csa_tree_add_8_49_groupi_g2813(csa_tree_add_8_49_groupi_n_142 ,in3[7] ,n_1884);
  or csa_tree_add_8_49_groupi_g2814(csa_tree_add_8_49_groupi_n_141 ,in3[17] ,n_1894);
  or csa_tree_add_8_49_groupi_g2815(csa_tree_add_8_49_groupi_n_140 ,in3[20] ,n_1897);
  or csa_tree_add_8_49_groupi_g2816(csa_tree_add_8_49_groupi_n_139 ,in3[11] ,n_1888);
  or csa_tree_add_8_49_groupi_g2817(csa_tree_add_8_49_groupi_n_138 ,in3[21] ,n_1898);
  and csa_tree_add_8_49_groupi_g2818(csa_tree_add_8_49_groupi_n_137 ,in3[27] ,n_1904);
  or csa_tree_add_8_49_groupi_g2819(csa_tree_add_8_49_groupi_n_136 ,in3[25] ,n_1902);
  and csa_tree_add_8_49_groupi_g2820(csa_tree_add_8_49_groupi_n_135 ,in3[11] ,n_1888);
  and csa_tree_add_8_49_groupi_g2821(csa_tree_add_8_49_groupi_n_134 ,in3[25] ,n_1902);
  or csa_tree_add_8_49_groupi_g2822(csa_tree_add_8_49_groupi_n_133 ,in3[24] ,n_1901);
  or csa_tree_add_8_49_groupi_g2823(csa_tree_add_8_49_groupi_n_132 ,in3[14] ,n_1891);
  and csa_tree_add_8_49_groupi_g2824(csa_tree_add_8_49_groupi_n_131 ,in3[31] ,n_1908);
  and csa_tree_add_8_49_groupi_g2825(csa_tree_add_8_49_groupi_n_130 ,in3[0] ,n_1813);
  or csa_tree_add_8_49_groupi_g2826(csa_tree_add_8_49_groupi_n_129 ,in3[0] ,n_1813);
  or csa_tree_add_8_49_groupi_g2827(csa_tree_add_8_49_groupi_n_128 ,in3[13] ,n_1890);
  or csa_tree_add_8_49_groupi_g2828(csa_tree_add_8_49_groupi_n_127 ,csa_tree_add_8_49_groupi_n_19 ,csa_tree_add_8_49_groupi_n_38);
  or csa_tree_add_8_49_groupi_g2829(csa_tree_add_8_49_groupi_n_189 ,csa_tree_add_8_49_groupi_n_60 ,csa_tree_add_8_49_groupi_n_17);
  or csa_tree_add_8_49_groupi_g2830(csa_tree_add_8_49_groupi_n_187 ,csa_tree_add_8_49_groupi_n_61 ,csa_tree_add_8_49_groupi_n_18);
  or csa_tree_add_8_49_groupi_g2831(csa_tree_add_8_49_groupi_n_185 ,csa_tree_add_8_49_groupi_n_22 ,csa_tree_add_8_49_groupi_n_42);
  or csa_tree_add_8_49_groupi_g2832(csa_tree_add_8_49_groupi_n_183 ,csa_tree_add_8_49_groupi_n_41 ,csa_tree_add_8_49_groupi_n_44);
  or csa_tree_add_8_49_groupi_g2833(csa_tree_add_8_49_groupi_n_181 ,csa_tree_add_8_49_groupi_n_49 ,csa_tree_add_8_49_groupi_n_10);
  or csa_tree_add_8_49_groupi_g2834(csa_tree_add_8_49_groupi_n_179 ,csa_tree_add_8_49_groupi_n_57 ,csa_tree_add_8_49_groupi_n_58);
  or csa_tree_add_8_49_groupi_g2835(csa_tree_add_8_49_groupi_n_177 ,csa_tree_add_8_49_groupi_n_56 ,csa_tree_add_8_49_groupi_n_62);
  or csa_tree_add_8_49_groupi_g2836(csa_tree_add_8_49_groupi_n_175 ,csa_tree_add_8_49_groupi_n_45 ,csa_tree_add_8_49_groupi_n_20);
  or csa_tree_add_8_49_groupi_g2837(csa_tree_add_8_49_groupi_n_173 ,csa_tree_add_8_49_groupi_n_11 ,csa_tree_add_8_49_groupi_n_2);
  or csa_tree_add_8_49_groupi_g2838(csa_tree_add_8_49_groupi_n_171 ,csa_tree_add_8_49_groupi_n_46 ,csa_tree_add_8_49_groupi_n_27);
  or csa_tree_add_8_49_groupi_g2839(csa_tree_add_8_49_groupi_n_169 ,csa_tree_add_8_49_groupi_n_23 ,csa_tree_add_8_49_groupi_n_15);
  or csa_tree_add_8_49_groupi_g2840(csa_tree_add_8_49_groupi_n_167 ,csa_tree_add_8_49_groupi_n_4 ,csa_tree_add_8_49_groupi_n_34);
  or csa_tree_add_8_49_groupi_g2841(csa_tree_add_8_49_groupi_n_165 ,csa_tree_add_8_49_groupi_n_24 ,csa_tree_add_8_49_groupi_n_53);
  or csa_tree_add_8_49_groupi_g2842(csa_tree_add_8_49_groupi_n_163 ,csa_tree_add_8_49_groupi_n_6 ,csa_tree_add_8_49_groupi_n_43);
  or csa_tree_add_8_49_groupi_g2843(csa_tree_add_8_49_groupi_n_161 ,csa_tree_add_8_49_groupi_n_33 ,csa_tree_add_8_49_groupi_n_48);
  or csa_tree_add_8_49_groupi_g2844(csa_tree_add_8_49_groupi_n_159 ,csa_tree_add_8_49_groupi_n_3 ,csa_tree_add_8_49_groupi_n_16);
  not csa_tree_add_8_49_groupi_g2845(csa_tree_add_8_49_groupi_n_125 ,csa_tree_add_8_49_groupi_n_126);
  not csa_tree_add_8_49_groupi_g2846(csa_tree_add_8_49_groupi_n_123 ,csa_tree_add_8_49_groupi_n_124);
  not csa_tree_add_8_49_groupi_g2847(csa_tree_add_8_49_groupi_n_121 ,csa_tree_add_8_49_groupi_n_122);
  not csa_tree_add_8_49_groupi_g2848(csa_tree_add_8_49_groupi_n_119 ,csa_tree_add_8_49_groupi_n_120);
  not csa_tree_add_8_49_groupi_g2849(csa_tree_add_8_49_groupi_n_117 ,csa_tree_add_8_49_groupi_n_118);
  not csa_tree_add_8_49_groupi_g2850(csa_tree_add_8_49_groupi_n_115 ,csa_tree_add_8_49_groupi_n_116);
  not csa_tree_add_8_49_groupi_g2851(csa_tree_add_8_49_groupi_n_113 ,csa_tree_add_8_49_groupi_n_114);
  not csa_tree_add_8_49_groupi_g2852(csa_tree_add_8_49_groupi_n_111 ,csa_tree_add_8_49_groupi_n_112);
  not csa_tree_add_8_49_groupi_g2853(csa_tree_add_8_49_groupi_n_109 ,csa_tree_add_8_49_groupi_n_110);
  not csa_tree_add_8_49_groupi_g2854(csa_tree_add_8_49_groupi_n_107 ,csa_tree_add_8_49_groupi_n_108);
  not csa_tree_add_8_49_groupi_g2855(csa_tree_add_8_49_groupi_n_105 ,csa_tree_add_8_49_groupi_n_106);
  not csa_tree_add_8_49_groupi_g2856(csa_tree_add_8_49_groupi_n_103 ,csa_tree_add_8_49_groupi_n_104);
  not csa_tree_add_8_49_groupi_g2857(csa_tree_add_8_49_groupi_n_101 ,csa_tree_add_8_49_groupi_n_102);
  not csa_tree_add_8_49_groupi_g2858(csa_tree_add_8_49_groupi_n_99 ,csa_tree_add_8_49_groupi_n_100);
  not csa_tree_add_8_49_groupi_g2859(csa_tree_add_8_49_groupi_n_97 ,csa_tree_add_8_49_groupi_n_98);
  and csa_tree_add_8_49_groupi_g2860(csa_tree_add_8_49_groupi_n_96 ,in3[2] ,n_1879);
  or csa_tree_add_8_49_groupi_g2861(csa_tree_add_8_49_groupi_n_95 ,n_1881 ,n_1817);
  and csa_tree_add_8_49_groupi_g2862(csa_tree_add_8_49_groupi_n_94 ,in3[22] ,n_1899);
  and csa_tree_add_8_49_groupi_g2863(csa_tree_add_8_49_groupi_n_93 ,in3[8] ,n_1885);
  and csa_tree_add_8_49_groupi_g2864(csa_tree_add_8_49_groupi_n_92 ,in3[6] ,n_1883);
  or csa_tree_add_8_49_groupi_g2865(csa_tree_add_8_49_groupi_n_91 ,in3[28] ,n_1905);
  or csa_tree_add_8_49_groupi_g2866(csa_tree_add_8_49_groupi_n_90 ,in3[8] ,n_1885);
  or csa_tree_add_8_49_groupi_g2867(csa_tree_add_8_49_groupi_n_89 ,in3[22] ,n_1899);
  or csa_tree_add_8_49_groupi_g2868(csa_tree_add_8_49_groupi_n_88 ,in3[6] ,n_1883);
  and csa_tree_add_8_49_groupi_g2869(csa_tree_add_8_49_groupi_n_87 ,in3[10] ,n_1887);
  and csa_tree_add_8_49_groupi_g2870(csa_tree_add_8_49_groupi_n_86 ,in3[23] ,n_1900);
  and csa_tree_add_8_49_groupi_g2871(csa_tree_add_8_49_groupi_n_85 ,in3[17] ,n_1894);
  and csa_tree_add_8_49_groupi_g2872(csa_tree_add_8_49_groupi_n_84 ,in3[5] ,n_1882);
  and csa_tree_add_8_49_groupi_g2873(csa_tree_add_8_49_groupi_n_83 ,in3[3] ,n_1816);
  and csa_tree_add_8_49_groupi_g2874(csa_tree_add_8_49_groupi_n_82 ,in3[19] ,n_1896);
  and csa_tree_add_8_49_groupi_g2875(csa_tree_add_8_49_groupi_n_81 ,in3[18] ,n_1895);
  or csa_tree_add_8_49_groupi_g2876(csa_tree_add_8_49_groupi_n_80 ,in3[27] ,n_1904);
  and csa_tree_add_8_49_groupi_g2877(csa_tree_add_8_49_groupi_n_79 ,in3[15] ,n_1892);
  and csa_tree_add_8_49_groupi_g2878(csa_tree_add_8_49_groupi_n_78 ,in3[29] ,n_1906);
  or csa_tree_add_8_49_groupi_g2879(csa_tree_add_8_49_groupi_n_77 ,in3[16] ,n_1893);
  or csa_tree_add_8_49_groupi_g2880(csa_tree_add_8_49_groupi_n_76 ,in3[15] ,n_1892);
  or csa_tree_add_8_49_groupi_g2881(csa_tree_add_8_49_groupi_n_75 ,in3[2] ,n_1879);
  or csa_tree_add_8_49_groupi_g2882(csa_tree_add_8_49_groupi_n_74 ,in3[26] ,n_1903);
  or csa_tree_add_8_49_groupi_g2883(csa_tree_add_8_49_groupi_n_73 ,in3[29] ,n_1906);
  or csa_tree_add_8_49_groupi_g2884(csa_tree_add_8_49_groupi_n_72 ,in3[3] ,n_1816);
  and csa_tree_add_8_49_groupi_g2885(csa_tree_add_8_49_groupi_n_71 ,in3[14] ,n_1891);
  and csa_tree_add_8_49_groupi_g2886(csa_tree_add_8_49_groupi_n_70 ,in3[7] ,n_1884);
  or csa_tree_add_8_49_groupi_g2887(csa_tree_add_8_49_groupi_n_69 ,in3[19] ,n_1896);
  or csa_tree_add_8_49_groupi_g2888(csa_tree_add_8_49_groupi_n_68 ,in3[18] ,n_1895);
  and csa_tree_add_8_49_groupi_g2889(csa_tree_add_8_49_groupi_n_67 ,n_1881 ,n_1817);
  and csa_tree_add_8_49_groupi_g2890(csa_tree_add_8_49_groupi_n_66 ,in3[20] ,n_1897);
  and csa_tree_add_8_49_groupi_g2891(csa_tree_add_8_49_groupi_n_65 ,in3[28] ,n_1905);
  or csa_tree_add_8_49_groupi_g2892(csa_tree_add_8_49_groupi_n_126 ,csa_tree_add_8_49_groupi_n_54 ,csa_tree_add_8_49_groupi_n_63);
  or csa_tree_add_8_49_groupi_g2893(csa_tree_add_8_49_groupi_n_124 ,csa_tree_add_8_49_groupi_n_39 ,csa_tree_add_8_49_groupi_n_12);
  or csa_tree_add_8_49_groupi_g2894(csa_tree_add_8_49_groupi_n_122 ,csa_tree_add_8_49_groupi_n_26 ,csa_tree_add_8_49_groupi_n_52);
  or csa_tree_add_8_49_groupi_g2895(csa_tree_add_8_49_groupi_n_120 ,csa_tree_add_8_49_groupi_n_31 ,csa_tree_add_8_49_groupi_n_21);
  or csa_tree_add_8_49_groupi_g2896(csa_tree_add_8_49_groupi_n_118 ,csa_tree_add_8_49_groupi_n_40 ,csa_tree_add_8_49_groupi_n_14);
  or csa_tree_add_8_49_groupi_g2897(csa_tree_add_8_49_groupi_n_116 ,csa_tree_add_8_49_groupi_n_36 ,csa_tree_add_8_49_groupi_n_32);
  or csa_tree_add_8_49_groupi_g2898(csa_tree_add_8_49_groupi_n_114 ,csa_tree_add_8_49_groupi_n_64 ,csa_tree_add_8_49_groupi_n_55);
  or csa_tree_add_8_49_groupi_g2899(csa_tree_add_8_49_groupi_n_112 ,csa_tree_add_8_49_groupi_n_1 ,csa_tree_add_8_49_groupi_n_7);
  or csa_tree_add_8_49_groupi_g2900(csa_tree_add_8_49_groupi_n_110 ,csa_tree_add_8_49_groupi_n_25 ,csa_tree_add_8_49_groupi_n_30);
  or csa_tree_add_8_49_groupi_g2901(csa_tree_add_8_49_groupi_n_108 ,csa_tree_add_8_49_groupi_n_35 ,csa_tree_add_8_49_groupi_n_37);
  or csa_tree_add_8_49_groupi_g2902(csa_tree_add_8_49_groupi_n_106 ,csa_tree_add_8_49_groupi_n_5 ,csa_tree_add_8_49_groupi_n_59);
  or csa_tree_add_8_49_groupi_g2903(csa_tree_add_8_49_groupi_n_104 ,csa_tree_add_8_49_groupi_n_29 ,csa_tree_add_8_49_groupi_n_51);
  or csa_tree_add_8_49_groupi_g2904(csa_tree_add_8_49_groupi_n_102 ,csa_tree_add_8_49_groupi_n_47 ,csa_tree_add_8_49_groupi_n_8);
  or csa_tree_add_8_49_groupi_g2905(csa_tree_add_8_49_groupi_n_100 ,csa_tree_add_8_49_groupi_n_13 ,csa_tree_add_8_49_groupi_n_9);
  or csa_tree_add_8_49_groupi_g2906(csa_tree_add_8_49_groupi_n_98 ,csa_tree_add_8_49_groupi_n_50 ,csa_tree_add_8_49_groupi_n_28);
  not csa_tree_add_8_49_groupi_g2907(csa_tree_add_8_49_groupi_n_64 ,n_1919);
  not csa_tree_add_8_49_groupi_g2908(csa_tree_add_8_49_groupi_n_63 ,n_1856);
  not csa_tree_add_8_49_groupi_g2909(csa_tree_add_8_49_groupi_n_62 ,n_1859);
  not csa_tree_add_8_49_groupi_g2910(csa_tree_add_8_49_groupi_n_61 ,n_1915);
  not csa_tree_add_8_49_groupi_g2911(csa_tree_add_8_49_groupi_n_60 ,n_1927);
  not csa_tree_add_8_49_groupi_g2912(csa_tree_add_8_49_groupi_n_59 ,n_1866);
  not csa_tree_add_8_49_groupi_g2913(csa_tree_add_8_49_groupi_n_58 ,n_1868);
  not csa_tree_add_8_49_groupi_g2914(csa_tree_add_8_49_groupi_n_57 ,n_1932);
  not csa_tree_add_8_49_groupi_g2915(csa_tree_add_8_49_groupi_n_56 ,n_1923);
  not csa_tree_add_8_49_groupi_g2916(csa_tree_add_8_49_groupi_n_55 ,n_1855);
  not csa_tree_add_8_49_groupi_g2917(csa_tree_add_8_49_groupi_n_54 ,n_1920);
  not csa_tree_add_8_49_groupi_g2918(csa_tree_add_8_49_groupi_n_53 ,n_1867);
  not csa_tree_add_8_49_groupi_g2919(csa_tree_add_8_49_groupi_n_52 ,n_1853);
  not csa_tree_add_8_49_groupi_g2920(csa_tree_add_8_49_groupi_n_51 ,n_1852);
  not csa_tree_add_8_49_groupi_g2921(csa_tree_add_8_49_groupi_n_50 ,n_1918);
  not csa_tree_add_8_49_groupi_g2922(csa_tree_add_8_49_groupi_n_49 ,n_1936);
  not csa_tree_add_8_49_groupi_g2923(csa_tree_add_8_49_groupi_n_48 ,n_1845);
  not csa_tree_add_8_49_groupi_g2924(csa_tree_add_8_49_groupi_n_47 ,n_1910);
  not csa_tree_add_8_49_groupi_g2925(csa_tree_add_8_49_groupi_n_46 ,n_1926);
  not csa_tree_add_8_49_groupi_g2926(csa_tree_add_8_49_groupi_n_45 ,n_1911);
  not csa_tree_add_8_49_groupi_g2927(csa_tree_add_8_49_groupi_n_44 ,n_1857);
  not csa_tree_add_8_49_groupi_g2928(csa_tree_add_8_49_groupi_n_43 ,n_1870);
  not csa_tree_add_8_49_groupi_g2929(csa_tree_add_8_49_groupi_n_42 ,n_1873);
  not csa_tree_add_8_49_groupi_g2930(csa_tree_add_8_49_groupi_n_41 ,n_1921);
  not csa_tree_add_8_49_groupi_g2931(csa_tree_add_8_49_groupi_n_40 ,n_1935);
  not csa_tree_add_8_49_groupi_g2932(csa_tree_add_8_49_groupi_n_39 ,n_1933);
  not csa_tree_add_8_49_groupi_g2933(csa_tree_add_8_49_groupi_n_38 ,n_1875);
  not csa_tree_add_8_49_groupi_g2934(csa_tree_add_8_49_groupi_n_37 ,n_1858);
  not csa_tree_add_8_49_groupi_g2935(csa_tree_add_8_49_groupi_n_36 ,n_1928);
  not csa_tree_add_8_49_groupi_g2936(csa_tree_add_8_49_groupi_n_35 ,n_1922);
  not csa_tree_add_8_49_groupi_g2937(csa_tree_add_8_49_groupi_n_34 ,n_1850);
  not csa_tree_add_8_49_groupi_g2938(csa_tree_add_8_49_groupi_n_33 ,n_1909);
  not csa_tree_add_8_49_groupi_g2939(csa_tree_add_8_49_groupi_n_32 ,n_1864);
  not csa_tree_add_8_49_groupi_g2940(csa_tree_add_8_49_groupi_n_31 ,n_1913);
  not csa_tree_add_8_49_groupi_g2941(csa_tree_add_8_49_groupi_n_30 ,n_1865);
  not csa_tree_add_8_49_groupi_g2942(csa_tree_add_8_49_groupi_n_29 ,n_1916);
  not csa_tree_add_8_49_groupi_g2943(csa_tree_add_8_49_groupi_n_28 ,n_1854);
  not csa_tree_add_8_49_groupi_g2944(csa_tree_add_8_49_groupi_n_27 ,n_1862);
  not csa_tree_add_8_49_groupi_g2945(csa_tree_add_8_49_groupi_n_26 ,n_1917);
  not csa_tree_add_8_49_groupi_g2946(csa_tree_add_8_49_groupi_n_25 ,n_1929);
  not csa_tree_add_8_49_groupi_g2947(csa_tree_add_8_49_groupi_n_24 ,n_1931);
  not csa_tree_add_8_49_groupi_g2948(csa_tree_add_8_49_groupi_n_23 ,n_1924);
  not csa_tree_add_8_49_groupi_g2949(csa_tree_add_8_49_groupi_n_22 ,n_1937);
  not csa_tree_add_8_49_groupi_g2950(csa_tree_add_8_49_groupi_n_21 ,n_1849);
  not csa_tree_add_8_49_groupi_g2951(csa_tree_add_8_49_groupi_n_20 ,n_1847);
  not csa_tree_add_8_49_groupi_g2952(csa_tree_add_8_49_groupi_n_19 ,n_1939);
  not csa_tree_add_8_49_groupi_g2953(csa_tree_add_8_49_groupi_n_18 ,n_1851);
  not csa_tree_add_8_49_groupi_g2954(csa_tree_add_8_49_groupi_n_17 ,n_1863);
  not csa_tree_add_8_49_groupi_g2955(csa_tree_add_8_49_groupi_n_16 ,n_1874);
  not csa_tree_add_8_49_groupi_g2956(csa_tree_add_8_49_groupi_n_15 ,n_1860);
  not csa_tree_add_8_49_groupi_g2957(csa_tree_add_8_49_groupi_n_14 ,n_1871);
  not csa_tree_add_8_49_groupi_g2958(csa_tree_add_8_49_groupi_n_13 ,n_1912);
  not csa_tree_add_8_49_groupi_g2959(csa_tree_add_8_49_groupi_n_12 ,n_1869);
  not csa_tree_add_8_49_groupi_g2960(csa_tree_add_8_49_groupi_n_11 ,in3[1]);
  not csa_tree_add_8_49_groupi_g2961(csa_tree_add_8_49_groupi_n_10 ,n_1872);
  not csa_tree_add_8_49_groupi_g2962(csa_tree_add_8_49_groupi_n_9 ,n_1848);
  not csa_tree_add_8_49_groupi_g2963(csa_tree_add_8_49_groupi_n_8 ,n_1846);
  not csa_tree_add_8_49_groupi_g2964(csa_tree_add_8_49_groupi_n_7 ,n_1861);
  not csa_tree_add_8_49_groupi_g2965(csa_tree_add_8_49_groupi_n_6 ,n_1934);
  not csa_tree_add_8_49_groupi_g2966(csa_tree_add_8_49_groupi_n_5 ,n_1930);
  not csa_tree_add_8_49_groupi_g2967(csa_tree_add_8_49_groupi_n_4 ,n_1914);
  not csa_tree_add_8_49_groupi_g2968(csa_tree_add_8_49_groupi_n_3 ,n_1938);
  not csa_tree_add_8_49_groupi_g2969(csa_tree_add_8_49_groupi_n_2 ,n_1814);
  not csa_tree_add_8_49_groupi_g2970(csa_tree_add_8_49_groupi_n_1 ,n_1925);
  not csa_tree_add_8_49_groupi_g2971(csa_tree_add_8_49_groupi_n_0 ,n_1878);

endmodule

module top(in1, in2, in3, out1);

  input [2:0] in1;

  input [3:0] in2;

  input [8:0] in3;

  output out1;
  wire [2:0] in1;
  wire [3:0] in2;
  wire [8:0] in3;
  wire out1;
  wire csa_tree_lt_8_21_groupi_n_0, csa_tree_lt_8_21_groupi_n_1, csa_tree_lt_8_21_groupi_n_2, csa_tree_lt_8_21_groupi_n_3, csa_tree_lt_8_21_groupi_n_4, csa_tree_lt_8_21_groupi_n_5, csa_tree_lt_8_21_groupi_n_6, csa_tree_lt_8_21_groupi_n_7;
  wire csa_tree_lt_8_21_groupi_n_8, csa_tree_lt_8_21_groupi_n_9, csa_tree_lt_8_21_groupi_n_10, csa_tree_lt_8_21_groupi_n_11, csa_tree_lt_8_21_groupi_n_12, csa_tree_lt_8_21_groupi_n_13, csa_tree_lt_8_21_groupi_n_14, csa_tree_lt_8_21_groupi_n_15;
  wire csa_tree_lt_8_21_groupi_n_16, csa_tree_lt_8_21_groupi_n_17, csa_tree_lt_8_21_groupi_n_18, csa_tree_lt_8_21_groupi_n_19, csa_tree_lt_8_21_groupi_n_20, csa_tree_lt_8_21_groupi_n_21, csa_tree_lt_8_21_groupi_n_22, csa_tree_lt_8_21_groupi_n_23;
  wire csa_tree_lt_8_21_groupi_n_24, csa_tree_lt_8_21_groupi_n_25, csa_tree_lt_8_21_groupi_n_26, csa_tree_lt_8_21_groupi_n_27, csa_tree_lt_8_21_groupi_n_28, csa_tree_lt_8_21_groupi_n_29, csa_tree_lt_8_21_groupi_n_30, csa_tree_lt_8_21_groupi_n_31;
  wire csa_tree_lt_8_21_groupi_n_32, csa_tree_lt_8_21_groupi_n_33, csa_tree_lt_8_21_groupi_n_34, csa_tree_lt_8_21_groupi_n_35, csa_tree_lt_8_21_groupi_n_36, csa_tree_lt_8_21_groupi_n_37, csa_tree_lt_8_21_groupi_n_38, csa_tree_lt_8_21_groupi_n_39;
  wire csa_tree_lt_8_21_groupi_n_40, csa_tree_lt_8_21_groupi_n_41, csa_tree_lt_8_21_groupi_n_42, csa_tree_lt_8_21_groupi_n_43, csa_tree_lt_8_21_groupi_n_44, csa_tree_lt_8_21_groupi_n_45, csa_tree_lt_8_21_groupi_n_46, csa_tree_lt_8_21_groupi_n_47;
  wire csa_tree_lt_8_21_groupi_n_48, csa_tree_lt_8_21_groupi_n_49, csa_tree_lt_8_21_groupi_n_50, csa_tree_lt_8_21_groupi_n_51, csa_tree_lt_8_21_groupi_n_52, csa_tree_lt_8_21_groupi_n_53, csa_tree_lt_8_21_groupi_n_54, csa_tree_lt_8_21_groupi_n_55;
  wire csa_tree_lt_8_21_groupi_n_56, csa_tree_lt_8_21_groupi_n_57, csa_tree_lt_8_21_groupi_n_58, csa_tree_lt_8_21_groupi_n_59, csa_tree_lt_8_21_groupi_n_60, csa_tree_lt_8_21_groupi_n_61, csa_tree_lt_8_21_groupi_n_62, csa_tree_lt_8_21_groupi_n_63;
  wire csa_tree_lt_8_21_groupi_n_64;
  and csa_tree_lt_8_21_groupi_g428__2398(out1 ,csa_tree_lt_8_21_groupi_n_63 ,csa_tree_lt_8_21_groupi_n_64);
  or csa_tree_lt_8_21_groupi_g429__5107(csa_tree_lt_8_21_groupi_n_64 ,csa_tree_lt_8_21_groupi_n_35 ,csa_tree_lt_8_21_groupi_n_62);
  nor csa_tree_lt_8_21_groupi_g430__6260(csa_tree_lt_8_21_groupi_n_63 ,csa_tree_lt_8_21_groupi_n_15 ,csa_tree_lt_8_21_groupi_n_60);
  or csa_tree_lt_8_21_groupi_g431__4319(csa_tree_lt_8_21_groupi_n_62 ,csa_tree_lt_8_21_groupi_n_42 ,csa_tree_lt_8_21_groupi_n_61);
  or csa_tree_lt_8_21_groupi_g432__8428(csa_tree_lt_8_21_groupi_n_61 ,csa_tree_lt_8_21_groupi_n_34 ,csa_tree_lt_8_21_groupi_n_59);
  or csa_tree_lt_8_21_groupi_g433__5526(csa_tree_lt_8_21_groupi_n_60 ,csa_tree_lt_8_21_groupi_n_37 ,csa_tree_lt_8_21_groupi_n_58);
  nor csa_tree_lt_8_21_groupi_g434__6783(csa_tree_lt_8_21_groupi_n_59 ,csa_tree_lt_8_21_groupi_n_53 ,csa_tree_lt_8_21_groupi_n_57);
  nor csa_tree_lt_8_21_groupi_g435__3680(csa_tree_lt_8_21_groupi_n_58 ,csa_tree_lt_8_21_groupi_n_27 ,csa_tree_lt_8_21_groupi_n_56);
  or csa_tree_lt_8_21_groupi_g436__1617(csa_tree_lt_8_21_groupi_n_57 ,csa_tree_lt_8_21_groupi_n_47 ,csa_tree_lt_8_21_groupi_n_54);
  nor csa_tree_lt_8_21_groupi_g437__2802(csa_tree_lt_8_21_groupi_n_56 ,csa_tree_lt_8_21_groupi_n_13 ,csa_tree_lt_8_21_groupi_n_55);
  or csa_tree_lt_8_21_groupi_g438__1705(csa_tree_lt_8_21_groupi_n_55 ,csa_tree_lt_8_21_groupi_n_38 ,csa_tree_lt_8_21_groupi_n_51);
  nor csa_tree_lt_8_21_groupi_g439__5122(csa_tree_lt_8_21_groupi_n_54 ,csa_tree_lt_8_21_groupi_n_12 ,csa_tree_lt_8_21_groupi_n_52);
  nor csa_tree_lt_8_21_groupi_g440__8246(csa_tree_lt_8_21_groupi_n_53 ,in1[0] ,csa_tree_lt_8_21_groupi_n_48);
  or csa_tree_lt_8_21_groupi_g441__7098(csa_tree_lt_8_21_groupi_n_52 ,csa_tree_lt_8_21_groupi_n_33 ,csa_tree_lt_8_21_groupi_n_50);
  nor csa_tree_lt_8_21_groupi_g442__6131(csa_tree_lt_8_21_groupi_n_51 ,csa_tree_lt_8_21_groupi_n_26 ,csa_tree_lt_8_21_groupi_n_49);
  or csa_tree_lt_8_21_groupi_g443__1881(csa_tree_lt_8_21_groupi_n_50 ,csa_tree_lt_8_21_groupi_n_46 ,csa_tree_lt_8_21_groupi_n_44);
  nor csa_tree_lt_8_21_groupi_g444__5115(csa_tree_lt_8_21_groupi_n_49 ,csa_tree_lt_8_21_groupi_n_31 ,csa_tree_lt_8_21_groupi_n_45);
  or csa_tree_lt_8_21_groupi_g445__7482(csa_tree_lt_8_21_groupi_n_48 ,csa_tree_lt_8_21_groupi_n_40 ,csa_tree_lt_8_21_groupi_n_44);
  nor csa_tree_lt_8_21_groupi_g446__4733(csa_tree_lt_8_21_groupi_n_47 ,csa_tree_lt_8_21_groupi_n_36 ,csa_tree_lt_8_21_groupi_n_41);
  and csa_tree_lt_8_21_groupi_g447__6161(csa_tree_lt_8_21_groupi_n_46 ,in1[0] ,csa_tree_lt_8_21_groupi_n_40);
  nor csa_tree_lt_8_21_groupi_g448__9315(csa_tree_lt_8_21_groupi_n_45 ,csa_tree_lt_8_21_groupi_n_28 ,csa_tree_lt_8_21_groupi_n_43);
  and csa_tree_lt_8_21_groupi_g449__9945(csa_tree_lt_8_21_groupi_n_44 ,csa_tree_lt_8_21_groupi_n_36 ,csa_tree_lt_8_21_groupi_n_41);
  or csa_tree_lt_8_21_groupi_g450__2883(csa_tree_lt_8_21_groupi_n_43 ,csa_tree_lt_8_21_groupi_n_34 ,csa_tree_lt_8_21_groupi_n_39);
  and csa_tree_lt_8_21_groupi_g451__2346(csa_tree_lt_8_21_groupi_n_42 ,csa_tree_lt_8_21_groupi_n_28 ,csa_tree_lt_8_21_groupi_n_39);
  xnor csa_tree_lt_8_21_groupi_g452__1666(csa_tree_lt_8_21_groupi_n_41 ,csa_tree_lt_8_21_groupi_n_24 ,in3[2]);
  xnor csa_tree_lt_8_21_groupi_g453__7410(csa_tree_lt_8_21_groupi_n_40 ,csa_tree_lt_8_21_groupi_n_23 ,in3[1]);
  and csa_tree_lt_8_21_groupi_g454__6417(csa_tree_lt_8_21_groupi_n_39 ,csa_tree_lt_8_21_groupi_n_20 ,csa_tree_lt_8_21_groupi_n_29);
  and csa_tree_lt_8_21_groupi_g455__5477(csa_tree_lt_8_21_groupi_n_38 ,in3[4] ,csa_tree_lt_8_21_groupi_n_30);
  and csa_tree_lt_8_21_groupi_g456__2398(csa_tree_lt_8_21_groupi_n_37 ,in3[6] ,csa_tree_lt_8_21_groupi_n_32);
  and csa_tree_lt_8_21_groupi_g457__5107(csa_tree_lt_8_21_groupi_n_36 ,csa_tree_lt_8_21_groupi_n_14 ,csa_tree_lt_8_21_groupi_n_25);
  or csa_tree_lt_8_21_groupi_g458__6260(csa_tree_lt_8_21_groupi_n_35 ,csa_tree_lt_8_21_groupi_n_27 ,csa_tree_lt_8_21_groupi_n_26);
  nor csa_tree_lt_8_21_groupi_g459__4319(csa_tree_lt_8_21_groupi_n_33 ,in2[0] ,csa_tree_lt_8_21_groupi_n_11);
  nor csa_tree_lt_8_21_groupi_g460__8428(csa_tree_lt_8_21_groupi_n_32 ,in3[7] ,csa_tree_lt_8_21_groupi_n_22);
  nor csa_tree_lt_8_21_groupi_g461__5526(csa_tree_lt_8_21_groupi_n_31 ,in3[4] ,csa_tree_lt_8_21_groupi_n_16);
  nor csa_tree_lt_8_21_groupi_g462__6783(csa_tree_lt_8_21_groupi_n_30 ,in3[5] ,csa_tree_lt_8_21_groupi_n_21);
  or csa_tree_lt_8_21_groupi_g463__3680(csa_tree_lt_8_21_groupi_n_29 ,csa_tree_lt_8_21_groupi_n_7 ,csa_tree_lt_8_21_groupi_n_18);
  and csa_tree_lt_8_21_groupi_g464__1617(csa_tree_lt_8_21_groupi_n_34 ,in3[4] ,csa_tree_lt_8_21_groupi_n_16);
  or csa_tree_lt_8_21_groupi_g465__2802(csa_tree_lt_8_21_groupi_n_25 ,csa_tree_lt_8_21_groupi_n_6 ,csa_tree_lt_8_21_groupi_n_17);
  xnor csa_tree_lt_8_21_groupi_g466__1705(csa_tree_lt_8_21_groupi_n_24 ,in1[2] ,in2[2]);
  xor csa_tree_lt_8_21_groupi_g467__5122(csa_tree_lt_8_21_groupi_n_28 ,in3[3] ,in2[3]);
  or csa_tree_lt_8_21_groupi_g468__8246(csa_tree_lt_8_21_groupi_n_27 ,csa_tree_lt_8_21_groupi_n_22 ,csa_tree_lt_8_21_groupi_n_19);
  xnor csa_tree_lt_8_21_groupi_g469__7098(csa_tree_lt_8_21_groupi_n_23 ,in1[1] ,in2[1]);
  or csa_tree_lt_8_21_groupi_g470__6131(csa_tree_lt_8_21_groupi_n_26 ,csa_tree_lt_8_21_groupi_n_21 ,csa_tree_lt_8_21_groupi_n_10);
  or csa_tree_lt_8_21_groupi_g471__1881(csa_tree_lt_8_21_groupi_n_20 ,csa_tree_lt_8_21_groupi_n_4 ,in1[2]);
  nor csa_tree_lt_8_21_groupi_g472__5115(csa_tree_lt_8_21_groupi_n_19 ,csa_tree_lt_8_21_groupi_n_1 ,in3[6]);
  nor csa_tree_lt_8_21_groupi_g473__7482(csa_tree_lt_8_21_groupi_n_18 ,csa_tree_lt_8_21_groupi_n_0 ,in3[2]);
  nor csa_tree_lt_8_21_groupi_g474__4733(csa_tree_lt_8_21_groupi_n_17 ,csa_tree_lt_8_21_groupi_n_2 ,in3[1]);
  and csa_tree_lt_8_21_groupi_g475__6161(csa_tree_lt_8_21_groupi_n_22 ,in3[8] ,csa_tree_lt_8_21_groupi_n_1);
  and csa_tree_lt_8_21_groupi_g476__9315(csa_tree_lt_8_21_groupi_n_21 ,in3[6] ,csa_tree_lt_8_21_groupi_n_3);
  nor csa_tree_lt_8_21_groupi_g477__9945(csa_tree_lt_8_21_groupi_n_15 ,csa_tree_lt_8_21_groupi_n_1 ,in3[8]);
  or csa_tree_lt_8_21_groupi_g478__2883(csa_tree_lt_8_21_groupi_n_14 ,csa_tree_lt_8_21_groupi_n_5 ,in1[1]);
  nor csa_tree_lt_8_21_groupi_g479__2346(csa_tree_lt_8_21_groupi_n_13 ,csa_tree_lt_8_21_groupi_n_3 ,in3[6]);
  nor csa_tree_lt_8_21_groupi_g480__1666(csa_tree_lt_8_21_groupi_n_12 ,in3[0] ,in1[0]);
  and csa_tree_lt_8_21_groupi_g481__7410(csa_tree_lt_8_21_groupi_n_11 ,in3[0] ,in1[0]);
  nor csa_tree_lt_8_21_groupi_g482__6417(csa_tree_lt_8_21_groupi_n_10 ,csa_tree_lt_8_21_groupi_n_3 ,in3[4]);
  and csa_tree_lt_8_21_groupi_g483__5477(csa_tree_lt_8_21_groupi_n_16 ,csa_tree_lt_8_21_groupi_n_9 ,csa_tree_lt_8_21_groupi_n_8);
  not csa_tree_lt_8_21_groupi_g484(csa_tree_lt_8_21_groupi_n_9 ,in3[3]);
  not csa_tree_lt_8_21_groupi_g485(csa_tree_lt_8_21_groupi_n_8 ,in2[3]);
  not csa_tree_lt_8_21_groupi_g486(csa_tree_lt_8_21_groupi_n_7 ,in2[2]);
  not csa_tree_lt_8_21_groupi_g487(csa_tree_lt_8_21_groupi_n_6 ,in2[1]);
  not csa_tree_lt_8_21_groupi_g488(csa_tree_lt_8_21_groupi_n_5 ,in3[1]);
  not csa_tree_lt_8_21_groupi_g489(csa_tree_lt_8_21_groupi_n_4 ,in3[2]);
  not csa_tree_lt_8_21_groupi_g490(csa_tree_lt_8_21_groupi_n_3 ,in3[5]);
  not csa_tree_lt_8_21_groupi_g491(csa_tree_lt_8_21_groupi_n_2 ,in1[1]);
  not csa_tree_lt_8_21_groupi_g492(csa_tree_lt_8_21_groupi_n_1 ,in3[7]);
  not csa_tree_lt_8_21_groupi_g493(csa_tree_lt_8_21_groupi_n_0 ,in1[2]);

endmodule
